module LED64Enc ( clk, rst, Plaintext, Key, Ciphertext );
  input [63:0] Plaintext;
  input [63:0] Key;
  output [63:0] Ciphertext;
  (* FIRMER="clock" *)input clk;
  (* FIRMER="control" *)input rst;
  wire   SubCellInst_LFInst_0_LFInst_3_n16 ,
         SubCellInst_LFInst_0_LFInst_3_n15 ,
         SubCellInst_LFInst_0_LFInst_3_n14 ,
         SubCellInst_LFInst_0_LFInst_3_n13 ,
         SubCellInst_LFInst_0_LFInst_3_n12 ,
         SubCellInst_LFInst_0_LFInst_3_n11 ,
         SubCellInst_LFInst_0_LFInst_2_n22 ,
         SubCellInst_LFInst_0_LFInst_2_n21 ,
         SubCellInst_LFInst_0_LFInst_2_n20 ,
         SubCellInst_LFInst_0_LFInst_2_n19 ,
         SubCellInst_LFInst_0_LFInst_2_n18 ,
         SubCellInst_LFInst_0_LFInst_2_n17 ,
         SubCellInst_LFInst_0_LFInst_2_n16 ,
         SubCellInst_LFInst_0_LFInst_2_n15 ,
         SubCellInst_LFInst_0_LFInst_1_n18 ,
         SubCellInst_LFInst_0_LFInst_1_n17 ,
         SubCellInst_LFInst_0_LFInst_1_n16 ,
         SubCellInst_LFInst_0_LFInst_1_n15 ,
         SubCellInst_LFInst_0_LFInst_1_n14 ,
         SubCellInst_LFInst_0_LFInst_1_n13 ,
         SubCellInst_LFInst_0_LFInst_1_n12 ,
         SubCellInst_LFInst_0_LFInst_1_n11 ,
         SubCellInst_LFInst_0_LFInst_1_n10 ,
         SubCellInst_LFInst_0_LFInst_0_n6 ,
         SubCellInst_LFInst_0_LFInst_0_n5 ,
         SubCellInst_LFInst_0_LFInst_0_n4 ,
         SubCellInst_LFInst_1_LFInst_3_n16 ,
         SubCellInst_LFInst_1_LFInst_3_n15 ,
         SubCellInst_LFInst_1_LFInst_3_n14 ,
         SubCellInst_LFInst_1_LFInst_3_n13 ,
         SubCellInst_LFInst_1_LFInst_3_n12 ,
         SubCellInst_LFInst_1_LFInst_3_n11 ,
         SubCellInst_LFInst_1_LFInst_2_n22 ,
         SubCellInst_LFInst_1_LFInst_2_n21 ,
         SubCellInst_LFInst_1_LFInst_2_n20 ,
         SubCellInst_LFInst_1_LFInst_2_n19 ,
         SubCellInst_LFInst_1_LFInst_2_n18 ,
         SubCellInst_LFInst_1_LFInst_2_n17 ,
         SubCellInst_LFInst_1_LFInst_2_n16 ,
         SubCellInst_LFInst_1_LFInst_2_n15 ,
         SubCellInst_LFInst_1_LFInst_1_n18 ,
         SubCellInst_LFInst_1_LFInst_1_n17 ,
         SubCellInst_LFInst_1_LFInst_1_n16 ,
         SubCellInst_LFInst_1_LFInst_1_n15 ,
         SubCellInst_LFInst_1_LFInst_1_n14 ,
         SubCellInst_LFInst_1_LFInst_1_n13 ,
         SubCellInst_LFInst_1_LFInst_1_n12 ,
         SubCellInst_LFInst_1_LFInst_1_n11 ,
         SubCellInst_LFInst_1_LFInst_1_n10 ,
         SubCellInst_LFInst_1_LFInst_0_n6 ,
         SubCellInst_LFInst_1_LFInst_0_n5 ,
         SubCellInst_LFInst_1_LFInst_0_n4 ,
         SubCellInst_LFInst_2_LFInst_3_n16 ,
         SubCellInst_LFInst_2_LFInst_3_n15 ,
         SubCellInst_LFInst_2_LFInst_3_n14 ,
         SubCellInst_LFInst_2_LFInst_3_n13 ,
         SubCellInst_LFInst_2_LFInst_3_n12 ,
         SubCellInst_LFInst_2_LFInst_3_n11 ,
         SubCellInst_LFInst_2_LFInst_2_n22 ,
         SubCellInst_LFInst_2_LFInst_2_n21 ,
         SubCellInst_LFInst_2_LFInst_2_n20 ,
         SubCellInst_LFInst_2_LFInst_2_n19 ,
         SubCellInst_LFInst_2_LFInst_2_n18 ,
         SubCellInst_LFInst_2_LFInst_2_n17 ,
         SubCellInst_LFInst_2_LFInst_2_n16 ,
         SubCellInst_LFInst_2_LFInst_2_n15 ,
         SubCellInst_LFInst_2_LFInst_1_n18 ,
         SubCellInst_LFInst_2_LFInst_1_n17 ,
         SubCellInst_LFInst_2_LFInst_1_n16 ,
         SubCellInst_LFInst_2_LFInst_1_n15 ,
         SubCellInst_LFInst_2_LFInst_1_n14 ,
         SubCellInst_LFInst_2_LFInst_1_n13 ,
         SubCellInst_LFInst_2_LFInst_1_n12 ,
         SubCellInst_LFInst_2_LFInst_1_n11 ,
         SubCellInst_LFInst_2_LFInst_1_n10 ,
         SubCellInst_LFInst_2_LFInst_0_n6 ,
         SubCellInst_LFInst_2_LFInst_0_n5 ,
         SubCellInst_LFInst_2_LFInst_0_n4 ,
         SubCellInst_LFInst_3_LFInst_3_n16 ,
         SubCellInst_LFInst_3_LFInst_3_n15 ,
         SubCellInst_LFInst_3_LFInst_3_n14 ,
         SubCellInst_LFInst_3_LFInst_3_n13 ,
         SubCellInst_LFInst_3_LFInst_3_n12 ,
         SubCellInst_LFInst_3_LFInst_3_n11 ,
         SubCellInst_LFInst_3_LFInst_2_n22 ,
         SubCellInst_LFInst_3_LFInst_2_n21 ,
         SubCellInst_LFInst_3_LFInst_2_n20 ,
         SubCellInst_LFInst_3_LFInst_2_n19 ,
         SubCellInst_LFInst_3_LFInst_2_n18 ,
         SubCellInst_LFInst_3_LFInst_2_n17 ,
         SubCellInst_LFInst_3_LFInst_2_n16 ,
         SubCellInst_LFInst_3_LFInst_2_n15 ,
         SubCellInst_LFInst_3_LFInst_1_n18 ,
         SubCellInst_LFInst_3_LFInst_1_n17 ,
         SubCellInst_LFInst_3_LFInst_1_n16 ,
         SubCellInst_LFInst_3_LFInst_1_n15 ,
         SubCellInst_LFInst_3_LFInst_1_n14 ,
         SubCellInst_LFInst_3_LFInst_1_n13 ,
         SubCellInst_LFInst_3_LFInst_1_n12 ,
         SubCellInst_LFInst_3_LFInst_1_n11 ,
         SubCellInst_LFInst_3_LFInst_1_n10 ,
         SubCellInst_LFInst_3_LFInst_0_n6 ,
         SubCellInst_LFInst_3_LFInst_0_n5 ,
         SubCellInst_LFInst_3_LFInst_0_n4 ,
         SubCellInst_LFInst_4_LFInst_3_n16 ,
         SubCellInst_LFInst_4_LFInst_3_n15 ,
         SubCellInst_LFInst_4_LFInst_3_n14 ,
         SubCellInst_LFInst_4_LFInst_3_n13 ,
         SubCellInst_LFInst_4_LFInst_3_n12 ,
         SubCellInst_LFInst_4_LFInst_3_n11 ,
         SubCellInst_LFInst_4_LFInst_2_n22 ,
         SubCellInst_LFInst_4_LFInst_2_n21 ,
         SubCellInst_LFInst_4_LFInst_2_n20 ,
         SubCellInst_LFInst_4_LFInst_2_n19 ,
         SubCellInst_LFInst_4_LFInst_2_n18 ,
         SubCellInst_LFInst_4_LFInst_2_n17 ,
         SubCellInst_LFInst_4_LFInst_2_n16 ,
         SubCellInst_LFInst_4_LFInst_2_n15 ,
         SubCellInst_LFInst_4_LFInst_1_n18 ,
         SubCellInst_LFInst_4_LFInst_1_n17 ,
         SubCellInst_LFInst_4_LFInst_1_n16 ,
         SubCellInst_LFInst_4_LFInst_1_n15 ,
         SubCellInst_LFInst_4_LFInst_1_n14 ,
         SubCellInst_LFInst_4_LFInst_1_n13 ,
         SubCellInst_LFInst_4_LFInst_1_n12 ,
         SubCellInst_LFInst_4_LFInst_1_n11 ,
         SubCellInst_LFInst_4_LFInst_1_n10 ,
         SubCellInst_LFInst_4_LFInst_0_n6 ,
         SubCellInst_LFInst_4_LFInst_0_n5 ,
         SubCellInst_LFInst_4_LFInst_0_n4 ,
         SubCellInst_LFInst_5_LFInst_3_n16 ,
         SubCellInst_LFInst_5_LFInst_3_n15 ,
         SubCellInst_LFInst_5_LFInst_3_n14 ,
         SubCellInst_LFInst_5_LFInst_3_n13 ,
         SubCellInst_LFInst_5_LFInst_3_n12 ,
         SubCellInst_LFInst_5_LFInst_3_n11 ,
         SubCellInst_LFInst_5_LFInst_2_n22 ,
         SubCellInst_LFInst_5_LFInst_2_n21 ,
         SubCellInst_LFInst_5_LFInst_2_n20 ,
         SubCellInst_LFInst_5_LFInst_2_n19 ,
         SubCellInst_LFInst_5_LFInst_2_n18 ,
         SubCellInst_LFInst_5_LFInst_2_n17 ,
         SubCellInst_LFInst_5_LFInst_2_n16 ,
         SubCellInst_LFInst_5_LFInst_2_n15 ,
         SubCellInst_LFInst_5_LFInst_1_n18 ,
         SubCellInst_LFInst_5_LFInst_1_n17 ,
         SubCellInst_LFInst_5_LFInst_1_n16 ,
         SubCellInst_LFInst_5_LFInst_1_n15 ,
         SubCellInst_LFInst_5_LFInst_1_n14 ,
         SubCellInst_LFInst_5_LFInst_1_n13 ,
         SubCellInst_LFInst_5_LFInst_1_n12 ,
         SubCellInst_LFInst_5_LFInst_1_n11 ,
         SubCellInst_LFInst_5_LFInst_1_n10 ,
         SubCellInst_LFInst_5_LFInst_0_n6 ,
         SubCellInst_LFInst_5_LFInst_0_n5 ,
         SubCellInst_LFInst_5_LFInst_0_n4 ,
         SubCellInst_LFInst_6_LFInst_3_n16 ,
         SubCellInst_LFInst_6_LFInst_3_n15 ,
         SubCellInst_LFInst_6_LFInst_3_n14 ,
         SubCellInst_LFInst_6_LFInst_3_n13 ,
         SubCellInst_LFInst_6_LFInst_3_n12 ,
         SubCellInst_LFInst_6_LFInst_3_n11 ,
         SubCellInst_LFInst_6_LFInst_2_n22 ,
         SubCellInst_LFInst_6_LFInst_2_n21 ,
         SubCellInst_LFInst_6_LFInst_2_n20 ,
         SubCellInst_LFInst_6_LFInst_2_n19 ,
         SubCellInst_LFInst_6_LFInst_2_n18 ,
         SubCellInst_LFInst_6_LFInst_2_n17 ,
         SubCellInst_LFInst_6_LFInst_2_n16 ,
         SubCellInst_LFInst_6_LFInst_2_n15 ,
         SubCellInst_LFInst_6_LFInst_1_n18 ,
         SubCellInst_LFInst_6_LFInst_1_n17 ,
         SubCellInst_LFInst_6_LFInst_1_n16 ,
         SubCellInst_LFInst_6_LFInst_1_n15 ,
         SubCellInst_LFInst_6_LFInst_1_n14 ,
         SubCellInst_LFInst_6_LFInst_1_n13 ,
         SubCellInst_LFInst_6_LFInst_1_n12 ,
         SubCellInst_LFInst_6_LFInst_1_n11 ,
         SubCellInst_LFInst_6_LFInst_1_n10 ,
         SubCellInst_LFInst_6_LFInst_0_n6 ,
         SubCellInst_LFInst_6_LFInst_0_n5 ,
         SubCellInst_LFInst_6_LFInst_0_n4 ,
         SubCellInst_LFInst_7_LFInst_3_n16 ,
         SubCellInst_LFInst_7_LFInst_3_n15 ,
         SubCellInst_LFInst_7_LFInst_3_n14 ,
         SubCellInst_LFInst_7_LFInst_3_n13 ,
         SubCellInst_LFInst_7_LFInst_3_n12 ,
         SubCellInst_LFInst_7_LFInst_3_n11 ,
         SubCellInst_LFInst_7_LFInst_2_n22 ,
         SubCellInst_LFInst_7_LFInst_2_n21 ,
         SubCellInst_LFInst_7_LFInst_2_n20 ,
         SubCellInst_LFInst_7_LFInst_2_n19 ,
         SubCellInst_LFInst_7_LFInst_2_n18 ,
         SubCellInst_LFInst_7_LFInst_2_n17 ,
         SubCellInst_LFInst_7_LFInst_2_n16 ,
         SubCellInst_LFInst_7_LFInst_2_n15 ,
         SubCellInst_LFInst_7_LFInst_1_n18 ,
         SubCellInst_LFInst_7_LFInst_1_n17 ,
         SubCellInst_LFInst_7_LFInst_1_n16 ,
         SubCellInst_LFInst_7_LFInst_1_n15 ,
         SubCellInst_LFInst_7_LFInst_1_n14 ,
         SubCellInst_LFInst_7_LFInst_1_n13 ,
         SubCellInst_LFInst_7_LFInst_1_n12 ,
         SubCellInst_LFInst_7_LFInst_1_n11 ,
         SubCellInst_LFInst_7_LFInst_1_n10 ,
         SubCellInst_LFInst_7_LFInst_0_n6 ,
         SubCellInst_LFInst_7_LFInst_0_n5 ,
         SubCellInst_LFInst_7_LFInst_0_n4 ,
         SubCellInst_LFInst_8_LFInst_3_n16 ,
         SubCellInst_LFInst_8_LFInst_3_n15 ,
         SubCellInst_LFInst_8_LFInst_3_n14 ,
         SubCellInst_LFInst_8_LFInst_3_n13 ,
         SubCellInst_LFInst_8_LFInst_3_n12 ,
         SubCellInst_LFInst_8_LFInst_3_n11 ,
         SubCellInst_LFInst_8_LFInst_2_n22 ,
         SubCellInst_LFInst_8_LFInst_2_n21 ,
         SubCellInst_LFInst_8_LFInst_2_n20 ,
         SubCellInst_LFInst_8_LFInst_2_n19 ,
         SubCellInst_LFInst_8_LFInst_2_n18 ,
         SubCellInst_LFInst_8_LFInst_2_n17 ,
         SubCellInst_LFInst_8_LFInst_2_n16 ,
         SubCellInst_LFInst_8_LFInst_2_n15 ,
         SubCellInst_LFInst_8_LFInst_1_n18 ,
         SubCellInst_LFInst_8_LFInst_1_n17 ,
         SubCellInst_LFInst_8_LFInst_1_n16 ,
         SubCellInst_LFInst_8_LFInst_1_n15 ,
         SubCellInst_LFInst_8_LFInst_1_n14 ,
         SubCellInst_LFInst_8_LFInst_1_n13 ,
         SubCellInst_LFInst_8_LFInst_1_n12 ,
         SubCellInst_LFInst_8_LFInst_1_n11 ,
         SubCellInst_LFInst_8_LFInst_1_n10 ,
         SubCellInst_LFInst_8_LFInst_0_n6 ,
         SubCellInst_LFInst_8_LFInst_0_n5 ,
         SubCellInst_LFInst_8_LFInst_0_n4 ,
         SubCellInst_LFInst_9_LFInst_3_n16 ,
         SubCellInst_LFInst_9_LFInst_3_n15 ,
         SubCellInst_LFInst_9_LFInst_3_n14 ,
         SubCellInst_LFInst_9_LFInst_3_n13 ,
         SubCellInst_LFInst_9_LFInst_3_n12 ,
         SubCellInst_LFInst_9_LFInst_3_n11 ,
         SubCellInst_LFInst_9_LFInst_2_n22 ,
         SubCellInst_LFInst_9_LFInst_2_n21 ,
         SubCellInst_LFInst_9_LFInst_2_n20 ,
         SubCellInst_LFInst_9_LFInst_2_n19 ,
         SubCellInst_LFInst_9_LFInst_2_n18 ,
         SubCellInst_LFInst_9_LFInst_2_n17 ,
         SubCellInst_LFInst_9_LFInst_2_n16 ,
         SubCellInst_LFInst_9_LFInst_2_n15 ,
         SubCellInst_LFInst_9_LFInst_1_n18 ,
         SubCellInst_LFInst_9_LFInst_1_n17 ,
         SubCellInst_LFInst_9_LFInst_1_n16 ,
         SubCellInst_LFInst_9_LFInst_1_n15 ,
         SubCellInst_LFInst_9_LFInst_1_n14 ,
         SubCellInst_LFInst_9_LFInst_1_n13 ,
         SubCellInst_LFInst_9_LFInst_1_n12 ,
         SubCellInst_LFInst_9_LFInst_1_n11 ,
         SubCellInst_LFInst_9_LFInst_1_n10 ,
         SubCellInst_LFInst_9_LFInst_0_n6 ,
         SubCellInst_LFInst_9_LFInst_0_n5 ,
         SubCellInst_LFInst_9_LFInst_0_n4 ,
         SubCellInst_LFInst_10_LFInst_3_n16 ,
         SubCellInst_LFInst_10_LFInst_3_n15 ,
         SubCellInst_LFInst_10_LFInst_3_n14 ,
         SubCellInst_LFInst_10_LFInst_3_n13 ,
         SubCellInst_LFInst_10_LFInst_3_n12 ,
         SubCellInst_LFInst_10_LFInst_3_n11 ,
         SubCellInst_LFInst_10_LFInst_2_n22 ,
         SubCellInst_LFInst_10_LFInst_2_n21 ,
         SubCellInst_LFInst_10_LFInst_2_n20 ,
         SubCellInst_LFInst_10_LFInst_2_n19 ,
         SubCellInst_LFInst_10_LFInst_2_n18 ,
         SubCellInst_LFInst_10_LFInst_2_n17 ,
         SubCellInst_LFInst_10_LFInst_2_n16 ,
         SubCellInst_LFInst_10_LFInst_2_n15 ,
         SubCellInst_LFInst_10_LFInst_1_n18 ,
         SubCellInst_LFInst_10_LFInst_1_n17 ,
         SubCellInst_LFInst_10_LFInst_1_n16 ,
         SubCellInst_LFInst_10_LFInst_1_n15 ,
         SubCellInst_LFInst_10_LFInst_1_n14 ,
         SubCellInst_LFInst_10_LFInst_1_n13 ,
         SubCellInst_LFInst_10_LFInst_1_n12 ,
         SubCellInst_LFInst_10_LFInst_1_n11 ,
         SubCellInst_LFInst_10_LFInst_1_n10 ,
         SubCellInst_LFInst_10_LFInst_0_n6 ,
         SubCellInst_LFInst_10_LFInst_0_n5 ,
         SubCellInst_LFInst_10_LFInst_0_n4 ,
         SubCellInst_LFInst_11_LFInst_3_n16 ,
         SubCellInst_LFInst_11_LFInst_3_n15 ,
         SubCellInst_LFInst_11_LFInst_3_n14 ,
         SubCellInst_LFInst_11_LFInst_3_n13 ,
         SubCellInst_LFInst_11_LFInst_3_n12 ,
         SubCellInst_LFInst_11_LFInst_3_n11 ,
         SubCellInst_LFInst_11_LFInst_2_n22 ,
         SubCellInst_LFInst_11_LFInst_2_n21 ,
         SubCellInst_LFInst_11_LFInst_2_n20 ,
         SubCellInst_LFInst_11_LFInst_2_n19 ,
         SubCellInst_LFInst_11_LFInst_2_n18 ,
         SubCellInst_LFInst_11_LFInst_2_n17 ,
         SubCellInst_LFInst_11_LFInst_2_n16 ,
         SubCellInst_LFInst_11_LFInst_2_n15 ,
         SubCellInst_LFInst_11_LFInst_1_n18 ,
         SubCellInst_LFInst_11_LFInst_1_n17 ,
         SubCellInst_LFInst_11_LFInst_1_n16 ,
         SubCellInst_LFInst_11_LFInst_1_n15 ,
         SubCellInst_LFInst_11_LFInst_1_n14 ,
         SubCellInst_LFInst_11_LFInst_1_n13 ,
         SubCellInst_LFInst_11_LFInst_1_n12 ,
         SubCellInst_LFInst_11_LFInst_1_n11 ,
         SubCellInst_LFInst_11_LFInst_1_n10 ,
         SubCellInst_LFInst_11_LFInst_0_n6 ,
         SubCellInst_LFInst_11_LFInst_0_n5 ,
         SubCellInst_LFInst_11_LFInst_0_n4 ,
         SubCellInst_LFInst_12_LFInst_3_n16 ,
         SubCellInst_LFInst_12_LFInst_3_n15 ,
         SubCellInst_LFInst_12_LFInst_3_n14 ,
         SubCellInst_LFInst_12_LFInst_3_n13 ,
         SubCellInst_LFInst_12_LFInst_3_n12 ,
         SubCellInst_LFInst_12_LFInst_3_n11 ,
         SubCellInst_LFInst_12_LFInst_2_n22 ,
         SubCellInst_LFInst_12_LFInst_2_n21 ,
         SubCellInst_LFInst_12_LFInst_2_n20 ,
         SubCellInst_LFInst_12_LFInst_2_n19 ,
         SubCellInst_LFInst_12_LFInst_2_n18 ,
         SubCellInst_LFInst_12_LFInst_2_n17 ,
         SubCellInst_LFInst_12_LFInst_2_n16 ,
         SubCellInst_LFInst_12_LFInst_2_n15 ,
         SubCellInst_LFInst_12_LFInst_1_n18 ,
         SubCellInst_LFInst_12_LFInst_1_n17 ,
         SubCellInst_LFInst_12_LFInst_1_n16 ,
         SubCellInst_LFInst_12_LFInst_1_n15 ,
         SubCellInst_LFInst_12_LFInst_1_n14 ,
         SubCellInst_LFInst_12_LFInst_1_n13 ,
         SubCellInst_LFInst_12_LFInst_1_n12 ,
         SubCellInst_LFInst_12_LFInst_1_n11 ,
         SubCellInst_LFInst_12_LFInst_1_n10 ,
         SubCellInst_LFInst_12_LFInst_0_n6 ,
         SubCellInst_LFInst_12_LFInst_0_n5 ,
         SubCellInst_LFInst_12_LFInst_0_n4 ,
         SubCellInst_LFInst_13_LFInst_3_n16 ,
         SubCellInst_LFInst_13_LFInst_3_n15 ,
         SubCellInst_LFInst_13_LFInst_3_n14 ,
         SubCellInst_LFInst_13_LFInst_3_n13 ,
         SubCellInst_LFInst_13_LFInst_3_n12 ,
         SubCellInst_LFInst_13_LFInst_3_n11 ,
         SubCellInst_LFInst_13_LFInst_2_n22 ,
         SubCellInst_LFInst_13_LFInst_2_n21 ,
         SubCellInst_LFInst_13_LFInst_2_n20 ,
         SubCellInst_LFInst_13_LFInst_2_n19 ,
         SubCellInst_LFInst_13_LFInst_2_n18 ,
         SubCellInst_LFInst_13_LFInst_2_n17 ,
         SubCellInst_LFInst_13_LFInst_2_n16 ,
         SubCellInst_LFInst_13_LFInst_2_n15 ,
         SubCellInst_LFInst_13_LFInst_1_n18 ,
         SubCellInst_LFInst_13_LFInst_1_n17 ,
         SubCellInst_LFInst_13_LFInst_1_n16 ,
         SubCellInst_LFInst_13_LFInst_1_n15 ,
         SubCellInst_LFInst_13_LFInst_1_n14 ,
         SubCellInst_LFInst_13_LFInst_1_n13 ,
         SubCellInst_LFInst_13_LFInst_1_n12 ,
         SubCellInst_LFInst_13_LFInst_1_n11 ,
         SubCellInst_LFInst_13_LFInst_1_n10 ,
         SubCellInst_LFInst_13_LFInst_0_n6 ,
         SubCellInst_LFInst_13_LFInst_0_n5 ,
         SubCellInst_LFInst_13_LFInst_0_n4 ,
         SubCellInst_LFInst_14_LFInst_3_n16 ,
         SubCellInst_LFInst_14_LFInst_3_n15 ,
         SubCellInst_LFInst_14_LFInst_3_n14 ,
         SubCellInst_LFInst_14_LFInst_3_n13 ,
         SubCellInst_LFInst_14_LFInst_3_n12 ,
         SubCellInst_LFInst_14_LFInst_3_n11 ,
         SubCellInst_LFInst_14_LFInst_2_n22 ,
         SubCellInst_LFInst_14_LFInst_2_n21 ,
         SubCellInst_LFInst_14_LFInst_2_n20 ,
         SubCellInst_LFInst_14_LFInst_2_n19 ,
         SubCellInst_LFInst_14_LFInst_2_n18 ,
         SubCellInst_LFInst_14_LFInst_2_n17 ,
         SubCellInst_LFInst_14_LFInst_2_n16 ,
         SubCellInst_LFInst_14_LFInst_2_n15 ,
         SubCellInst_LFInst_14_LFInst_1_n18 ,
         SubCellInst_LFInst_14_LFInst_1_n17 ,
         SubCellInst_LFInst_14_LFInst_1_n16 ,
         SubCellInst_LFInst_14_LFInst_1_n15 ,
         SubCellInst_LFInst_14_LFInst_1_n14 ,
         SubCellInst_LFInst_14_LFInst_1_n13 ,
         SubCellInst_LFInst_14_LFInst_1_n12 ,
         SubCellInst_LFInst_14_LFInst_1_n11 ,
         SubCellInst_LFInst_14_LFInst_1_n10 ,
         SubCellInst_LFInst_14_LFInst_0_n6 ,
         SubCellInst_LFInst_14_LFInst_0_n5 ,
         SubCellInst_LFInst_14_LFInst_0_n4 ,
         SubCellInst_LFInst_15_LFInst_3_n16 ,
         SubCellInst_LFInst_15_LFInst_3_n15 ,
         SubCellInst_LFInst_15_LFInst_3_n14 ,
         SubCellInst_LFInst_15_LFInst_3_n13 ,
         SubCellInst_LFInst_15_LFInst_3_n12 ,
         SubCellInst_LFInst_15_LFInst_3_n11 ,
         SubCellInst_LFInst_15_LFInst_2_n22 ,
         SubCellInst_LFInst_15_LFInst_2_n21 ,
         SubCellInst_LFInst_15_LFInst_2_n20 ,
         SubCellInst_LFInst_15_LFInst_2_n19 ,
         SubCellInst_LFInst_15_LFInst_2_n18 ,
         SubCellInst_LFInst_15_LFInst_2_n17 ,
         SubCellInst_LFInst_15_LFInst_2_n16 ,
         SubCellInst_LFInst_15_LFInst_2_n15 ,
         SubCellInst_LFInst_15_LFInst_1_n18 ,
         SubCellInst_LFInst_15_LFInst_1_n17 ,
         SubCellInst_LFInst_15_LFInst_1_n16 ,
         SubCellInst_LFInst_15_LFInst_1_n15 ,
         SubCellInst_LFInst_15_LFInst_1_n14 ,
         SubCellInst_LFInst_15_LFInst_1_n13 ,
         SubCellInst_LFInst_15_LFInst_1_n12 ,
         SubCellInst_LFInst_15_LFInst_1_n11 ,
         SubCellInst_LFInst_15_LFInst_1_n10 ,
         SubCellInst_LFInst_15_LFInst_0_n6 ,
         SubCellInst_LFInst_15_LFInst_0_n5 ,
         SubCellInst_LFInst_15_LFInst_0_n4 , MCInst1_MC0_v0_2Inst_0_n2 ,
         MCInst1_MC0_v1_2Inst_0_n2 , MCInst1_MC0_v2_3Inst_0_n4 ,
         MCInst1_MC0_v2_3Inst_0_n3 , MCInst1_MC0_v3_3Inst_0_n2 ,
         MCInst1_MC0_v0_2Inst_1_n2 , MCInst1_MC0_v2_1Inst_1_n2 ,
         MCInst1_MC0_v2_2Inst_1_n4 , MCInst1_MC0_v2_2Inst_1_n3 ,
         MCInst1_MC0_v3_3Inst_1_n2 , MCInst1_MC0_v1_1Inst_2_n2 ,
         MCInst1_MC0_v1_2Inst_2_n2 , MCInst1_MC0_v2_1Inst_2_n2 ,
         MCInst1_MC0_v2_2Inst_2_n2 , MCInst1_MC0_v3_1Inst_2_n2 ,
         MCInst1_MC0_v1_2Inst_3_n4 , MCInst1_MC0_v1_2Inst_3_n3 ,
         MCInst1_MC0_v2_2Inst_3_n2 , MCInst1_MC0_v2_3Inst_3_n2 ,
         MCInst1_MC0_r0Inst_XORInst_0_0_n5 ,
         MCInst1_MC0_r0Inst_XORInst_0_0_n4 ,
         MCInst1_MC0_r0Inst_XORInst_0_1_n5 ,
         MCInst1_MC0_r0Inst_XORInst_0_1_n4 ,
         MCInst1_MC0_r0Inst_XORInst_0_2_n5 ,
         MCInst1_MC0_r0Inst_XORInst_0_2_n4 ,
         MCInst1_MC0_r0Inst_XORInst_0_3_n5 ,
         MCInst1_MC0_r0Inst_XORInst_0_3_n4 ,
         MCInst1_MC0_r1Inst_XORInst_0_0_n5 ,
         MCInst1_MC0_r1Inst_XORInst_0_0_n4 ,
         MCInst1_MC0_r1Inst_XORInst_0_1_n5 ,
         MCInst1_MC0_r1Inst_XORInst_0_1_n4 ,
         MCInst1_MC0_r1Inst_XORInst_0_2_n5 ,
         MCInst1_MC0_r1Inst_XORInst_0_2_n4 ,
         MCInst1_MC0_r1Inst_XORInst_0_3_n5 ,
         MCInst1_MC0_r1Inst_XORInst_0_3_n4 ,
         MCInst1_MC0_r2Inst_XORInst_0_0_n5 ,
         MCInst1_MC0_r2Inst_XORInst_0_0_n4 ,
         MCInst1_MC0_r2Inst_XORInst_0_1_n5 ,
         MCInst1_MC0_r2Inst_XORInst_0_1_n4 ,
         MCInst1_MC0_r2Inst_XORInst_0_2_n5 ,
         MCInst1_MC0_r2Inst_XORInst_0_2_n4 ,
         MCInst1_MC0_r2Inst_XORInst_0_3_n5 ,
         MCInst1_MC0_r2Inst_XORInst_0_3_n4 ,
         MCInst1_MC0_r3Inst_XORInst_0_0_n5 ,
         MCInst1_MC0_r3Inst_XORInst_0_0_n4 ,
         MCInst1_MC0_r3Inst_XORInst_0_1_n5 ,
         MCInst1_MC0_r3Inst_XORInst_0_1_n4 ,
         MCInst1_MC0_r3Inst_XORInst_0_2_n5 ,
         MCInst1_MC0_r3Inst_XORInst_0_2_n4 ,
         MCInst1_MC0_r3Inst_XORInst_0_3_n5 ,
         MCInst1_MC0_r3Inst_XORInst_0_3_n4 , MCInst1_MC1_v0_2Inst_0_n2 ,
         MCInst1_MC1_v1_2Inst_0_n2 , MCInst1_MC1_v2_3Inst_0_n4 ,
         MCInst1_MC1_v2_3Inst_0_n3 , MCInst1_MC1_v3_3Inst_0_n2 ,
         MCInst1_MC1_v0_2Inst_1_n2 , MCInst1_MC1_v2_1Inst_1_n2 ,
         MCInst1_MC1_v2_2Inst_1_n4 , MCInst1_MC1_v2_2Inst_1_n3 ,
         MCInst1_MC1_v3_3Inst_1_n2 , MCInst1_MC1_v1_1Inst_2_n2 ,
         MCInst1_MC1_v1_2Inst_2_n2 , MCInst1_MC1_v2_1Inst_2_n2 ,
         MCInst1_MC1_v2_2Inst_2_n2 , MCInst1_MC1_v3_1Inst_2_n2 ,
         MCInst1_MC1_v1_2Inst_3_n4 , MCInst1_MC1_v1_2Inst_3_n3 ,
         MCInst1_MC1_v2_2Inst_3_n2 , MCInst1_MC1_v2_3Inst_3_n2 ,
         MCInst1_MC1_r0Inst_XORInst_0_0_n5 ,
         MCInst1_MC1_r0Inst_XORInst_0_0_n4 ,
         MCInst1_MC1_r0Inst_XORInst_0_1_n5 ,
         MCInst1_MC1_r0Inst_XORInst_0_1_n4 ,
         MCInst1_MC1_r0Inst_XORInst_0_2_n5 ,
         MCInst1_MC1_r0Inst_XORInst_0_2_n4 ,
         MCInst1_MC1_r0Inst_XORInst_0_3_n5 ,
         MCInst1_MC1_r0Inst_XORInst_0_3_n4 ,
         MCInst1_MC1_r1Inst_XORInst_0_0_n5 ,
         MCInst1_MC1_r1Inst_XORInst_0_0_n4 ,
         MCInst1_MC1_r1Inst_XORInst_0_1_n5 ,
         MCInst1_MC1_r1Inst_XORInst_0_1_n4 ,
         MCInst1_MC1_r1Inst_XORInst_0_2_n5 ,
         MCInst1_MC1_r1Inst_XORInst_0_2_n4 ,
         MCInst1_MC1_r1Inst_XORInst_0_3_n5 ,
         MCInst1_MC1_r1Inst_XORInst_0_3_n4 ,
         MCInst1_MC1_r2Inst_XORInst_0_0_n5 ,
         MCInst1_MC1_r2Inst_XORInst_0_0_n4 ,
         MCInst1_MC1_r2Inst_XORInst_0_1_n5 ,
         MCInst1_MC1_r2Inst_XORInst_0_1_n4 ,
         MCInst1_MC1_r2Inst_XORInst_0_2_n5 ,
         MCInst1_MC1_r2Inst_XORInst_0_2_n4 ,
         MCInst1_MC1_r2Inst_XORInst_0_3_n5 ,
         MCInst1_MC1_r2Inst_XORInst_0_3_n4 ,
         MCInst1_MC1_r3Inst_XORInst_0_0_n5 ,
         MCInst1_MC1_r3Inst_XORInst_0_0_n4 ,
         MCInst1_MC1_r3Inst_XORInst_0_1_n5 ,
         MCInst1_MC1_r3Inst_XORInst_0_1_n4 ,
         MCInst1_MC1_r3Inst_XORInst_0_2_n5 ,
         MCInst1_MC1_r3Inst_XORInst_0_2_n4 ,
         MCInst1_MC1_r3Inst_XORInst_0_3_n5 ,
         MCInst1_MC1_r3Inst_XORInst_0_3_n4 , MCInst1_MC2_v0_2Inst_0_n2 ,
         MCInst1_MC2_v1_2Inst_0_n2 , MCInst1_MC2_v2_3Inst_0_n4 ,
         MCInst1_MC2_v2_3Inst_0_n3 , MCInst1_MC2_v3_3Inst_0_n2 ,
         MCInst1_MC2_v0_2Inst_1_n2 , MCInst1_MC2_v2_1Inst_1_n2 ,
         MCInst1_MC2_v2_2Inst_1_n4 , MCInst1_MC2_v2_2Inst_1_n3 ,
         MCInst1_MC2_v3_3Inst_1_n2 , MCInst1_MC2_v1_1Inst_2_n2 ,
         MCInst1_MC2_v1_2Inst_2_n2 , MCInst1_MC2_v2_1Inst_2_n2 ,
         MCInst1_MC2_v2_2Inst_2_n2 , MCInst1_MC2_v3_1Inst_2_n2 ,
         MCInst1_MC2_v1_2Inst_3_n4 , MCInst1_MC2_v1_2Inst_3_n3 ,
         MCInst1_MC2_v2_2Inst_3_n2 , MCInst1_MC2_v2_3Inst_3_n2 ,
         MCInst1_MC2_r0Inst_XORInst_0_0_n5 ,
         MCInst1_MC2_r0Inst_XORInst_0_0_n4 ,
         MCInst1_MC2_r0Inst_XORInst_0_1_n5 ,
         MCInst1_MC2_r0Inst_XORInst_0_1_n4 ,
         MCInst1_MC2_r0Inst_XORInst_0_2_n5 ,
         MCInst1_MC2_r0Inst_XORInst_0_2_n4 ,
         MCInst1_MC2_r0Inst_XORInst_0_3_n5 ,
         MCInst1_MC2_r0Inst_XORInst_0_3_n4 ,
         MCInst1_MC2_r1Inst_XORInst_0_0_n5 ,
         MCInst1_MC2_r1Inst_XORInst_0_0_n4 ,
         MCInst1_MC2_r1Inst_XORInst_0_1_n5 ,
         MCInst1_MC2_r1Inst_XORInst_0_1_n4 ,
         MCInst1_MC2_r1Inst_XORInst_0_2_n5 ,
         MCInst1_MC2_r1Inst_XORInst_0_2_n4 ,
         MCInst1_MC2_r1Inst_XORInst_0_3_n5 ,
         MCInst1_MC2_r1Inst_XORInst_0_3_n4 ,
         MCInst1_MC2_r2Inst_XORInst_0_0_n5 ,
         MCInst1_MC2_r2Inst_XORInst_0_0_n4 ,
         MCInst1_MC2_r2Inst_XORInst_0_1_n5 ,
         MCInst1_MC2_r2Inst_XORInst_0_1_n4 ,
         MCInst1_MC2_r2Inst_XORInst_0_2_n5 ,
         MCInst1_MC2_r2Inst_XORInst_0_2_n4 ,
         MCInst1_MC2_r2Inst_XORInst_0_3_n5 ,
         MCInst1_MC2_r2Inst_XORInst_0_3_n4 ,
         MCInst1_MC2_r3Inst_XORInst_0_0_n5 ,
         MCInst1_MC2_r3Inst_XORInst_0_0_n4 ,
         MCInst1_MC2_r3Inst_XORInst_0_1_n5 ,
         MCInst1_MC2_r3Inst_XORInst_0_1_n4 ,
         MCInst1_MC2_r3Inst_XORInst_0_2_n5 ,
         MCInst1_MC2_r3Inst_XORInst_0_2_n4 ,
         MCInst1_MC2_r3Inst_XORInst_0_3_n5 ,
         MCInst1_MC2_r3Inst_XORInst_0_3_n4 , MCInst1_MC3_v0_2Inst_0_n2 ,
         MCInst1_MC3_v1_2Inst_0_n2 , MCInst1_MC3_v2_3Inst_0_n4 ,
         MCInst1_MC3_v2_3Inst_0_n3 , MCInst1_MC3_v3_3Inst_0_n2 ,
         MCInst1_MC3_v0_2Inst_1_n2 , MCInst1_MC3_v2_1Inst_1_n2 ,
         MCInst1_MC3_v2_2Inst_1_n4 , MCInst1_MC3_v2_2Inst_1_n3 ,
         MCInst1_MC3_v3_3Inst_1_n2 , MCInst1_MC3_v1_1Inst_2_n2 ,
         MCInst1_MC3_v1_2Inst_2_n2 , MCInst1_MC3_v2_1Inst_2_n2 ,
         MCInst1_MC3_v2_2Inst_2_n2 , MCInst1_MC3_v3_1Inst_2_n2 ,
         MCInst1_MC3_v1_2Inst_3_n4 , MCInst1_MC3_v1_2Inst_3_n3 ,
         MCInst1_MC3_v2_2Inst_3_n2 , MCInst1_MC3_v2_3Inst_3_n2 ,
         MCInst1_MC3_r0Inst_XORInst_0_0_n5 ,
         MCInst1_MC3_r0Inst_XORInst_0_0_n4 ,
         MCInst1_MC3_r0Inst_XORInst_0_1_n5 ,
         MCInst1_MC3_r0Inst_XORInst_0_1_n4 ,
         MCInst1_MC3_r0Inst_XORInst_0_2_n5 ,
         MCInst1_MC3_r0Inst_XORInst_0_2_n4 ,
         MCInst1_MC3_r0Inst_XORInst_0_3_n5 ,
         MCInst1_MC3_r0Inst_XORInst_0_3_n4 ,
         MCInst1_MC3_r1Inst_XORInst_0_0_n5 ,
         MCInst1_MC3_r1Inst_XORInst_0_0_n4 ,
         MCInst1_MC3_r1Inst_XORInst_0_1_n5 ,
         MCInst1_MC3_r1Inst_XORInst_0_1_n4 ,
         MCInst1_MC3_r1Inst_XORInst_0_2_n5 ,
         MCInst1_MC3_r1Inst_XORInst_0_2_n4 ,
         MCInst1_MC3_r1Inst_XORInst_0_3_n5 ,
         MCInst1_MC3_r1Inst_XORInst_0_3_n4 ,
         MCInst1_MC3_r2Inst_XORInst_0_0_n5 ,
         MCInst1_MC3_r2Inst_XORInst_0_0_n4 ,
         MCInst1_MC3_r2Inst_XORInst_0_1_n5 ,
         MCInst1_MC3_r2Inst_XORInst_0_1_n4 ,
         MCInst1_MC3_r2Inst_XORInst_0_2_n5 ,
         MCInst1_MC3_r2Inst_XORInst_0_2_n4 ,
         MCInst1_MC3_r2Inst_XORInst_0_3_n5 ,
         MCInst1_MC3_r2Inst_XORInst_0_3_n4 ,
         MCInst1_MC3_r3Inst_XORInst_0_0_n5 ,
         MCInst1_MC3_r3Inst_XORInst_0_0_n4 ,
         MCInst1_MC3_r3Inst_XORInst_0_1_n5 ,
         MCInst1_MC3_r3Inst_XORInst_0_1_n4 ,
         MCInst1_MC3_r3Inst_XORInst_0_2_n5 ,
         MCInst1_MC3_r3Inst_XORInst_0_2_n4 ,
         MCInst1_MC3_r3Inst_XORInst_0_3_n5 ,
         MCInst1_MC3_r3Inst_XORInst_0_3_n4 ,
         SubCellInst2_LFInst_0_LFInst_3_n16 ,
         SubCellInst2_LFInst_0_LFInst_3_n15 ,
         SubCellInst2_LFInst_0_LFInst_3_n14 ,
         SubCellInst2_LFInst_0_LFInst_3_n13 ,
         SubCellInst2_LFInst_0_LFInst_3_n12 ,
         SubCellInst2_LFInst_0_LFInst_3_n11 ,
         SubCellInst2_LFInst_0_LFInst_2_n22 ,
         SubCellInst2_LFInst_0_LFInst_2_n21 ,
         SubCellInst2_LFInst_0_LFInst_2_n20 ,
         SubCellInst2_LFInst_0_LFInst_2_n19 ,
         SubCellInst2_LFInst_0_LFInst_2_n18 ,
         SubCellInst2_LFInst_0_LFInst_2_n17 ,
         SubCellInst2_LFInst_0_LFInst_2_n16 ,
         SubCellInst2_LFInst_0_LFInst_2_n15 ,
         SubCellInst2_LFInst_0_LFInst_1_n18 ,
         SubCellInst2_LFInst_0_LFInst_1_n17 ,
         SubCellInst2_LFInst_0_LFInst_1_n16 ,
         SubCellInst2_LFInst_0_LFInst_1_n15 ,
         SubCellInst2_LFInst_0_LFInst_1_n14 ,
         SubCellInst2_LFInst_0_LFInst_1_n13 ,
         SubCellInst2_LFInst_0_LFInst_1_n12 ,
         SubCellInst2_LFInst_0_LFInst_1_n11 ,
         SubCellInst2_LFInst_0_LFInst_1_n10 ,
         SubCellInst2_LFInst_0_LFInst_0_n6 ,
         SubCellInst2_LFInst_0_LFInst_0_n5 ,
         SubCellInst2_LFInst_0_LFInst_0_n4 ,
         SubCellInst2_LFInst_1_LFInst_3_n16 ,
         SubCellInst2_LFInst_1_LFInst_3_n15 ,
         SubCellInst2_LFInst_1_LFInst_3_n14 ,
         SubCellInst2_LFInst_1_LFInst_3_n13 ,
         SubCellInst2_LFInst_1_LFInst_3_n12 ,
         SubCellInst2_LFInst_1_LFInst_3_n11 ,
         SubCellInst2_LFInst_1_LFInst_2_n22 ,
         SubCellInst2_LFInst_1_LFInst_2_n21 ,
         SubCellInst2_LFInst_1_LFInst_2_n20 ,
         SubCellInst2_LFInst_1_LFInst_2_n19 ,
         SubCellInst2_LFInst_1_LFInst_2_n18 ,
         SubCellInst2_LFInst_1_LFInst_2_n17 ,
         SubCellInst2_LFInst_1_LFInst_2_n16 ,
         SubCellInst2_LFInst_1_LFInst_2_n15 ,
         SubCellInst2_LFInst_1_LFInst_1_n18 ,
         SubCellInst2_LFInst_1_LFInst_1_n17 ,
         SubCellInst2_LFInst_1_LFInst_1_n16 ,
         SubCellInst2_LFInst_1_LFInst_1_n15 ,
         SubCellInst2_LFInst_1_LFInst_1_n14 ,
         SubCellInst2_LFInst_1_LFInst_1_n13 ,
         SubCellInst2_LFInst_1_LFInst_1_n12 ,
         SubCellInst2_LFInst_1_LFInst_1_n11 ,
         SubCellInst2_LFInst_1_LFInst_1_n10 ,
         SubCellInst2_LFInst_1_LFInst_0_n6 ,
         SubCellInst2_LFInst_1_LFInst_0_n5 ,
         SubCellInst2_LFInst_1_LFInst_0_n4 ,
         SubCellInst2_LFInst_2_LFInst_3_n16 ,
         SubCellInst2_LFInst_2_LFInst_3_n15 ,
         SubCellInst2_LFInst_2_LFInst_3_n14 ,
         SubCellInst2_LFInst_2_LFInst_3_n13 ,
         SubCellInst2_LFInst_2_LFInst_3_n12 ,
         SubCellInst2_LFInst_2_LFInst_3_n11 ,
         SubCellInst2_LFInst_2_LFInst_2_n22 ,
         SubCellInst2_LFInst_2_LFInst_2_n21 ,
         SubCellInst2_LFInst_2_LFInst_2_n20 ,
         SubCellInst2_LFInst_2_LFInst_2_n19 ,
         SubCellInst2_LFInst_2_LFInst_2_n18 ,
         SubCellInst2_LFInst_2_LFInst_2_n17 ,
         SubCellInst2_LFInst_2_LFInst_2_n16 ,
         SubCellInst2_LFInst_2_LFInst_2_n15 ,
         SubCellInst2_LFInst_2_LFInst_1_n18 ,
         SubCellInst2_LFInst_2_LFInst_1_n17 ,
         SubCellInst2_LFInst_2_LFInst_1_n16 ,
         SubCellInst2_LFInst_2_LFInst_1_n15 ,
         SubCellInst2_LFInst_2_LFInst_1_n14 ,
         SubCellInst2_LFInst_2_LFInst_1_n13 ,
         SubCellInst2_LFInst_2_LFInst_1_n12 ,
         SubCellInst2_LFInst_2_LFInst_1_n11 ,
         SubCellInst2_LFInst_2_LFInst_1_n10 ,
         SubCellInst2_LFInst_2_LFInst_0_n6 ,
         SubCellInst2_LFInst_2_LFInst_0_n5 ,
         SubCellInst2_LFInst_2_LFInst_0_n4 ,
         SubCellInst2_LFInst_3_LFInst_3_n16 ,
         SubCellInst2_LFInst_3_LFInst_3_n15 ,
         SubCellInst2_LFInst_3_LFInst_3_n14 ,
         SubCellInst2_LFInst_3_LFInst_3_n13 ,
         SubCellInst2_LFInst_3_LFInst_3_n12 ,
         SubCellInst2_LFInst_3_LFInst_3_n11 ,
         SubCellInst2_LFInst_3_LFInst_2_n22 ,
         SubCellInst2_LFInst_3_LFInst_2_n21 ,
         SubCellInst2_LFInst_3_LFInst_2_n20 ,
         SubCellInst2_LFInst_3_LFInst_2_n19 ,
         SubCellInst2_LFInst_3_LFInst_2_n18 ,
         SubCellInst2_LFInst_3_LFInst_2_n17 ,
         SubCellInst2_LFInst_3_LFInst_2_n16 ,
         SubCellInst2_LFInst_3_LFInst_2_n15 ,
         SubCellInst2_LFInst_3_LFInst_1_n18 ,
         SubCellInst2_LFInst_3_LFInst_1_n17 ,
         SubCellInst2_LFInst_3_LFInst_1_n16 ,
         SubCellInst2_LFInst_3_LFInst_1_n15 ,
         SubCellInst2_LFInst_3_LFInst_1_n14 ,
         SubCellInst2_LFInst_3_LFInst_1_n13 ,
         SubCellInst2_LFInst_3_LFInst_1_n12 ,
         SubCellInst2_LFInst_3_LFInst_1_n11 ,
         SubCellInst2_LFInst_3_LFInst_1_n10 ,
         SubCellInst2_LFInst_3_LFInst_0_n6 ,
         SubCellInst2_LFInst_3_LFInst_0_n5 ,
         SubCellInst2_LFInst_3_LFInst_0_n4 ,
         SubCellInst2_LFInst_4_LFInst_3_n16 ,
         SubCellInst2_LFInst_4_LFInst_3_n15 ,
         SubCellInst2_LFInst_4_LFInst_3_n14 ,
         SubCellInst2_LFInst_4_LFInst_3_n13 ,
         SubCellInst2_LFInst_4_LFInst_3_n12 ,
         SubCellInst2_LFInst_4_LFInst_3_n11 ,
         SubCellInst2_LFInst_4_LFInst_2_n22 ,
         SubCellInst2_LFInst_4_LFInst_2_n21 ,
         SubCellInst2_LFInst_4_LFInst_2_n20 ,
         SubCellInst2_LFInst_4_LFInst_2_n19 ,
         SubCellInst2_LFInst_4_LFInst_2_n18 ,
         SubCellInst2_LFInst_4_LFInst_2_n17 ,
         SubCellInst2_LFInst_4_LFInst_2_n16 ,
         SubCellInst2_LFInst_4_LFInst_2_n15 ,
         SubCellInst2_LFInst_4_LFInst_1_n18 ,
         SubCellInst2_LFInst_4_LFInst_1_n17 ,
         SubCellInst2_LFInst_4_LFInst_1_n16 ,
         SubCellInst2_LFInst_4_LFInst_1_n15 ,
         SubCellInst2_LFInst_4_LFInst_1_n14 ,
         SubCellInst2_LFInst_4_LFInst_1_n13 ,
         SubCellInst2_LFInst_4_LFInst_1_n12 ,
         SubCellInst2_LFInst_4_LFInst_1_n11 ,
         SubCellInst2_LFInst_4_LFInst_1_n10 ,
         SubCellInst2_LFInst_4_LFInst_0_n6 ,
         SubCellInst2_LFInst_4_LFInst_0_n5 ,
         SubCellInst2_LFInst_4_LFInst_0_n4 ,
         SubCellInst2_LFInst_5_LFInst_3_n16 ,
         SubCellInst2_LFInst_5_LFInst_3_n15 ,
         SubCellInst2_LFInst_5_LFInst_3_n14 ,
         SubCellInst2_LFInst_5_LFInst_3_n13 ,
         SubCellInst2_LFInst_5_LFInst_3_n12 ,
         SubCellInst2_LFInst_5_LFInst_3_n11 ,
         SubCellInst2_LFInst_5_LFInst_2_n22 ,
         SubCellInst2_LFInst_5_LFInst_2_n21 ,
         SubCellInst2_LFInst_5_LFInst_2_n20 ,
         SubCellInst2_LFInst_5_LFInst_2_n19 ,
         SubCellInst2_LFInst_5_LFInst_2_n18 ,
         SubCellInst2_LFInst_5_LFInst_2_n17 ,
         SubCellInst2_LFInst_5_LFInst_2_n16 ,
         SubCellInst2_LFInst_5_LFInst_2_n15 ,
         SubCellInst2_LFInst_5_LFInst_1_n18 ,
         SubCellInst2_LFInst_5_LFInst_1_n17 ,
         SubCellInst2_LFInst_5_LFInst_1_n16 ,
         SubCellInst2_LFInst_5_LFInst_1_n15 ,
         SubCellInst2_LFInst_5_LFInst_1_n14 ,
         SubCellInst2_LFInst_5_LFInst_1_n13 ,
         SubCellInst2_LFInst_5_LFInst_1_n12 ,
         SubCellInst2_LFInst_5_LFInst_1_n11 ,
         SubCellInst2_LFInst_5_LFInst_1_n10 ,
         SubCellInst2_LFInst_5_LFInst_0_n6 ,
         SubCellInst2_LFInst_5_LFInst_0_n5 ,
         SubCellInst2_LFInst_5_LFInst_0_n4 ,
         SubCellInst2_LFInst_6_LFInst_3_n16 ,
         SubCellInst2_LFInst_6_LFInst_3_n15 ,
         SubCellInst2_LFInst_6_LFInst_3_n14 ,
         SubCellInst2_LFInst_6_LFInst_3_n13 ,
         SubCellInst2_LFInst_6_LFInst_3_n12 ,
         SubCellInst2_LFInst_6_LFInst_3_n11 ,
         SubCellInst2_LFInst_6_LFInst_2_n22 ,
         SubCellInst2_LFInst_6_LFInst_2_n21 ,
         SubCellInst2_LFInst_6_LFInst_2_n20 ,
         SubCellInst2_LFInst_6_LFInst_2_n19 ,
         SubCellInst2_LFInst_6_LFInst_2_n18 ,
         SubCellInst2_LFInst_6_LFInst_2_n17 ,
         SubCellInst2_LFInst_6_LFInst_2_n16 ,
         SubCellInst2_LFInst_6_LFInst_2_n15 ,
         SubCellInst2_LFInst_6_LFInst_1_n18 ,
         SubCellInst2_LFInst_6_LFInst_1_n17 ,
         SubCellInst2_LFInst_6_LFInst_1_n16 ,
         SubCellInst2_LFInst_6_LFInst_1_n15 ,
         SubCellInst2_LFInst_6_LFInst_1_n14 ,
         SubCellInst2_LFInst_6_LFInst_1_n13 ,
         SubCellInst2_LFInst_6_LFInst_1_n12 ,
         SubCellInst2_LFInst_6_LFInst_1_n11 ,
         SubCellInst2_LFInst_6_LFInst_1_n10 ,
         SubCellInst2_LFInst_6_LFInst_0_n6 ,
         SubCellInst2_LFInst_6_LFInst_0_n5 ,
         SubCellInst2_LFInst_6_LFInst_0_n4 ,
         SubCellInst2_LFInst_7_LFInst_3_n16 ,
         SubCellInst2_LFInst_7_LFInst_3_n15 ,
         SubCellInst2_LFInst_7_LFInst_3_n14 ,
         SubCellInst2_LFInst_7_LFInst_3_n13 ,
         SubCellInst2_LFInst_7_LFInst_3_n12 ,
         SubCellInst2_LFInst_7_LFInst_3_n11 ,
         SubCellInst2_LFInst_7_LFInst_2_n22 ,
         SubCellInst2_LFInst_7_LFInst_2_n21 ,
         SubCellInst2_LFInst_7_LFInst_2_n20 ,
         SubCellInst2_LFInst_7_LFInst_2_n19 ,
         SubCellInst2_LFInst_7_LFInst_2_n18 ,
         SubCellInst2_LFInst_7_LFInst_2_n17 ,
         SubCellInst2_LFInst_7_LFInst_2_n16 ,
         SubCellInst2_LFInst_7_LFInst_2_n15 ,
         SubCellInst2_LFInst_7_LFInst_1_n18 ,
         SubCellInst2_LFInst_7_LFInst_1_n17 ,
         SubCellInst2_LFInst_7_LFInst_1_n16 ,
         SubCellInst2_LFInst_7_LFInst_1_n15 ,
         SubCellInst2_LFInst_7_LFInst_1_n14 ,
         SubCellInst2_LFInst_7_LFInst_1_n13 ,
         SubCellInst2_LFInst_7_LFInst_1_n12 ,
         SubCellInst2_LFInst_7_LFInst_1_n11 ,
         SubCellInst2_LFInst_7_LFInst_1_n10 ,
         SubCellInst2_LFInst_7_LFInst_0_n6 ,
         SubCellInst2_LFInst_7_LFInst_0_n5 ,
         SubCellInst2_LFInst_7_LFInst_0_n4 ,
         SubCellInst2_LFInst_8_LFInst_3_n16 ,
         SubCellInst2_LFInst_8_LFInst_3_n15 ,
         SubCellInst2_LFInst_8_LFInst_3_n14 ,
         SubCellInst2_LFInst_8_LFInst_3_n13 ,
         SubCellInst2_LFInst_8_LFInst_3_n12 ,
         SubCellInst2_LFInst_8_LFInst_3_n11 ,
         SubCellInst2_LFInst_8_LFInst_2_n22 ,
         SubCellInst2_LFInst_8_LFInst_2_n21 ,
         SubCellInst2_LFInst_8_LFInst_2_n20 ,
         SubCellInst2_LFInst_8_LFInst_2_n19 ,
         SubCellInst2_LFInst_8_LFInst_2_n18 ,
         SubCellInst2_LFInst_8_LFInst_2_n17 ,
         SubCellInst2_LFInst_8_LFInst_2_n16 ,
         SubCellInst2_LFInst_8_LFInst_2_n15 ,
         SubCellInst2_LFInst_8_LFInst_1_n18 ,
         SubCellInst2_LFInst_8_LFInst_1_n17 ,
         SubCellInst2_LFInst_8_LFInst_1_n16 ,
         SubCellInst2_LFInst_8_LFInst_1_n15 ,
         SubCellInst2_LFInst_8_LFInst_1_n14 ,
         SubCellInst2_LFInst_8_LFInst_1_n13 ,
         SubCellInst2_LFInst_8_LFInst_1_n12 ,
         SubCellInst2_LFInst_8_LFInst_1_n11 ,
         SubCellInst2_LFInst_8_LFInst_1_n10 ,
         SubCellInst2_LFInst_8_LFInst_0_n6 ,
         SubCellInst2_LFInst_8_LFInst_0_n5 ,
         SubCellInst2_LFInst_8_LFInst_0_n4 ,
         SubCellInst2_LFInst_9_LFInst_3_n16 ,
         SubCellInst2_LFInst_9_LFInst_3_n15 ,
         SubCellInst2_LFInst_9_LFInst_3_n14 ,
         SubCellInst2_LFInst_9_LFInst_3_n13 ,
         SubCellInst2_LFInst_9_LFInst_3_n12 ,
         SubCellInst2_LFInst_9_LFInst_3_n11 ,
         SubCellInst2_LFInst_9_LFInst_2_n22 ,
         SubCellInst2_LFInst_9_LFInst_2_n21 ,
         SubCellInst2_LFInst_9_LFInst_2_n20 ,
         SubCellInst2_LFInst_9_LFInst_2_n19 ,
         SubCellInst2_LFInst_9_LFInst_2_n18 ,
         SubCellInst2_LFInst_9_LFInst_2_n17 ,
         SubCellInst2_LFInst_9_LFInst_2_n16 ,
         SubCellInst2_LFInst_9_LFInst_2_n15 ,
         SubCellInst2_LFInst_9_LFInst_1_n18 ,
         SubCellInst2_LFInst_9_LFInst_1_n17 ,
         SubCellInst2_LFInst_9_LFInst_1_n16 ,
         SubCellInst2_LFInst_9_LFInst_1_n15 ,
         SubCellInst2_LFInst_9_LFInst_1_n14 ,
         SubCellInst2_LFInst_9_LFInst_1_n13 ,
         SubCellInst2_LFInst_9_LFInst_1_n12 ,
         SubCellInst2_LFInst_9_LFInst_1_n11 ,
         SubCellInst2_LFInst_9_LFInst_1_n10 ,
         SubCellInst2_LFInst_9_LFInst_0_n6 ,
         SubCellInst2_LFInst_9_LFInst_0_n5 ,
         SubCellInst2_LFInst_9_LFInst_0_n4 ,
         SubCellInst2_LFInst_10_LFInst_3_n16 ,
         SubCellInst2_LFInst_10_LFInst_3_n15 ,
         SubCellInst2_LFInst_10_LFInst_3_n14 ,
         SubCellInst2_LFInst_10_LFInst_3_n13 ,
         SubCellInst2_LFInst_10_LFInst_3_n12 ,
         SubCellInst2_LFInst_10_LFInst_3_n11 ,
         SubCellInst2_LFInst_10_LFInst_2_n22 ,
         SubCellInst2_LFInst_10_LFInst_2_n21 ,
         SubCellInst2_LFInst_10_LFInst_2_n20 ,
         SubCellInst2_LFInst_10_LFInst_2_n19 ,
         SubCellInst2_LFInst_10_LFInst_2_n18 ,
         SubCellInst2_LFInst_10_LFInst_2_n17 ,
         SubCellInst2_LFInst_10_LFInst_2_n16 ,
         SubCellInst2_LFInst_10_LFInst_2_n15 ,
         SubCellInst2_LFInst_10_LFInst_1_n18 ,
         SubCellInst2_LFInst_10_LFInst_1_n17 ,
         SubCellInst2_LFInst_10_LFInst_1_n16 ,
         SubCellInst2_LFInst_10_LFInst_1_n15 ,
         SubCellInst2_LFInst_10_LFInst_1_n14 ,
         SubCellInst2_LFInst_10_LFInst_1_n13 ,
         SubCellInst2_LFInst_10_LFInst_1_n12 ,
         SubCellInst2_LFInst_10_LFInst_1_n11 ,
         SubCellInst2_LFInst_10_LFInst_1_n10 ,
         SubCellInst2_LFInst_10_LFInst_0_n6 ,
         SubCellInst2_LFInst_10_LFInst_0_n5 ,
         SubCellInst2_LFInst_10_LFInst_0_n4 ,
         SubCellInst2_LFInst_11_LFInst_3_n16 ,
         SubCellInst2_LFInst_11_LFInst_3_n15 ,
         SubCellInst2_LFInst_11_LFInst_3_n14 ,
         SubCellInst2_LFInst_11_LFInst_3_n13 ,
         SubCellInst2_LFInst_11_LFInst_3_n12 ,
         SubCellInst2_LFInst_11_LFInst_3_n11 ,
         SubCellInst2_LFInst_11_LFInst_2_n22 ,
         SubCellInst2_LFInst_11_LFInst_2_n21 ,
         SubCellInst2_LFInst_11_LFInst_2_n20 ,
         SubCellInst2_LFInst_11_LFInst_2_n19 ,
         SubCellInst2_LFInst_11_LFInst_2_n18 ,
         SubCellInst2_LFInst_11_LFInst_2_n17 ,
         SubCellInst2_LFInst_11_LFInst_2_n16 ,
         SubCellInst2_LFInst_11_LFInst_2_n15 ,
         SubCellInst2_LFInst_11_LFInst_1_n18 ,
         SubCellInst2_LFInst_11_LFInst_1_n17 ,
         SubCellInst2_LFInst_11_LFInst_1_n16 ,
         SubCellInst2_LFInst_11_LFInst_1_n15 ,
         SubCellInst2_LFInst_11_LFInst_1_n14 ,
         SubCellInst2_LFInst_11_LFInst_1_n13 ,
         SubCellInst2_LFInst_11_LFInst_1_n12 ,
         SubCellInst2_LFInst_11_LFInst_1_n11 ,
         SubCellInst2_LFInst_11_LFInst_1_n10 ,
         SubCellInst2_LFInst_11_LFInst_0_n6 ,
         SubCellInst2_LFInst_11_LFInst_0_n5 ,
         SubCellInst2_LFInst_11_LFInst_0_n4 ,
         SubCellInst2_LFInst_12_LFInst_3_n16 ,
         SubCellInst2_LFInst_12_LFInst_3_n15 ,
         SubCellInst2_LFInst_12_LFInst_3_n14 ,
         SubCellInst2_LFInst_12_LFInst_3_n13 ,
         SubCellInst2_LFInst_12_LFInst_3_n12 ,
         SubCellInst2_LFInst_12_LFInst_3_n11 ,
         SubCellInst2_LFInst_12_LFInst_2_n22 ,
         SubCellInst2_LFInst_12_LFInst_2_n21 ,
         SubCellInst2_LFInst_12_LFInst_2_n20 ,
         SubCellInst2_LFInst_12_LFInst_2_n19 ,
         SubCellInst2_LFInst_12_LFInst_2_n18 ,
         SubCellInst2_LFInst_12_LFInst_2_n17 ,
         SubCellInst2_LFInst_12_LFInst_2_n16 ,
         SubCellInst2_LFInst_12_LFInst_2_n15 ,
         SubCellInst2_LFInst_12_LFInst_1_n18 ,
         SubCellInst2_LFInst_12_LFInst_1_n17 ,
         SubCellInst2_LFInst_12_LFInst_1_n16 ,
         SubCellInst2_LFInst_12_LFInst_1_n15 ,
         SubCellInst2_LFInst_12_LFInst_1_n14 ,
         SubCellInst2_LFInst_12_LFInst_1_n13 ,
         SubCellInst2_LFInst_12_LFInst_1_n12 ,
         SubCellInst2_LFInst_12_LFInst_1_n11 ,
         SubCellInst2_LFInst_12_LFInst_1_n10 ,
         SubCellInst2_LFInst_12_LFInst_0_n6 ,
         SubCellInst2_LFInst_12_LFInst_0_n5 ,
         SubCellInst2_LFInst_12_LFInst_0_n4 ,
         SubCellInst2_LFInst_13_LFInst_3_n16 ,
         SubCellInst2_LFInst_13_LFInst_3_n15 ,
         SubCellInst2_LFInst_13_LFInst_3_n14 ,
         SubCellInst2_LFInst_13_LFInst_3_n13 ,
         SubCellInst2_LFInst_13_LFInst_3_n12 ,
         SubCellInst2_LFInst_13_LFInst_3_n11 ,
         SubCellInst2_LFInst_13_LFInst_2_n22 ,
         SubCellInst2_LFInst_13_LFInst_2_n21 ,
         SubCellInst2_LFInst_13_LFInst_2_n20 ,
         SubCellInst2_LFInst_13_LFInst_2_n19 ,
         SubCellInst2_LFInst_13_LFInst_2_n18 ,
         SubCellInst2_LFInst_13_LFInst_2_n17 ,
         SubCellInst2_LFInst_13_LFInst_2_n16 ,
         SubCellInst2_LFInst_13_LFInst_2_n15 ,
         SubCellInst2_LFInst_13_LFInst_1_n18 ,
         SubCellInst2_LFInst_13_LFInst_1_n17 ,
         SubCellInst2_LFInst_13_LFInst_1_n16 ,
         SubCellInst2_LFInst_13_LFInst_1_n15 ,
         SubCellInst2_LFInst_13_LFInst_1_n14 ,
         SubCellInst2_LFInst_13_LFInst_1_n13 ,
         SubCellInst2_LFInst_13_LFInst_1_n12 ,
         SubCellInst2_LFInst_13_LFInst_1_n11 ,
         SubCellInst2_LFInst_13_LFInst_1_n10 ,
         SubCellInst2_LFInst_13_LFInst_0_n6 ,
         SubCellInst2_LFInst_13_LFInst_0_n5 ,
         SubCellInst2_LFInst_13_LFInst_0_n4 ,
         SubCellInst2_LFInst_14_LFInst_3_n16 ,
         SubCellInst2_LFInst_14_LFInst_3_n15 ,
         SubCellInst2_LFInst_14_LFInst_3_n14 ,
         SubCellInst2_LFInst_14_LFInst_3_n13 ,
         SubCellInst2_LFInst_14_LFInst_3_n12 ,
         SubCellInst2_LFInst_14_LFInst_3_n11 ,
         SubCellInst2_LFInst_14_LFInst_2_n22 ,
         SubCellInst2_LFInst_14_LFInst_2_n21 ,
         SubCellInst2_LFInst_14_LFInst_2_n20 ,
         SubCellInst2_LFInst_14_LFInst_2_n19 ,
         SubCellInst2_LFInst_14_LFInst_2_n18 ,
         SubCellInst2_LFInst_14_LFInst_2_n17 ,
         SubCellInst2_LFInst_14_LFInst_2_n16 ,
         SubCellInst2_LFInst_14_LFInst_2_n15 ,
         SubCellInst2_LFInst_14_LFInst_1_n18 ,
         SubCellInst2_LFInst_14_LFInst_1_n17 ,
         SubCellInst2_LFInst_14_LFInst_1_n16 ,
         SubCellInst2_LFInst_14_LFInst_1_n15 ,
         SubCellInst2_LFInst_14_LFInst_1_n14 ,
         SubCellInst2_LFInst_14_LFInst_1_n13 ,
         SubCellInst2_LFInst_14_LFInst_1_n12 ,
         SubCellInst2_LFInst_14_LFInst_1_n11 ,
         SubCellInst2_LFInst_14_LFInst_1_n10 ,
         SubCellInst2_LFInst_14_LFInst_0_n6 ,
         SubCellInst2_LFInst_14_LFInst_0_n5 ,
         SubCellInst2_LFInst_14_LFInst_0_n4 ,
         SubCellInst2_LFInst_15_LFInst_3_n16 ,
         SubCellInst2_LFInst_15_LFInst_3_n15 ,
         SubCellInst2_LFInst_15_LFInst_3_n14 ,
         SubCellInst2_LFInst_15_LFInst_3_n13 ,
         SubCellInst2_LFInst_15_LFInst_3_n12 ,
         SubCellInst2_LFInst_15_LFInst_3_n11 ,
         SubCellInst2_LFInst_15_LFInst_2_n22 ,
         SubCellInst2_LFInst_15_LFInst_2_n21 ,
         SubCellInst2_LFInst_15_LFInst_2_n20 ,
         SubCellInst2_LFInst_15_LFInst_2_n19 ,
         SubCellInst2_LFInst_15_LFInst_2_n18 ,
         SubCellInst2_LFInst_15_LFInst_2_n17 ,
         SubCellInst2_LFInst_15_LFInst_2_n16 ,
         SubCellInst2_LFInst_15_LFInst_2_n15 ,
         SubCellInst2_LFInst_15_LFInst_1_n18 ,
         SubCellInst2_LFInst_15_LFInst_1_n17 ,
         SubCellInst2_LFInst_15_LFInst_1_n16 ,
         SubCellInst2_LFInst_15_LFInst_1_n15 ,
         SubCellInst2_LFInst_15_LFInst_1_n14 ,
         SubCellInst2_LFInst_15_LFInst_1_n13 ,
         SubCellInst2_LFInst_15_LFInst_1_n12 ,
         SubCellInst2_LFInst_15_LFInst_1_n11 ,
         SubCellInst2_LFInst_15_LFInst_1_n10 ,
         SubCellInst2_LFInst_15_LFInst_0_n6 ,
         SubCellInst2_LFInst_15_LFInst_0_n5 ,
         SubCellInst2_LFInst_15_LFInst_0_n4 , MCInst2_MC0_v0_2Inst_0_n2 ,
         MCInst2_MC0_v1_2Inst_0_n2 , MCInst2_MC0_v2_3Inst_0_n4 ,
         MCInst2_MC0_v2_3Inst_0_n3 , MCInst2_MC0_v3_3Inst_0_n2 ,
         MCInst2_MC0_v0_2Inst_1_n2 , MCInst2_MC0_v2_1Inst_1_n2 ,
         MCInst2_MC0_v2_2Inst_1_n4 , MCInst2_MC0_v2_2Inst_1_n3 ,
         MCInst2_MC0_v3_3Inst_1_n2 , MCInst2_MC0_v1_1Inst_2_n2 ,
         MCInst2_MC0_v1_2Inst_2_n2 , MCInst2_MC0_v2_1Inst_2_n2 ,
         MCInst2_MC0_v2_2Inst_2_n2 , MCInst2_MC0_v3_1Inst_2_n2 ,
         MCInst2_MC0_v1_2Inst_3_n4 , MCInst2_MC0_v1_2Inst_3_n3 ,
         MCInst2_MC0_v2_2Inst_3_n2 , MCInst2_MC0_v2_3Inst_3_n2 ,
         MCInst2_MC0_r0Inst_XORInst_0_0_n5 ,
         MCInst2_MC0_r0Inst_XORInst_0_0_n4 ,
         MCInst2_MC0_r0Inst_XORInst_0_1_n5 ,
         MCInst2_MC0_r0Inst_XORInst_0_1_n4 ,
         MCInst2_MC0_r0Inst_XORInst_0_2_n5 ,
         MCInst2_MC0_r0Inst_XORInst_0_2_n4 ,
         MCInst2_MC0_r0Inst_XORInst_0_3_n5 ,
         MCInst2_MC0_r0Inst_XORInst_0_3_n4 ,
         MCInst2_MC0_r1Inst_XORInst_0_0_n5 ,
         MCInst2_MC0_r1Inst_XORInst_0_0_n4 ,
         MCInst2_MC0_r1Inst_XORInst_0_1_n5 ,
         MCInst2_MC0_r1Inst_XORInst_0_1_n4 ,
         MCInst2_MC0_r1Inst_XORInst_0_2_n5 ,
         MCInst2_MC0_r1Inst_XORInst_0_2_n4 ,
         MCInst2_MC0_r1Inst_XORInst_0_3_n5 ,
         MCInst2_MC0_r1Inst_XORInst_0_3_n4 ,
         MCInst2_MC0_r2Inst_XORInst_0_0_n5 ,
         MCInst2_MC0_r2Inst_XORInst_0_0_n4 ,
         MCInst2_MC0_r2Inst_XORInst_0_1_n5 ,
         MCInst2_MC0_r2Inst_XORInst_0_1_n4 ,
         MCInst2_MC0_r2Inst_XORInst_0_2_n5 ,
         MCInst2_MC0_r2Inst_XORInst_0_2_n4 ,
         MCInst2_MC0_r2Inst_XORInst_0_3_n5 ,
         MCInst2_MC0_r2Inst_XORInst_0_3_n4 ,
         MCInst2_MC0_r3Inst_XORInst_0_0_n5 ,
         MCInst2_MC0_r3Inst_XORInst_0_0_n4 ,
         MCInst2_MC0_r3Inst_XORInst_0_1_n5 ,
         MCInst2_MC0_r3Inst_XORInst_0_1_n4 ,
         MCInst2_MC0_r3Inst_XORInst_0_2_n5 ,
         MCInst2_MC0_r3Inst_XORInst_0_2_n4 ,
         MCInst2_MC0_r3Inst_XORInst_0_3_n5 ,
         MCInst2_MC0_r3Inst_XORInst_0_3_n4 , MCInst2_MC1_v0_2Inst_0_n2 ,
         MCInst2_MC1_v1_2Inst_0_n2 , MCInst2_MC1_v2_3Inst_0_n4 ,
         MCInst2_MC1_v2_3Inst_0_n3 , MCInst2_MC1_v3_3Inst_0_n2 ,
         MCInst2_MC1_v0_2Inst_1_n2 , MCInst2_MC1_v2_1Inst_1_n2 ,
         MCInst2_MC1_v2_2Inst_1_n4 , MCInst2_MC1_v2_2Inst_1_n3 ,
         MCInst2_MC1_v3_3Inst_1_n2 , MCInst2_MC1_v1_1Inst_2_n2 ,
         MCInst2_MC1_v1_2Inst_2_n2 , MCInst2_MC1_v2_1Inst_2_n2 ,
         MCInst2_MC1_v2_2Inst_2_n2 , MCInst2_MC1_v3_1Inst_2_n2 ,
         MCInst2_MC1_v1_2Inst_3_n4 , MCInst2_MC1_v1_2Inst_3_n3 ,
         MCInst2_MC1_v2_2Inst_3_n2 , MCInst2_MC1_v2_3Inst_3_n2 ,
         MCInst2_MC1_r0Inst_XORInst_0_0_n5 ,
         MCInst2_MC1_r0Inst_XORInst_0_0_n4 ,
         MCInst2_MC1_r0Inst_XORInst_0_1_n5 ,
         MCInst2_MC1_r0Inst_XORInst_0_1_n4 ,
         MCInst2_MC1_r0Inst_XORInst_0_2_n5 ,
         MCInst2_MC1_r0Inst_XORInst_0_2_n4 ,
         MCInst2_MC1_r0Inst_XORInst_0_3_n5 ,
         MCInst2_MC1_r0Inst_XORInst_0_3_n4 ,
         MCInst2_MC1_r1Inst_XORInst_0_0_n5 ,
         MCInst2_MC1_r1Inst_XORInst_0_0_n4 ,
         MCInst2_MC1_r1Inst_XORInst_0_1_n5 ,
         MCInst2_MC1_r1Inst_XORInst_0_1_n4 ,
         MCInst2_MC1_r1Inst_XORInst_0_2_n5 ,
         MCInst2_MC1_r1Inst_XORInst_0_2_n4 ,
         MCInst2_MC1_r1Inst_XORInst_0_3_n5 ,
         MCInst2_MC1_r1Inst_XORInst_0_3_n4 ,
         MCInst2_MC1_r2Inst_XORInst_0_0_n5 ,
         MCInst2_MC1_r2Inst_XORInst_0_0_n4 ,
         MCInst2_MC1_r2Inst_XORInst_0_1_n5 ,
         MCInst2_MC1_r2Inst_XORInst_0_1_n4 ,
         MCInst2_MC1_r2Inst_XORInst_0_2_n5 ,
         MCInst2_MC1_r2Inst_XORInst_0_2_n4 ,
         MCInst2_MC1_r2Inst_XORInst_0_3_n5 ,
         MCInst2_MC1_r2Inst_XORInst_0_3_n4 ,
         MCInst2_MC1_r3Inst_XORInst_0_0_n5 ,
         MCInst2_MC1_r3Inst_XORInst_0_0_n4 ,
         MCInst2_MC1_r3Inst_XORInst_0_1_n5 ,
         MCInst2_MC1_r3Inst_XORInst_0_1_n4 ,
         MCInst2_MC1_r3Inst_XORInst_0_2_n5 ,
         MCInst2_MC1_r3Inst_XORInst_0_2_n4 ,
         MCInst2_MC1_r3Inst_XORInst_0_3_n5 ,
         MCInst2_MC1_r3Inst_XORInst_0_3_n4 , MCInst2_MC2_v0_2Inst_0_n2 ,
         MCInst2_MC2_v1_2Inst_0_n2 , MCInst2_MC2_v2_3Inst_0_n4 ,
         MCInst2_MC2_v2_3Inst_0_n3 , MCInst2_MC2_v3_3Inst_0_n2 ,
         MCInst2_MC2_v0_2Inst_1_n2 , MCInst2_MC2_v2_1Inst_1_n2 ,
         MCInst2_MC2_v2_2Inst_1_n4 , MCInst2_MC2_v2_2Inst_1_n3 ,
         MCInst2_MC2_v3_3Inst_1_n2 , MCInst2_MC2_v1_1Inst_2_n2 ,
         MCInst2_MC2_v1_2Inst_2_n2 , MCInst2_MC2_v2_1Inst_2_n2 ,
         MCInst2_MC2_v2_2Inst_2_n2 , MCInst2_MC2_v3_1Inst_2_n2 ,
         MCInst2_MC2_v1_2Inst_3_n4 , MCInst2_MC2_v1_2Inst_3_n3 ,
         MCInst2_MC2_v2_2Inst_3_n2 , MCInst2_MC2_v2_3Inst_3_n2 ,
         MCInst2_MC2_r0Inst_XORInst_0_0_n5 ,
         MCInst2_MC2_r0Inst_XORInst_0_0_n4 ,
         MCInst2_MC2_r0Inst_XORInst_0_1_n5 ,
         MCInst2_MC2_r0Inst_XORInst_0_1_n4 ,
         MCInst2_MC2_r0Inst_XORInst_0_2_n5 ,
         MCInst2_MC2_r0Inst_XORInst_0_2_n4 ,
         MCInst2_MC2_r0Inst_XORInst_0_3_n5 ,
         MCInst2_MC2_r0Inst_XORInst_0_3_n4 ,
         MCInst2_MC2_r1Inst_XORInst_0_0_n5 ,
         MCInst2_MC2_r1Inst_XORInst_0_0_n4 ,
         MCInst2_MC2_r1Inst_XORInst_0_1_n5 ,
         MCInst2_MC2_r1Inst_XORInst_0_1_n4 ,
         MCInst2_MC2_r1Inst_XORInst_0_2_n5 ,
         MCInst2_MC2_r1Inst_XORInst_0_2_n4 ,
         MCInst2_MC2_r1Inst_XORInst_0_3_n5 ,
         MCInst2_MC2_r1Inst_XORInst_0_3_n4 ,
         MCInst2_MC2_r2Inst_XORInst_0_0_n5 ,
         MCInst2_MC2_r2Inst_XORInst_0_0_n4 ,
         MCInst2_MC2_r2Inst_XORInst_0_1_n5 ,
         MCInst2_MC2_r2Inst_XORInst_0_1_n4 ,
         MCInst2_MC2_r2Inst_XORInst_0_2_n5 ,
         MCInst2_MC2_r2Inst_XORInst_0_2_n4 ,
         MCInst2_MC2_r2Inst_XORInst_0_3_n5 ,
         MCInst2_MC2_r2Inst_XORInst_0_3_n4 ,
         MCInst2_MC2_r3Inst_XORInst_0_0_n5 ,
         MCInst2_MC2_r3Inst_XORInst_0_0_n4 ,
         MCInst2_MC2_r3Inst_XORInst_0_1_n5 ,
         MCInst2_MC2_r3Inst_XORInst_0_1_n4 ,
         MCInst2_MC2_r3Inst_XORInst_0_2_n5 ,
         MCInst2_MC2_r3Inst_XORInst_0_2_n4 ,
         MCInst2_MC2_r3Inst_XORInst_0_3_n5 ,
         MCInst2_MC2_r3Inst_XORInst_0_3_n4 , MCInst2_MC3_v0_2Inst_0_n2 ,
         MCInst2_MC3_v1_2Inst_0_n2 , MCInst2_MC3_v2_3Inst_0_n4 ,
         MCInst2_MC3_v2_3Inst_0_n3 , MCInst2_MC3_v3_3Inst_0_n2 ,
         MCInst2_MC3_v0_2Inst_1_n2 , MCInst2_MC3_v2_1Inst_1_n2 ,
         MCInst2_MC3_v2_2Inst_1_n4 , MCInst2_MC3_v2_2Inst_1_n3 ,
         MCInst2_MC3_v3_3Inst_1_n2 , MCInst2_MC3_v1_1Inst_2_n2 ,
         MCInst2_MC3_v1_2Inst_2_n2 , MCInst2_MC3_v2_1Inst_2_n2 ,
         MCInst2_MC3_v2_2Inst_2_n2 , MCInst2_MC3_v3_1Inst_2_n2 ,
         MCInst2_MC3_v1_2Inst_3_n4 , MCInst2_MC3_v1_2Inst_3_n3 ,
         MCInst2_MC3_v2_2Inst_3_n2 , MCInst2_MC3_v2_3Inst_3_n2 ,
         MCInst2_MC3_r0Inst_XORInst_0_0_n5 ,
         MCInst2_MC3_r0Inst_XORInst_0_0_n4 ,
         MCInst2_MC3_r0Inst_XORInst_0_1_n5 ,
         MCInst2_MC3_r0Inst_XORInst_0_1_n4 ,
         MCInst2_MC3_r0Inst_XORInst_0_2_n5 ,
         MCInst2_MC3_r0Inst_XORInst_0_2_n4 ,
         MCInst2_MC3_r0Inst_XORInst_0_3_n5 ,
         MCInst2_MC3_r0Inst_XORInst_0_3_n4 ,
         MCInst2_MC3_r1Inst_XORInst_0_0_n5 ,
         MCInst2_MC3_r1Inst_XORInst_0_0_n4 ,
         MCInst2_MC3_r1Inst_XORInst_0_1_n5 ,
         MCInst2_MC3_r1Inst_XORInst_0_1_n4 ,
         MCInst2_MC3_r1Inst_XORInst_0_2_n5 ,
         MCInst2_MC3_r1Inst_XORInst_0_2_n4 ,
         MCInst2_MC3_r1Inst_XORInst_0_3_n5 ,
         MCInst2_MC3_r1Inst_XORInst_0_3_n4 ,
         MCInst2_MC3_r2Inst_XORInst_0_0_n5 ,
         MCInst2_MC3_r2Inst_XORInst_0_0_n4 ,
         MCInst2_MC3_r2Inst_XORInst_0_1_n5 ,
         MCInst2_MC3_r2Inst_XORInst_0_1_n4 ,
         MCInst2_MC3_r2Inst_XORInst_0_2_n5 ,
         MCInst2_MC3_r2Inst_XORInst_0_2_n4 ,
         MCInst2_MC3_r2Inst_XORInst_0_3_n5 ,
         MCInst2_MC3_r2Inst_XORInst_0_3_n4 ,
         MCInst2_MC3_r3Inst_XORInst_0_0_n5 ,
         MCInst2_MC3_r3Inst_XORInst_0_0_n4 ,
         MCInst2_MC3_r3Inst_XORInst_0_1_n5 ,
         MCInst2_MC3_r3Inst_XORInst_0_1_n4 ,
         MCInst2_MC3_r3Inst_XORInst_0_2_n5 ,
         MCInst2_MC3_r3Inst_XORInst_0_2_n4 ,
         MCInst2_MC3_r3Inst_XORInst_0_3_n5 ,
         MCInst2_MC3_r3Inst_XORInst_0_3_n4 ;
  wire   [63:0] AddRoundKeyOutput;
  wire   [63:0] ShiftRowsOutput;
  wire   [63:0] Feedback;
  wire   [63:0] SubCellInput;
  wire   [63:0] ShiftRowsOutput2;
  wire   [3:0] MCInst1_MC0_v3_3 ;
  wire   [3:0] MCInst1_MC0_v3_2 ;
  wire   [3:0] MCInst1_MC0_v3_1 ;
  wire   [3:0] MCInst1_MC0_v3_0 ;
  wire   [3:0] MCInst1_MC0_v2_3 ;
  wire   [3:0] MCInst1_MC0_v2_2 ;
  wire   [3:0] MCInst1_MC0_v2_1 ;
  wire   [3:0] MCInst1_MC0_v2_0 ;
  wire   [3:0] MCInst1_MC0_v1_3 ;
  wire   [3:0] MCInst1_MC0_v1_2 ;
  wire   [3:0] MCInst1_MC0_v1_1 ;
  wire   [3:0] MCInst1_MC0_v0_3 ;
  wire   [3:0] MCInst1_MC0_v0_2 ;
  wire   [3:0] MCInst1_MC0_v0_1 ;
  wire   [3:0] MCInst1_MC0_v0_0 ;
  wire   [3:0] MCInst1_MC1_v3_3 ;
  wire   [3:0] MCInst1_MC1_v3_2 ;
  wire   [3:0] MCInst1_MC1_v3_1 ;
  wire   [3:0] MCInst1_MC1_v3_0 ;
  wire   [3:0] MCInst1_MC1_v2_3 ;
  wire   [3:0] MCInst1_MC1_v2_2 ;
  wire   [3:0] MCInst1_MC1_v2_1 ;
  wire   [3:0] MCInst1_MC1_v2_0 ;
  wire   [3:0] MCInst1_MC1_v1_3 ;
  wire   [3:0] MCInst1_MC1_v1_2 ;
  wire   [3:0] MCInst1_MC1_v1_1 ;
  wire   [3:0] MCInst1_MC1_v0_3 ;
  wire   [3:0] MCInst1_MC1_v0_2 ;
  wire   [3:0] MCInst1_MC1_v0_1 ;
  wire   [3:0] MCInst1_MC1_v0_0 ;
  wire   [3:0] MCInst1_MC2_v3_3 ;
  wire   [3:0] MCInst1_MC2_v3_2 ;
  wire   [3:0] MCInst1_MC2_v3_1 ;
  wire   [3:0] MCInst1_MC2_v3_0 ;
  wire   [3:0] MCInst1_MC2_v2_3 ;
  wire   [3:0] MCInst1_MC2_v2_2 ;
  wire   [3:0] MCInst1_MC2_v2_1 ;
  wire   [3:0] MCInst1_MC2_v2_0 ;
  wire   [3:0] MCInst1_MC2_v1_3 ;
  wire   [3:0] MCInst1_MC2_v1_2 ;
  wire   [3:0] MCInst1_MC2_v1_1 ;
  wire   [3:0] MCInst1_MC2_v0_3 ;
  wire   [3:0] MCInst1_MC2_v0_2 ;
  wire   [3:0] MCInst1_MC2_v0_1 ;
  wire   [3:0] MCInst1_MC2_v0_0 ;
  wire   [3:0] MCInst1_MC3_v3_3 ;
  wire   [3:0] MCInst1_MC3_v3_2 ;
  wire   [3:0] MCInst1_MC3_v3_1 ;
  wire   [3:0] MCInst1_MC3_v3_0 ;
  wire   [3:0] MCInst1_MC3_v2_3 ;
  wire   [3:0] MCInst1_MC3_v2_2 ;
  wire   [3:0] MCInst1_MC3_v2_1 ;
  wire   [3:0] MCInst1_MC3_v2_0 ;
  wire   [3:0] MCInst1_MC3_v1_3 ;
  wire   [3:0] MCInst1_MC3_v1_2 ;
  wire   [3:0] MCInst1_MC3_v1_1 ;
  wire   [3:0] MCInst1_MC3_v0_3 ;
  wire   [3:0] MCInst1_MC3_v0_2 ;
  wire   [3:0] MCInst1_MC3_v0_1 ;
  wire   [3:0] MCInst1_MC3_v0_0 ;
  wire   [3:0] MCInst2_MC0_v3_3 ;
  wire   [3:0] MCInst2_MC0_v3_2 ;
  wire   [3:0] MCInst2_MC0_v3_1 ;
  wire   [3:0] MCInst2_MC0_v3_0 ;
  wire   [3:0] MCInst2_MC0_v2_3 ;
  wire   [3:0] MCInst2_MC0_v2_2 ;
  wire   [3:0] MCInst2_MC0_v2_1 ;
  wire   [3:0] MCInst2_MC0_v2_0 ;
  wire   [3:0] MCInst2_MC0_v1_3 ;
  wire   [3:0] MCInst2_MC0_v1_2 ;
  wire   [3:0] MCInst2_MC0_v1_1 ;
  wire   [3:0] MCInst2_MC0_v0_3 ;
  wire   [3:0] MCInst2_MC0_v0_2 ;
  wire   [3:0] MCInst2_MC0_v0_1 ;
  wire   [3:0] MCInst2_MC0_v0_0 ;
  wire   [3:0] MCInst2_MC1_v3_3 ;
  wire   [3:0] MCInst2_MC1_v3_2 ;
  wire   [3:0] MCInst2_MC1_v3_1 ;
  wire   [3:0] MCInst2_MC1_v3_0 ;
  wire   [3:0] MCInst2_MC1_v2_3 ;
  wire   [3:0] MCInst2_MC1_v2_2 ;
  wire   [3:0] MCInst2_MC1_v2_1 ;
  wire   [3:0] MCInst2_MC1_v2_0 ;
  wire   [3:0] MCInst2_MC1_v1_3 ;
  wire   [3:0] MCInst2_MC1_v1_2 ;
  wire   [3:0] MCInst2_MC1_v1_1 ;
  wire   [3:0] MCInst2_MC1_v0_3 ;
  wire   [3:0] MCInst2_MC1_v0_2 ;
  wire   [3:0] MCInst2_MC1_v0_1 ;
  wire   [3:0] MCInst2_MC1_v0_0 ;
  wire   [3:0] MCInst2_MC2_v3_3 ;
  wire   [3:0] MCInst2_MC2_v3_2 ;
  wire   [3:0] MCInst2_MC2_v3_1 ;
  wire   [3:0] MCInst2_MC2_v3_0 ;
  wire   [3:0] MCInst2_MC2_v2_3 ;
  wire   [3:0] MCInst2_MC2_v2_2 ;
  wire   [3:0] MCInst2_MC2_v2_1 ;
  wire   [3:0] MCInst2_MC2_v2_0 ;
  wire   [3:0] MCInst2_MC2_v1_3 ;
  wire   [3:0] MCInst2_MC2_v1_2 ;
  wire   [3:0] MCInst2_MC2_v1_1 ;
  wire   [3:0] MCInst2_MC2_v0_3 ;
  wire   [3:0] MCInst2_MC2_v0_2 ;
  wire   [3:0] MCInst2_MC2_v0_1 ;
  wire   [3:0] MCInst2_MC2_v0_0 ;
  wire   [3:0] MCInst2_MC3_v3_3 ;
  wire   [3:0] MCInst2_MC3_v3_2 ;
  wire   [3:0] MCInst2_MC3_v3_1 ;
  wire   [3:0] MCInst2_MC3_v3_0 ;
  wire   [3:0] MCInst2_MC3_v2_3 ;
  wire   [3:0] MCInst2_MC3_v2_2 ;
  wire   [3:0] MCInst2_MC3_v2_1 ;
  wire   [3:0] MCInst2_MC3_v2_0 ;
  wire   [3:0] MCInst2_MC3_v1_3 ;
  wire   [3:0] MCInst2_MC3_v1_2 ;
  wire   [3:0] MCInst2_MC3_v1_1 ;
  wire   [3:0] MCInst2_MC3_v0_3 ;
  wire   [3:0] MCInst2_MC3_v0_2 ;
  wire   [3:0] MCInst2_MC3_v0_1 ;
  wire   [3:0] MCInst2_MC3_v0_0 ;

  XOR2_X1 AddKeyXOR_XORInst_0_0_U1  ( .A(Plaintext[0]), .B(Key[0]), .Z(
        AddRoundKeyOutput[0]) );
  XOR2_X1 AddKeyXOR_XORInst_0_1_U1  ( .A(Plaintext[1]), .B(Key[1]), .Z(
        AddRoundKeyOutput[1]) );
  XOR2_X1 AddKeyXOR_XORInst_0_2_U1  ( .A(Plaintext[2]), .B(Key[2]), .Z(
        AddRoundKeyOutput[2]) );
  XOR2_X1 AddKeyXOR_XORInst_0_3_U1  ( .A(Plaintext[3]), .B(Key[3]), .Z(
        AddRoundKeyOutput[3]) );
  XOR2_X1 AddKeyXOR_XORInst_1_0_U1  ( .A(Plaintext[4]), .B(Key[4]), .Z(
        AddRoundKeyOutput[4]) );
  XOR2_X1 AddKeyXOR_XORInst_1_1_U1  ( .A(Plaintext[5]), .B(Key[5]), .Z(
        AddRoundKeyOutput[5]) );
  XOR2_X1 AddKeyXOR_XORInst_1_2_U1  ( .A(Plaintext[6]), .B(Key[6]), .Z(
        AddRoundKeyOutput[6]) );
  XOR2_X1 AddKeyXOR_XORInst_1_3_U1  ( .A(Plaintext[7]), .B(Key[7]), .Z(
        AddRoundKeyOutput[7]) );
  XOR2_X1 AddKeyXOR_XORInst_2_0_U1  ( .A(Plaintext[8]), .B(Key[8]), .Z(
        AddRoundKeyOutput[8]) );
  XOR2_X1 AddKeyXOR_XORInst_2_1_U1  ( .A(Plaintext[9]), .B(Key[9]), .Z(
        AddRoundKeyOutput[9]) );
  XOR2_X1 AddKeyXOR_XORInst_2_2_U1  ( .A(Plaintext[10]), .B(Key[10]), .Z(
        AddRoundKeyOutput[10]) );
  XOR2_X1 AddKeyXOR_XORInst_2_3_U1  ( .A(Plaintext[11]), .B(Key[11]), .Z(
        AddRoundKeyOutput[11]) );
  XOR2_X1 AddKeyXOR_XORInst_3_0_U1  ( .A(Plaintext[12]), .B(Key[12]), .Z(
        AddRoundKeyOutput[12]) );
  XOR2_X1 AddKeyXOR_XORInst_3_1_U1  ( .A(Plaintext[13]), .B(Key[13]), .Z(
        AddRoundKeyOutput[13]) );
  XOR2_X1 AddKeyXOR_XORInst_3_2_U1  ( .A(Plaintext[14]), .B(Key[14]), .Z(
        AddRoundKeyOutput[14]) );
  XOR2_X1 AddKeyXOR_XORInst_3_3_U1  ( .A(Plaintext[15]), .B(Key[15]), .Z(
        AddRoundKeyOutput[15]) );
  XOR2_X1 AddKeyXOR_XORInst_4_0_U1  ( .A(Plaintext[16]), .B(Key[16]), .Z(
        AddRoundKeyOutput[16]) );
  XOR2_X1 AddKeyXOR_XORInst_4_1_U1  ( .A(Plaintext[17]), .B(Key[17]), .Z(
        AddRoundKeyOutput[17]) );
  XOR2_X1 AddKeyXOR_XORInst_4_2_U1  ( .A(Plaintext[18]), .B(Key[18]), .Z(
        AddRoundKeyOutput[18]) );
  XOR2_X1 AddKeyXOR_XORInst_4_3_U1  ( .A(Plaintext[19]), .B(Key[19]), .Z(
        AddRoundKeyOutput[19]) );
  XOR2_X1 AddKeyXOR_XORInst_5_0_U1  ( .A(Plaintext[20]), .B(Key[20]), .Z(
        AddRoundKeyOutput[20]) );
  XOR2_X1 AddKeyXOR_XORInst_5_1_U1  ( .A(Plaintext[21]), .B(Key[21]), .Z(
        AddRoundKeyOutput[21]) );
  XOR2_X1 AddKeyXOR_XORInst_5_2_U1  ( .A(Plaintext[22]), .B(Key[22]), .Z(
        AddRoundKeyOutput[22]) );
  XOR2_X1 AddKeyXOR_XORInst_5_3_U1  ( .A(Plaintext[23]), .B(Key[23]), .Z(
        AddRoundKeyOutput[23]) );
  XOR2_X1 AddKeyXOR_XORInst_6_0_U1  ( .A(Plaintext[24]), .B(Key[24]), .Z(
        AddRoundKeyOutput[24]) );
  XOR2_X1 AddKeyXOR_XORInst_6_1_U1  ( .A(Plaintext[25]), .B(Key[25]), .Z(
        AddRoundKeyOutput[25]) );
  XOR2_X1 AddKeyXOR_XORInst_6_2_U1  ( .A(Plaintext[26]), .B(Key[26]), .Z(
        AddRoundKeyOutput[26]) );
  XOR2_X1 AddKeyXOR_XORInst_6_3_U1  ( .A(Plaintext[27]), .B(Key[27]), .Z(
        AddRoundKeyOutput[27]) );
  XOR2_X1 AddKeyXOR_XORInst_7_0_U1  ( .A(Plaintext[28]), .B(Key[28]), .Z(
        AddRoundKeyOutput[28]) );
  XOR2_X1 AddKeyXOR_XORInst_7_1_U1  ( .A(Plaintext[29]), .B(Key[29]), .Z(
        AddRoundKeyOutput[29]) );
  XOR2_X1 AddKeyXOR_XORInst_7_2_U1  ( .A(Plaintext[30]), .B(Key[30]), .Z(
        AddRoundKeyOutput[30]) );
  XOR2_X1 AddKeyXOR_XORInst_7_3_U1  ( .A(Plaintext[31]), .B(Key[31]), .Z(
        AddRoundKeyOutput[31]) );
  XOR2_X1 AddKeyXOR_XORInst_8_0_U1  ( .A(Plaintext[32]), .B(Key[32]), .Z(
        AddRoundKeyOutput[32]) );
  XOR2_X1 AddKeyXOR_XORInst_8_1_U1  ( .A(Plaintext[33]), .B(Key[33]), .Z(
        AddRoundKeyOutput[33]) );
  XOR2_X1 AddKeyXOR_XORInst_8_2_U1  ( .A(Plaintext[34]), .B(Key[34]), .Z(
        AddRoundKeyOutput[34]) );
  XOR2_X1 AddKeyXOR_XORInst_8_3_U1  ( .A(Plaintext[35]), .B(Key[35]), .Z(
        AddRoundKeyOutput[35]) );
  XOR2_X1 AddKeyXOR_XORInst_9_0_U1  ( .A(Plaintext[36]), .B(Key[36]), .Z(
        AddRoundKeyOutput[36]) );
  XOR2_X1 AddKeyXOR_XORInst_9_1_U1  ( .A(Plaintext[37]), .B(Key[37]), .Z(
        AddRoundKeyOutput[37]) );
  XOR2_X1 AddKeyXOR_XORInst_9_2_U1  ( .A(Plaintext[38]), .B(Key[38]), .Z(
        AddRoundKeyOutput[38]) );
  XOR2_X1 AddKeyXOR_XORInst_9_3_U1  ( .A(Plaintext[39]), .B(Key[39]), .Z(
        AddRoundKeyOutput[39]) );
  XOR2_X1 AddKeyXOR_XORInst_10_0_U1  ( .A(Plaintext[40]), .B(Key[40]), .Z(
        AddRoundKeyOutput[40]) );
  XOR2_X1 AddKeyXOR_XORInst_10_1_U1  ( .A(Plaintext[41]), .B(Key[41]), .Z(
        AddRoundKeyOutput[41]) );
  XOR2_X1 AddKeyXOR_XORInst_10_2_U1  ( .A(Plaintext[42]), .B(Key[42]), .Z(
        AddRoundKeyOutput[42]) );
  XOR2_X1 AddKeyXOR_XORInst_10_3_U1  ( .A(Plaintext[43]), .B(Key[43]), .Z(
        AddRoundKeyOutput[43]) );
  XOR2_X1 AddKeyXOR_XORInst_11_0_U1  ( .A(Plaintext[44]), .B(Key[44]), .Z(
        AddRoundKeyOutput[44]) );
  XOR2_X1 AddKeyXOR_XORInst_11_1_U1  ( .A(Plaintext[45]), .B(Key[45]), .Z(
        AddRoundKeyOutput[45]) );
  XOR2_X1 AddKeyXOR_XORInst_11_2_U1  ( .A(Plaintext[46]), .B(Key[46]), .Z(
        AddRoundKeyOutput[46]) );
  XOR2_X1 AddKeyXOR_XORInst_11_3_U1  ( .A(Plaintext[47]), .B(Key[47]), .Z(
        AddRoundKeyOutput[47]) );
  XOR2_X1 AddKeyXOR_XORInst_12_0_U1  ( .A(Plaintext[48]), .B(Key[48]), .Z(
        AddRoundKeyOutput[48]) );
  XOR2_X1 AddKeyXOR_XORInst_12_1_U1  ( .A(Plaintext[49]), .B(Key[49]), .Z(
        AddRoundKeyOutput[49]) );
  XOR2_X1 AddKeyXOR_XORInst_12_2_U1  ( .A(Plaintext[50]), .B(Key[50]), .Z(
        AddRoundKeyOutput[50]) );
  XOR2_X1 AddKeyXOR_XORInst_12_3_U1  ( .A(Plaintext[51]), .B(Key[51]), .Z(
        AddRoundKeyOutput[51]) );
  XOR2_X1 AddKeyXOR_XORInst_13_0_U1  ( .A(Plaintext[52]), .B(Key[52]), .Z(
        AddRoundKeyOutput[52]) );
  XOR2_X1 AddKeyXOR_XORInst_13_1_U1  ( .A(Plaintext[53]), .B(Key[53]), .Z(
        AddRoundKeyOutput[53]) );
  XOR2_X1 AddKeyXOR_XORInst_13_2_U1  ( .A(Plaintext[54]), .B(Key[54]), .Z(
        AddRoundKeyOutput[54]) );
  XOR2_X1 AddKeyXOR_XORInst_13_3_U1  ( .A(Plaintext[55]), .B(Key[55]), .Z(
        AddRoundKeyOutput[55]) );
  XOR2_X1 AddKeyXOR_XORInst_14_0_U1  ( .A(Plaintext[56]), .B(Key[56]), .Z(
        AddRoundKeyOutput[56]) );
  XOR2_X1 AddKeyXOR_XORInst_14_1_U1  ( .A(Plaintext[57]), .B(Key[57]), .Z(
        AddRoundKeyOutput[57]) );
  XOR2_X1 AddKeyXOR_XORInst_14_2_U1  ( .A(Plaintext[58]), .B(Key[58]), .Z(
        AddRoundKeyOutput[58]) );
  XOR2_X1 AddKeyXOR_XORInst_14_3_U1  ( .A(Plaintext[59]), .B(Key[59]), .Z(
        AddRoundKeyOutput[59]) );
  XOR2_X1 AddKeyXOR_XORInst_15_0_U1  ( .A(Plaintext[60]), .B(Key[60]), .Z(
        AddRoundKeyOutput[60]) );
  XOR2_X1 AddKeyXOR_XORInst_15_1_U1  ( .A(Plaintext[61]), .B(Key[61]), .Z(
        AddRoundKeyOutput[61]) );
  XOR2_X1 AddKeyXOR_XORInst_15_2_U1  ( .A(Plaintext[62]), .B(Key[62]), .Z(
        AddRoundKeyOutput[62]) );
  XOR2_X1 AddKeyXOR_XORInst_15_3_U1  ( .A(Plaintext[63]), .B(Key[63]), .Z(
        AddRoundKeyOutput[63]) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_3_U9  ( .A1(
        SubCellInst_LFInst_0_LFInst_3_n16 ), .A2(
        SubCellInst_LFInst_0_LFInst_3_n15 ), .ZN(MCInst1_MC0_v3_2 [2]) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_3_U8  ( .A1(AddRoundKeyOutput[1]), 
        .A2(SubCellInst_LFInst_0_LFInst_3_n14 ), .ZN(
        SubCellInst_LFInst_0_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst_LFInst_0_LFInst_3_U7  ( .A(AddRoundKeyOutput[3]), .B(
        AddRoundKeyOutput[2]), .Z(SubCellInst_LFInst_0_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_3_U6  ( .A1(
        SubCellInst_LFInst_0_LFInst_3_n13 ), .A2(
        SubCellInst_LFInst_0_LFInst_3_n12 ), .ZN(
        SubCellInst_LFInst_0_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_3_U5  ( .A1(AddRoundKeyOutput[0]), 
        .A2(AddRoundKeyOutput[2]), .ZN(SubCellInst_LFInst_0_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst_LFInst_0_LFInst_3_U4  ( .A(AddRoundKeyOutput[0]), .B(
        SubCellInst_LFInst_0_LFInst_3_n11 ), .ZN(
        SubCellInst_LFInst_0_LFInst_3_n13 ) );
  OR2_X1 SubCellInst_LFInst_0_LFInst_3_U3  ( .A1(AddRoundKeyOutput[3]), .A2(
        AddRoundKeyOutput[1]), .ZN(SubCellInst_LFInst_0_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_2_U11  ( .A1(
        SubCellInst_LFInst_0_LFInst_2_n22 ), .A2(
        SubCellInst_LFInst_0_LFInst_2_n21 ), .ZN(MCInst1_MC0_v3_0 [3]) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_2_U10  ( .A1(AddRoundKeyOutput[2]), 
        .A2(SubCellInst_LFInst_0_LFInst_2_n20 ), .ZN(
        SubCellInst_LFInst_0_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst_LFInst_0_LFInst_2_U9  ( .A1(AddRoundKeyOutput[1]), .A2(
        SubCellInst_LFInst_0_LFInst_2_n19 ), .ZN(
        SubCellInst_LFInst_0_LFInst_2_n20 ) );
  INV_X1 SubCellInst_LFInst_0_LFInst_2_U8  ( .A(AddRoundKeyOutput[3]), .ZN(
        SubCellInst_LFInst_0_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_2_U7  ( .A1(
        SubCellInst_LFInst_0_LFInst_2_n18 ), .A2(
        SubCellInst_LFInst_0_LFInst_2_n17 ), .ZN(
        SubCellInst_LFInst_0_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst_LFInst_0_LFInst_2_U6  ( .A(
        SubCellInst_LFInst_0_LFInst_2_n16 ), .B(AddRoundKeyOutput[2]), .Z(
        SubCellInst_LFInst_0_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_2_U5  ( .A1(AddRoundKeyOutput[0]), 
        .A2(AddRoundKeyOutput[1]), .ZN(SubCellInst_LFInst_0_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_2_U4  ( .A1(
        SubCellInst_LFInst_0_LFInst_2_n15 ), .A2(AddRoundKeyOutput[3]), .ZN(
        SubCellInst_LFInst_0_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst_LFInst_0_LFInst_2_U3  ( .A(AddRoundKeyOutput[0]), .B(
        AddRoundKeyOutput[1]), .ZN(SubCellInst_LFInst_0_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_1_U12  ( .A1(
        SubCellInst_LFInst_0_LFInst_1_n18 ), .A2(
        SubCellInst_LFInst_0_LFInst_1_n17 ), .ZN(MCInst1_MC0_v3_0 [2]) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_1_U11  ( .A1(AddRoundKeyOutput[1]), 
        .A2(SubCellInst_LFInst_0_LFInst_1_n16 ), .ZN(
        SubCellInst_LFInst_0_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst_LFInst_0_LFInst_1_U10  ( .A1(AddRoundKeyOutput[3]), 
        .A2(SubCellInst_LFInst_0_LFInst_1_n15 ), .ZN(
        SubCellInst_LFInst_0_LFInst_1_n16 ) );
  AND2_X1 SubCellInst_LFInst_0_LFInst_1_U9  ( .A1(AddRoundKeyOutput[0]), .A2(
        AddRoundKeyOutput[2]), .ZN(SubCellInst_LFInst_0_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_1_U8  ( .A1(AddRoundKeyOutput[3]), 
        .A2(SubCellInst_LFInst_0_LFInst_1_n14 ), .ZN(
        SubCellInst_LFInst_0_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_1_U7  ( .A1(
        SubCellInst_LFInst_0_LFInst_1_n13 ), .A2(
        SubCellInst_LFInst_0_LFInst_1_n12 ), .ZN(
        SubCellInst_LFInst_0_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_1_U6  ( .A1(AddRoundKeyOutput[0]), 
        .A2(AddRoundKeyOutput[2]), .ZN(SubCellInst_LFInst_0_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_1_U5  ( .A1(
        SubCellInst_LFInst_0_LFInst_1_n11 ), .A2(
        SubCellInst_LFInst_0_LFInst_1_n10 ), .ZN(
        SubCellInst_LFInst_0_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_1_U4  ( .A1(AddRoundKeyOutput[0]), 
        .A2(AddRoundKeyOutput[1]), .ZN(SubCellInst_LFInst_0_LFInst_1_n10 ) );
  INV_X1 SubCellInst_LFInst_0_LFInst_1_U3  ( .A(AddRoundKeyOutput[2]), .ZN(
        SubCellInst_LFInst_0_LFInst_1_n11 ) );
  XNOR2_X1 SubCellInst_LFInst_0_LFInst_0_U6  ( .A(
        SubCellInst_LFInst_0_LFInst_0_n6 ), .B(
        SubCellInst_LFInst_0_LFInst_0_n5 ), .ZN(MCInst1_MC0_v3_2 [3]) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_0_U5  ( .A1(AddRoundKeyOutput[2]), 
        .A2(SubCellInst_LFInst_0_LFInst_0_n4 ), .ZN(
        SubCellInst_LFInst_0_LFInst_0_n5 ) );
  INV_X1 SubCellInst_LFInst_0_LFInst_0_U4  ( .A(AddRoundKeyOutput[1]), .ZN(
        SubCellInst_LFInst_0_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst_LFInst_0_LFInst_0_U3  ( .A(AddRoundKeyOutput[0]), .B(
        AddRoundKeyOutput[3]), .Z(SubCellInst_LFInst_0_LFInst_0_n6 ) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_3_U9  ( .A1(
        SubCellInst_LFInst_1_LFInst_3_n16 ), .A2(
        SubCellInst_LFInst_1_LFInst_3_n15 ), .ZN(MCInst1_MC3_v3_2 [2]) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_3_U8  ( .A1(AddRoundKeyOutput[5]), 
        .A2(SubCellInst_LFInst_1_LFInst_3_n14 ), .ZN(
        SubCellInst_LFInst_1_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst_LFInst_1_LFInst_3_U7  ( .A(AddRoundKeyOutput[7]), .B(
        AddRoundKeyOutput[6]), .Z(SubCellInst_LFInst_1_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_3_U6  ( .A1(
        SubCellInst_LFInst_1_LFInst_3_n13 ), .A2(
        SubCellInst_LFInst_1_LFInst_3_n12 ), .ZN(
        SubCellInst_LFInst_1_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_3_U5  ( .A1(AddRoundKeyOutput[4]), 
        .A2(AddRoundKeyOutput[6]), .ZN(SubCellInst_LFInst_1_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst_LFInst_1_LFInst_3_U4  ( .A(AddRoundKeyOutput[4]), .B(
        SubCellInst_LFInst_1_LFInst_3_n11 ), .ZN(
        SubCellInst_LFInst_1_LFInst_3_n13 ) );
  OR2_X1 SubCellInst_LFInst_1_LFInst_3_U3  ( .A1(AddRoundKeyOutput[7]), .A2(
        AddRoundKeyOutput[5]), .ZN(SubCellInst_LFInst_1_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_2_U11  ( .A1(
        SubCellInst_LFInst_1_LFInst_2_n22 ), .A2(
        SubCellInst_LFInst_1_LFInst_2_n21 ), .ZN(MCInst1_MC3_v3_0 [3]) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_2_U10  ( .A1(AddRoundKeyOutput[6]), 
        .A2(SubCellInst_LFInst_1_LFInst_2_n20 ), .ZN(
        SubCellInst_LFInst_1_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst_LFInst_1_LFInst_2_U9  ( .A1(AddRoundKeyOutput[5]), .A2(
        SubCellInst_LFInst_1_LFInst_2_n19 ), .ZN(
        SubCellInst_LFInst_1_LFInst_2_n20 ) );
  INV_X1 SubCellInst_LFInst_1_LFInst_2_U8  ( .A(AddRoundKeyOutput[7]), .ZN(
        SubCellInst_LFInst_1_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_2_U7  ( .A1(
        SubCellInst_LFInst_1_LFInst_2_n18 ), .A2(
        SubCellInst_LFInst_1_LFInst_2_n17 ), .ZN(
        SubCellInst_LFInst_1_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst_LFInst_1_LFInst_2_U6  ( .A(
        SubCellInst_LFInst_1_LFInst_2_n16 ), .B(AddRoundKeyOutput[6]), .Z(
        SubCellInst_LFInst_1_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_2_U5  ( .A1(AddRoundKeyOutput[4]), 
        .A2(AddRoundKeyOutput[5]), .ZN(SubCellInst_LFInst_1_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_2_U4  ( .A1(
        SubCellInst_LFInst_1_LFInst_2_n15 ), .A2(AddRoundKeyOutput[7]), .ZN(
        SubCellInst_LFInst_1_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst_LFInst_1_LFInst_2_U3  ( .A(AddRoundKeyOutput[4]), .B(
        AddRoundKeyOutput[5]), .ZN(SubCellInst_LFInst_1_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_1_U12  ( .A1(
        SubCellInst_LFInst_1_LFInst_1_n18 ), .A2(
        SubCellInst_LFInst_1_LFInst_1_n17 ), .ZN(MCInst1_MC3_v3_0 [2]) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_1_U11  ( .A1(AddRoundKeyOutput[5]), 
        .A2(SubCellInst_LFInst_1_LFInst_1_n16 ), .ZN(
        SubCellInst_LFInst_1_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst_LFInst_1_LFInst_1_U10  ( .A1(AddRoundKeyOutput[7]), 
        .A2(SubCellInst_LFInst_1_LFInst_1_n15 ), .ZN(
        SubCellInst_LFInst_1_LFInst_1_n16 ) );
  AND2_X1 SubCellInst_LFInst_1_LFInst_1_U9  ( .A1(AddRoundKeyOutput[4]), .A2(
        AddRoundKeyOutput[6]), .ZN(SubCellInst_LFInst_1_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_1_U8  ( .A1(AddRoundKeyOutput[7]), 
        .A2(SubCellInst_LFInst_1_LFInst_1_n14 ), .ZN(
        SubCellInst_LFInst_1_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_1_U7  ( .A1(
        SubCellInst_LFInst_1_LFInst_1_n13 ), .A2(
        SubCellInst_LFInst_1_LFInst_1_n12 ), .ZN(
        SubCellInst_LFInst_1_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_1_U6  ( .A1(AddRoundKeyOutput[4]), 
        .A2(AddRoundKeyOutput[6]), .ZN(SubCellInst_LFInst_1_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_1_U5  ( .A1(
        SubCellInst_LFInst_1_LFInst_1_n11 ), .A2(
        SubCellInst_LFInst_1_LFInst_1_n10 ), .ZN(
        SubCellInst_LFInst_1_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_1_U4  ( .A1(AddRoundKeyOutput[4]), 
        .A2(AddRoundKeyOutput[5]), .ZN(SubCellInst_LFInst_1_LFInst_1_n10 ) );
  INV_X1 SubCellInst_LFInst_1_LFInst_1_U3  ( .A(AddRoundKeyOutput[6]), .ZN(
        SubCellInst_LFInst_1_LFInst_1_n11 ) );
  XNOR2_X1 SubCellInst_LFInst_1_LFInst_0_U6  ( .A(
        SubCellInst_LFInst_1_LFInst_0_n6 ), .B(
        SubCellInst_LFInst_1_LFInst_0_n5 ), .ZN(MCInst1_MC3_v3_2 [3]) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_0_U5  ( .A1(AddRoundKeyOutput[6]), 
        .A2(SubCellInst_LFInst_1_LFInst_0_n4 ), .ZN(
        SubCellInst_LFInst_1_LFInst_0_n5 ) );
  INV_X1 SubCellInst_LFInst_1_LFInst_0_U4  ( .A(AddRoundKeyOutput[5]), .ZN(
        SubCellInst_LFInst_1_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst_LFInst_1_LFInst_0_U3  ( .A(AddRoundKeyOutput[4]), .B(
        AddRoundKeyOutput[7]), .Z(SubCellInst_LFInst_1_LFInst_0_n6 ) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_3_U9  ( .A1(
        SubCellInst_LFInst_2_LFInst_3_n16 ), .A2(
        SubCellInst_LFInst_2_LFInst_3_n15 ), .ZN(MCInst1_MC2_v3_2 [2]) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_3_U8  ( .A1(AddRoundKeyOutput[9]), 
        .A2(SubCellInst_LFInst_2_LFInst_3_n14 ), .ZN(
        SubCellInst_LFInst_2_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst_LFInst_2_LFInst_3_U7  ( .A(AddRoundKeyOutput[11]), .B(
        AddRoundKeyOutput[10]), .Z(SubCellInst_LFInst_2_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_3_U6  ( .A1(
        SubCellInst_LFInst_2_LFInst_3_n13 ), .A2(
        SubCellInst_LFInst_2_LFInst_3_n12 ), .ZN(
        SubCellInst_LFInst_2_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_3_U5  ( .A1(AddRoundKeyOutput[8]), 
        .A2(AddRoundKeyOutput[10]), .ZN(SubCellInst_LFInst_2_LFInst_3_n12 )
         );
  XNOR2_X1 SubCellInst_LFInst_2_LFInst_3_U4  ( .A(AddRoundKeyOutput[8]), .B(
        SubCellInst_LFInst_2_LFInst_3_n11 ), .ZN(
        SubCellInst_LFInst_2_LFInst_3_n13 ) );
  OR2_X1 SubCellInst_LFInst_2_LFInst_3_U3  ( .A1(AddRoundKeyOutput[11]), .A2(
        AddRoundKeyOutput[9]), .ZN(SubCellInst_LFInst_2_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_2_U11  ( .A1(
        SubCellInst_LFInst_2_LFInst_2_n22 ), .A2(
        SubCellInst_LFInst_2_LFInst_2_n21 ), .ZN(MCInst1_MC2_v3_0 [3]) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_2_U10  ( .A1(AddRoundKeyOutput[10]), 
        .A2(SubCellInst_LFInst_2_LFInst_2_n20 ), .ZN(
        SubCellInst_LFInst_2_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst_LFInst_2_LFInst_2_U9  ( .A1(AddRoundKeyOutput[9]), .A2(
        SubCellInst_LFInst_2_LFInst_2_n19 ), .ZN(
        SubCellInst_LFInst_2_LFInst_2_n20 ) );
  INV_X1 SubCellInst_LFInst_2_LFInst_2_U8  ( .A(AddRoundKeyOutput[11]), .ZN(
        SubCellInst_LFInst_2_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_2_U7  ( .A1(
        SubCellInst_LFInst_2_LFInst_2_n18 ), .A2(
        SubCellInst_LFInst_2_LFInst_2_n17 ), .ZN(
        SubCellInst_LFInst_2_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst_LFInst_2_LFInst_2_U6  ( .A(
        SubCellInst_LFInst_2_LFInst_2_n16 ), .B(AddRoundKeyOutput[10]), .Z(
        SubCellInst_LFInst_2_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_2_U5  ( .A1(AddRoundKeyOutput[8]), 
        .A2(AddRoundKeyOutput[9]), .ZN(SubCellInst_LFInst_2_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_2_U4  ( .A1(
        SubCellInst_LFInst_2_LFInst_2_n15 ), .A2(AddRoundKeyOutput[11]), .ZN(
        SubCellInst_LFInst_2_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst_LFInst_2_LFInst_2_U3  ( .A(AddRoundKeyOutput[8]), .B(
        AddRoundKeyOutput[9]), .ZN(SubCellInst_LFInst_2_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_1_U12  ( .A1(
        SubCellInst_LFInst_2_LFInst_1_n18 ), .A2(
        SubCellInst_LFInst_2_LFInst_1_n17 ), .ZN(MCInst1_MC2_v3_0 [2]) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_1_U11  ( .A1(AddRoundKeyOutput[9]), 
        .A2(SubCellInst_LFInst_2_LFInst_1_n16 ), .ZN(
        SubCellInst_LFInst_2_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst_LFInst_2_LFInst_1_U10  ( .A1(AddRoundKeyOutput[11]), 
        .A2(SubCellInst_LFInst_2_LFInst_1_n15 ), .ZN(
        SubCellInst_LFInst_2_LFInst_1_n16 ) );
  AND2_X1 SubCellInst_LFInst_2_LFInst_1_U9  ( .A1(AddRoundKeyOutput[8]), .A2(
        AddRoundKeyOutput[10]), .ZN(SubCellInst_LFInst_2_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_1_U8  ( .A1(AddRoundKeyOutput[11]), 
        .A2(SubCellInst_LFInst_2_LFInst_1_n14 ), .ZN(
        SubCellInst_LFInst_2_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_1_U7  ( .A1(
        SubCellInst_LFInst_2_LFInst_1_n13 ), .A2(
        SubCellInst_LFInst_2_LFInst_1_n12 ), .ZN(
        SubCellInst_LFInst_2_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_1_U6  ( .A1(AddRoundKeyOutput[8]), 
        .A2(AddRoundKeyOutput[10]), .ZN(SubCellInst_LFInst_2_LFInst_1_n12 )
         );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_1_U5  ( .A1(
        SubCellInst_LFInst_2_LFInst_1_n11 ), .A2(
        SubCellInst_LFInst_2_LFInst_1_n10 ), .ZN(
        SubCellInst_LFInst_2_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_1_U4  ( .A1(AddRoundKeyOutput[8]), 
        .A2(AddRoundKeyOutput[9]), .ZN(SubCellInst_LFInst_2_LFInst_1_n10 ) );
  INV_X1 SubCellInst_LFInst_2_LFInst_1_U3  ( .A(AddRoundKeyOutput[10]), .ZN(
        SubCellInst_LFInst_2_LFInst_1_n11 ) );
  XNOR2_X1 SubCellInst_LFInst_2_LFInst_0_U6  ( .A(
        SubCellInst_LFInst_2_LFInst_0_n6 ), .B(
        SubCellInst_LFInst_2_LFInst_0_n5 ), .ZN(MCInst1_MC2_v3_2 [3]) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_0_U5  ( .A1(AddRoundKeyOutput[10]), 
        .A2(SubCellInst_LFInst_2_LFInst_0_n4 ), .ZN(
        SubCellInst_LFInst_2_LFInst_0_n5 ) );
  INV_X1 SubCellInst_LFInst_2_LFInst_0_U4  ( .A(AddRoundKeyOutput[9]), .ZN(
        SubCellInst_LFInst_2_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst_LFInst_2_LFInst_0_U3  ( .A(AddRoundKeyOutput[8]), .B(
        AddRoundKeyOutput[11]), .Z(SubCellInst_LFInst_2_LFInst_0_n6 ) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_3_U9  ( .A1(
        SubCellInst_LFInst_3_LFInst_3_n16 ), .A2(
        SubCellInst_LFInst_3_LFInst_3_n15 ), .ZN(MCInst1_MC1_v3_2 [2]) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_3_U8  ( .A1(AddRoundKeyOutput[13]), 
        .A2(SubCellInst_LFInst_3_LFInst_3_n14 ), .ZN(
        SubCellInst_LFInst_3_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst_LFInst_3_LFInst_3_U7  ( .A(AddRoundKeyOutput[15]), .B(
        AddRoundKeyOutput[14]), .Z(SubCellInst_LFInst_3_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_3_U6  ( .A1(
        SubCellInst_LFInst_3_LFInst_3_n13 ), .A2(
        SubCellInst_LFInst_3_LFInst_3_n12 ), .ZN(
        SubCellInst_LFInst_3_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_3_U5  ( .A1(AddRoundKeyOutput[12]), 
        .A2(AddRoundKeyOutput[14]), .ZN(SubCellInst_LFInst_3_LFInst_3_n12 )
         );
  XNOR2_X1 SubCellInst_LFInst_3_LFInst_3_U4  ( .A(AddRoundKeyOutput[12]), .B(
        SubCellInst_LFInst_3_LFInst_3_n11 ), .ZN(
        SubCellInst_LFInst_3_LFInst_3_n13 ) );
  OR2_X1 SubCellInst_LFInst_3_LFInst_3_U3  ( .A1(AddRoundKeyOutput[15]), .A2(
        AddRoundKeyOutput[13]), .ZN(SubCellInst_LFInst_3_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_2_U11  ( .A1(
        SubCellInst_LFInst_3_LFInst_2_n22 ), .A2(
        SubCellInst_LFInst_3_LFInst_2_n21 ), .ZN(MCInst1_MC1_v3_0 [3]) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_2_U10  ( .A1(AddRoundKeyOutput[14]), 
        .A2(SubCellInst_LFInst_3_LFInst_2_n20 ), .ZN(
        SubCellInst_LFInst_3_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst_LFInst_3_LFInst_2_U9  ( .A1(AddRoundKeyOutput[13]), 
        .A2(SubCellInst_LFInst_3_LFInst_2_n19 ), .ZN(
        SubCellInst_LFInst_3_LFInst_2_n20 ) );
  INV_X1 SubCellInst_LFInst_3_LFInst_2_U8  ( .A(AddRoundKeyOutput[15]), .ZN(
        SubCellInst_LFInst_3_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_2_U7  ( .A1(
        SubCellInst_LFInst_3_LFInst_2_n18 ), .A2(
        SubCellInst_LFInst_3_LFInst_2_n17 ), .ZN(
        SubCellInst_LFInst_3_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst_LFInst_3_LFInst_2_U6  ( .A(
        SubCellInst_LFInst_3_LFInst_2_n16 ), .B(AddRoundKeyOutput[14]), .Z(
        SubCellInst_LFInst_3_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_2_U5  ( .A1(AddRoundKeyOutput[12]), 
        .A2(AddRoundKeyOutput[13]), .ZN(SubCellInst_LFInst_3_LFInst_2_n16 )
         );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_2_U4  ( .A1(
        SubCellInst_LFInst_3_LFInst_2_n15 ), .A2(AddRoundKeyOutput[15]), .ZN(
        SubCellInst_LFInst_3_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst_LFInst_3_LFInst_2_U3  ( .A(AddRoundKeyOutput[12]), .B(
        AddRoundKeyOutput[13]), .ZN(SubCellInst_LFInst_3_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_1_U12  ( .A1(
        SubCellInst_LFInst_3_LFInst_1_n18 ), .A2(
        SubCellInst_LFInst_3_LFInst_1_n17 ), .ZN(MCInst1_MC1_v3_0 [2]) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_1_U11  ( .A1(AddRoundKeyOutput[13]), 
        .A2(SubCellInst_LFInst_3_LFInst_1_n16 ), .ZN(
        SubCellInst_LFInst_3_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst_LFInst_3_LFInst_1_U10  ( .A1(AddRoundKeyOutput[15]), 
        .A2(SubCellInst_LFInst_3_LFInst_1_n15 ), .ZN(
        SubCellInst_LFInst_3_LFInst_1_n16 ) );
  AND2_X1 SubCellInst_LFInst_3_LFInst_1_U9  ( .A1(AddRoundKeyOutput[12]), 
        .A2(AddRoundKeyOutput[14]), .ZN(SubCellInst_LFInst_3_LFInst_1_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_1_U8  ( .A1(AddRoundKeyOutput[15]), 
        .A2(SubCellInst_LFInst_3_LFInst_1_n14 ), .ZN(
        SubCellInst_LFInst_3_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_1_U7  ( .A1(
        SubCellInst_LFInst_3_LFInst_1_n13 ), .A2(
        SubCellInst_LFInst_3_LFInst_1_n12 ), .ZN(
        SubCellInst_LFInst_3_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_1_U6  ( .A1(AddRoundKeyOutput[12]), 
        .A2(AddRoundKeyOutput[14]), .ZN(SubCellInst_LFInst_3_LFInst_1_n12 )
         );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_1_U5  ( .A1(
        SubCellInst_LFInst_3_LFInst_1_n11 ), .A2(
        SubCellInst_LFInst_3_LFInst_1_n10 ), .ZN(
        SubCellInst_LFInst_3_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_1_U4  ( .A1(AddRoundKeyOutput[12]), 
        .A2(AddRoundKeyOutput[13]), .ZN(SubCellInst_LFInst_3_LFInst_1_n10 )
         );
  INV_X1 SubCellInst_LFInst_3_LFInst_1_U3  ( .A(AddRoundKeyOutput[14]), .ZN(
        SubCellInst_LFInst_3_LFInst_1_n11 ) );
  XNOR2_X1 SubCellInst_LFInst_3_LFInst_0_U6  ( .A(
        SubCellInst_LFInst_3_LFInst_0_n6 ), .B(
        SubCellInst_LFInst_3_LFInst_0_n5 ), .ZN(MCInst1_MC1_v3_2 [3]) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_0_U5  ( .A1(AddRoundKeyOutput[14]), 
        .A2(SubCellInst_LFInst_3_LFInst_0_n4 ), .ZN(
        SubCellInst_LFInst_3_LFInst_0_n5 ) );
  INV_X1 SubCellInst_LFInst_3_LFInst_0_U4  ( .A(AddRoundKeyOutput[13]), .ZN(
        SubCellInst_LFInst_3_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst_LFInst_3_LFInst_0_U3  ( .A(AddRoundKeyOutput[12]), .B(
        AddRoundKeyOutput[15]), .Z(SubCellInst_LFInst_3_LFInst_0_n6 ) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_3_U9  ( .A1(
        SubCellInst_LFInst_4_LFInst_3_n16 ), .A2(
        SubCellInst_LFInst_4_LFInst_3_n15 ), .ZN(MCInst1_MC1_v2_0 [0]) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_3_U8  ( .A1(AddRoundKeyOutput[17]), 
        .A2(SubCellInst_LFInst_4_LFInst_3_n14 ), .ZN(
        SubCellInst_LFInst_4_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst_LFInst_4_LFInst_3_U7  ( .A(AddRoundKeyOutput[19]), .B(
        AddRoundKeyOutput[18]), .Z(SubCellInst_LFInst_4_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_3_U6  ( .A1(
        SubCellInst_LFInst_4_LFInst_3_n13 ), .A2(
        SubCellInst_LFInst_4_LFInst_3_n12 ), .ZN(
        SubCellInst_LFInst_4_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_3_U5  ( .A1(AddRoundKeyOutput[16]), 
        .A2(AddRoundKeyOutput[18]), .ZN(SubCellInst_LFInst_4_LFInst_3_n12 )
         );
  XNOR2_X1 SubCellInst_LFInst_4_LFInst_3_U4  ( .A(AddRoundKeyOutput[16]), .B(
        SubCellInst_LFInst_4_LFInst_3_n11 ), .ZN(
        SubCellInst_LFInst_4_LFInst_3_n13 ) );
  OR2_X1 SubCellInst_LFInst_4_LFInst_3_U3  ( .A1(AddRoundKeyOutput[19]), .A2(
        AddRoundKeyOutput[17]), .ZN(SubCellInst_LFInst_4_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_2_U11  ( .A1(
        SubCellInst_LFInst_4_LFInst_2_n22 ), .A2(
        SubCellInst_LFInst_4_LFInst_2_n21 ), .ZN(MCInst1_MC1_v2_0 [3]) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_2_U10  ( .A1(AddRoundKeyOutput[18]), 
        .A2(SubCellInst_LFInst_4_LFInst_2_n20 ), .ZN(
        SubCellInst_LFInst_4_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst_LFInst_4_LFInst_2_U9  ( .A1(AddRoundKeyOutput[17]), 
        .A2(SubCellInst_LFInst_4_LFInst_2_n19 ), .ZN(
        SubCellInst_LFInst_4_LFInst_2_n20 ) );
  INV_X1 SubCellInst_LFInst_4_LFInst_2_U8  ( .A(AddRoundKeyOutput[19]), .ZN(
        SubCellInst_LFInst_4_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_2_U7  ( .A1(
        SubCellInst_LFInst_4_LFInst_2_n18 ), .A2(
        SubCellInst_LFInst_4_LFInst_2_n17 ), .ZN(
        SubCellInst_LFInst_4_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst_LFInst_4_LFInst_2_U6  ( .A(
        SubCellInst_LFInst_4_LFInst_2_n16 ), .B(AddRoundKeyOutput[18]), .Z(
        SubCellInst_LFInst_4_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_2_U5  ( .A1(AddRoundKeyOutput[16]), 
        .A2(AddRoundKeyOutput[17]), .ZN(SubCellInst_LFInst_4_LFInst_2_n16 )
         );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_2_U4  ( .A1(
        SubCellInst_LFInst_4_LFInst_2_n15 ), .A2(AddRoundKeyOutput[19]), .ZN(
        SubCellInst_LFInst_4_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst_LFInst_4_LFInst_2_U3  ( .A(AddRoundKeyOutput[16]), .B(
        AddRoundKeyOutput[17]), .ZN(SubCellInst_LFInst_4_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_1_U12  ( .A1(
        SubCellInst_LFInst_4_LFInst_1_n18 ), .A2(
        SubCellInst_LFInst_4_LFInst_1_n17 ), .ZN(MCInst1_MC1_v2_0 [2]) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_1_U11  ( .A1(AddRoundKeyOutput[17]), 
        .A2(SubCellInst_LFInst_4_LFInst_1_n16 ), .ZN(
        SubCellInst_LFInst_4_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst_LFInst_4_LFInst_1_U10  ( .A1(AddRoundKeyOutput[19]), 
        .A2(SubCellInst_LFInst_4_LFInst_1_n15 ), .ZN(
        SubCellInst_LFInst_4_LFInst_1_n16 ) );
  AND2_X1 SubCellInst_LFInst_4_LFInst_1_U9  ( .A1(AddRoundKeyOutput[16]), 
        .A2(AddRoundKeyOutput[18]), .ZN(SubCellInst_LFInst_4_LFInst_1_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_1_U8  ( .A1(AddRoundKeyOutput[19]), 
        .A2(SubCellInst_LFInst_4_LFInst_1_n14 ), .ZN(
        SubCellInst_LFInst_4_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_1_U7  ( .A1(
        SubCellInst_LFInst_4_LFInst_1_n13 ), .A2(
        SubCellInst_LFInst_4_LFInst_1_n12 ), .ZN(
        SubCellInst_LFInst_4_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_1_U6  ( .A1(AddRoundKeyOutput[16]), 
        .A2(AddRoundKeyOutput[18]), .ZN(SubCellInst_LFInst_4_LFInst_1_n12 )
         );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_1_U5  ( .A1(
        SubCellInst_LFInst_4_LFInst_1_n11 ), .A2(
        SubCellInst_LFInst_4_LFInst_1_n10 ), .ZN(
        SubCellInst_LFInst_4_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_1_U4  ( .A1(AddRoundKeyOutput[16]), 
        .A2(AddRoundKeyOutput[17]), .ZN(SubCellInst_LFInst_4_LFInst_1_n10 )
         );
  INV_X1 SubCellInst_LFInst_4_LFInst_1_U3  ( .A(AddRoundKeyOutput[18]), .ZN(
        SubCellInst_LFInst_4_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_0_U6  ( .A1(AddRoundKeyOutput[18]), 
        .A2(SubCellInst_LFInst_4_LFInst_0_n4 ), .ZN(
        SubCellInst_LFInst_4_LFInst_0_n5 ) );
  INV_X1 SubCellInst_LFInst_4_LFInst_0_U5  ( .A(AddRoundKeyOutput[17]), .ZN(
        SubCellInst_LFInst_4_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst_LFInst_4_LFInst_0_U4  ( .A(AddRoundKeyOutput[16]), .B(
        AddRoundKeyOutput[19]), .Z(SubCellInst_LFInst_4_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst_LFInst_4_LFInst_0_U3  ( .A(
        SubCellInst_LFInst_4_LFInst_0_n6 ), .B(
        SubCellInst_LFInst_4_LFInst_0_n5 ), .ZN(MCInst1_MC1_v2_3 [1]) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_3_U9  ( .A1(
        SubCellInst_LFInst_5_LFInst_3_n16 ), .A2(
        SubCellInst_LFInst_5_LFInst_3_n15 ), .ZN(MCInst1_MC0_v2_0 [0]) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_3_U8  ( .A1(AddRoundKeyOutput[21]), 
        .A2(SubCellInst_LFInst_5_LFInst_3_n14 ), .ZN(
        SubCellInst_LFInst_5_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst_LFInst_5_LFInst_3_U7  ( .A(AddRoundKeyOutput[23]), .B(
        AddRoundKeyOutput[22]), .Z(SubCellInst_LFInst_5_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_3_U6  ( .A1(
        SubCellInst_LFInst_5_LFInst_3_n13 ), .A2(
        SubCellInst_LFInst_5_LFInst_3_n12 ), .ZN(
        SubCellInst_LFInst_5_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_3_U5  ( .A1(AddRoundKeyOutput[20]), 
        .A2(AddRoundKeyOutput[22]), .ZN(SubCellInst_LFInst_5_LFInst_3_n12 )
         );
  XNOR2_X1 SubCellInst_LFInst_5_LFInst_3_U4  ( .A(AddRoundKeyOutput[20]), .B(
        SubCellInst_LFInst_5_LFInst_3_n11 ), .ZN(
        SubCellInst_LFInst_5_LFInst_3_n13 ) );
  OR2_X1 SubCellInst_LFInst_5_LFInst_3_U3  ( .A1(AddRoundKeyOutput[23]), .A2(
        AddRoundKeyOutput[21]), .ZN(SubCellInst_LFInst_5_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_2_U11  ( .A1(
        SubCellInst_LFInst_5_LFInst_2_n22 ), .A2(
        SubCellInst_LFInst_5_LFInst_2_n21 ), .ZN(MCInst1_MC0_v2_0 [3]) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_2_U10  ( .A1(AddRoundKeyOutput[22]), 
        .A2(SubCellInst_LFInst_5_LFInst_2_n20 ), .ZN(
        SubCellInst_LFInst_5_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst_LFInst_5_LFInst_2_U9  ( .A1(AddRoundKeyOutput[21]), 
        .A2(SubCellInst_LFInst_5_LFInst_2_n19 ), .ZN(
        SubCellInst_LFInst_5_LFInst_2_n20 ) );
  INV_X1 SubCellInst_LFInst_5_LFInst_2_U8  ( .A(AddRoundKeyOutput[23]), .ZN(
        SubCellInst_LFInst_5_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_2_U7  ( .A1(
        SubCellInst_LFInst_5_LFInst_2_n18 ), .A2(
        SubCellInst_LFInst_5_LFInst_2_n17 ), .ZN(
        SubCellInst_LFInst_5_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst_LFInst_5_LFInst_2_U6  ( .A(
        SubCellInst_LFInst_5_LFInst_2_n16 ), .B(AddRoundKeyOutput[22]), .Z(
        SubCellInst_LFInst_5_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_2_U5  ( .A1(AddRoundKeyOutput[20]), 
        .A2(AddRoundKeyOutput[21]), .ZN(SubCellInst_LFInst_5_LFInst_2_n16 )
         );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_2_U4  ( .A1(
        SubCellInst_LFInst_5_LFInst_2_n15 ), .A2(AddRoundKeyOutput[23]), .ZN(
        SubCellInst_LFInst_5_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst_LFInst_5_LFInst_2_U3  ( .A(AddRoundKeyOutput[20]), .B(
        AddRoundKeyOutput[21]), .ZN(SubCellInst_LFInst_5_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_1_U12  ( .A1(
        SubCellInst_LFInst_5_LFInst_1_n18 ), .A2(
        SubCellInst_LFInst_5_LFInst_1_n17 ), .ZN(MCInst1_MC0_v2_0 [2]) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_1_U11  ( .A1(AddRoundKeyOutput[21]), 
        .A2(SubCellInst_LFInst_5_LFInst_1_n16 ), .ZN(
        SubCellInst_LFInst_5_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst_LFInst_5_LFInst_1_U10  ( .A1(AddRoundKeyOutput[23]), 
        .A2(SubCellInst_LFInst_5_LFInst_1_n15 ), .ZN(
        SubCellInst_LFInst_5_LFInst_1_n16 ) );
  AND2_X1 SubCellInst_LFInst_5_LFInst_1_U9  ( .A1(AddRoundKeyOutput[20]), 
        .A2(AddRoundKeyOutput[22]), .ZN(SubCellInst_LFInst_5_LFInst_1_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_1_U8  ( .A1(AddRoundKeyOutput[23]), 
        .A2(SubCellInst_LFInst_5_LFInst_1_n14 ), .ZN(
        SubCellInst_LFInst_5_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_1_U7  ( .A1(
        SubCellInst_LFInst_5_LFInst_1_n13 ), .A2(
        SubCellInst_LFInst_5_LFInst_1_n12 ), .ZN(
        SubCellInst_LFInst_5_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_1_U6  ( .A1(AddRoundKeyOutput[20]), 
        .A2(AddRoundKeyOutput[22]), .ZN(SubCellInst_LFInst_5_LFInst_1_n12 )
         );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_1_U5  ( .A1(
        SubCellInst_LFInst_5_LFInst_1_n11 ), .A2(
        SubCellInst_LFInst_5_LFInst_1_n10 ), .ZN(
        SubCellInst_LFInst_5_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_1_U4  ( .A1(AddRoundKeyOutput[20]), 
        .A2(AddRoundKeyOutput[21]), .ZN(SubCellInst_LFInst_5_LFInst_1_n10 )
         );
  INV_X1 SubCellInst_LFInst_5_LFInst_1_U3  ( .A(AddRoundKeyOutput[22]), .ZN(
        SubCellInst_LFInst_5_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_0_U6  ( .A1(AddRoundKeyOutput[22]), 
        .A2(SubCellInst_LFInst_5_LFInst_0_n4 ), .ZN(
        SubCellInst_LFInst_5_LFInst_0_n5 ) );
  INV_X1 SubCellInst_LFInst_5_LFInst_0_U5  ( .A(AddRoundKeyOutput[21]), .ZN(
        SubCellInst_LFInst_5_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst_LFInst_5_LFInst_0_U4  ( .A(AddRoundKeyOutput[20]), .B(
        AddRoundKeyOutput[23]), .Z(SubCellInst_LFInst_5_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst_LFInst_5_LFInst_0_U3  ( .A(
        SubCellInst_LFInst_5_LFInst_0_n6 ), .B(
        SubCellInst_LFInst_5_LFInst_0_n5 ), .ZN(MCInst1_MC0_v2_3 [1]) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_3_U9  ( .A1(
        SubCellInst_LFInst_6_LFInst_3_n16 ), .A2(
        SubCellInst_LFInst_6_LFInst_3_n15 ), .ZN(MCInst1_MC3_v2_0 [0]) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_3_U8  ( .A1(AddRoundKeyOutput[25]), 
        .A2(SubCellInst_LFInst_6_LFInst_3_n14 ), .ZN(
        SubCellInst_LFInst_6_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst_LFInst_6_LFInst_3_U7  ( .A(AddRoundKeyOutput[27]), .B(
        AddRoundKeyOutput[26]), .Z(SubCellInst_LFInst_6_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_3_U6  ( .A1(
        SubCellInst_LFInst_6_LFInst_3_n13 ), .A2(
        SubCellInst_LFInst_6_LFInst_3_n12 ), .ZN(
        SubCellInst_LFInst_6_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_3_U5  ( .A1(AddRoundKeyOutput[24]), 
        .A2(AddRoundKeyOutput[26]), .ZN(SubCellInst_LFInst_6_LFInst_3_n12 )
         );
  XNOR2_X1 SubCellInst_LFInst_6_LFInst_3_U4  ( .A(AddRoundKeyOutput[24]), .B(
        SubCellInst_LFInst_6_LFInst_3_n11 ), .ZN(
        SubCellInst_LFInst_6_LFInst_3_n13 ) );
  OR2_X1 SubCellInst_LFInst_6_LFInst_3_U3  ( .A1(AddRoundKeyOutput[27]), .A2(
        AddRoundKeyOutput[25]), .ZN(SubCellInst_LFInst_6_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_2_U11  ( .A1(
        SubCellInst_LFInst_6_LFInst_2_n22 ), .A2(
        SubCellInst_LFInst_6_LFInst_2_n21 ), .ZN(MCInst1_MC3_v2_0 [3]) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_2_U10  ( .A1(AddRoundKeyOutput[26]), 
        .A2(SubCellInst_LFInst_6_LFInst_2_n20 ), .ZN(
        SubCellInst_LFInst_6_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst_LFInst_6_LFInst_2_U9  ( .A1(AddRoundKeyOutput[25]), 
        .A2(SubCellInst_LFInst_6_LFInst_2_n19 ), .ZN(
        SubCellInst_LFInst_6_LFInst_2_n20 ) );
  INV_X1 SubCellInst_LFInst_6_LFInst_2_U8  ( .A(AddRoundKeyOutput[27]), .ZN(
        SubCellInst_LFInst_6_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_2_U7  ( .A1(
        SubCellInst_LFInst_6_LFInst_2_n18 ), .A2(
        SubCellInst_LFInst_6_LFInst_2_n17 ), .ZN(
        SubCellInst_LFInst_6_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst_LFInst_6_LFInst_2_U6  ( .A(
        SubCellInst_LFInst_6_LFInst_2_n16 ), .B(AddRoundKeyOutput[26]), .Z(
        SubCellInst_LFInst_6_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_2_U5  ( .A1(AddRoundKeyOutput[24]), 
        .A2(AddRoundKeyOutput[25]), .ZN(SubCellInst_LFInst_6_LFInst_2_n16 )
         );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_2_U4  ( .A1(
        SubCellInst_LFInst_6_LFInst_2_n15 ), .A2(AddRoundKeyOutput[27]), .ZN(
        SubCellInst_LFInst_6_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst_LFInst_6_LFInst_2_U3  ( .A(AddRoundKeyOutput[24]), .B(
        AddRoundKeyOutput[25]), .ZN(SubCellInst_LFInst_6_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_1_U12  ( .A1(
        SubCellInst_LFInst_6_LFInst_1_n18 ), .A2(
        SubCellInst_LFInst_6_LFInst_1_n17 ), .ZN(MCInst1_MC3_v2_0 [2]) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_1_U11  ( .A1(AddRoundKeyOutput[25]), 
        .A2(SubCellInst_LFInst_6_LFInst_1_n16 ), .ZN(
        SubCellInst_LFInst_6_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst_LFInst_6_LFInst_1_U10  ( .A1(AddRoundKeyOutput[27]), 
        .A2(SubCellInst_LFInst_6_LFInst_1_n15 ), .ZN(
        SubCellInst_LFInst_6_LFInst_1_n16 ) );
  AND2_X1 SubCellInst_LFInst_6_LFInst_1_U9  ( .A1(AddRoundKeyOutput[24]), 
        .A2(AddRoundKeyOutput[26]), .ZN(SubCellInst_LFInst_6_LFInst_1_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_1_U8  ( .A1(AddRoundKeyOutput[27]), 
        .A2(SubCellInst_LFInst_6_LFInst_1_n14 ), .ZN(
        SubCellInst_LFInst_6_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_1_U7  ( .A1(
        SubCellInst_LFInst_6_LFInst_1_n13 ), .A2(
        SubCellInst_LFInst_6_LFInst_1_n12 ), .ZN(
        SubCellInst_LFInst_6_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_1_U6  ( .A1(AddRoundKeyOutput[24]), 
        .A2(AddRoundKeyOutput[26]), .ZN(SubCellInst_LFInst_6_LFInst_1_n12 )
         );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_1_U5  ( .A1(
        SubCellInst_LFInst_6_LFInst_1_n11 ), .A2(
        SubCellInst_LFInst_6_LFInst_1_n10 ), .ZN(
        SubCellInst_LFInst_6_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_1_U4  ( .A1(AddRoundKeyOutput[24]), 
        .A2(AddRoundKeyOutput[25]), .ZN(SubCellInst_LFInst_6_LFInst_1_n10 )
         );
  INV_X1 SubCellInst_LFInst_6_LFInst_1_U3  ( .A(AddRoundKeyOutput[26]), .ZN(
        SubCellInst_LFInst_6_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_0_U6  ( .A1(AddRoundKeyOutput[26]), 
        .A2(SubCellInst_LFInst_6_LFInst_0_n4 ), .ZN(
        SubCellInst_LFInst_6_LFInst_0_n5 ) );
  INV_X1 SubCellInst_LFInst_6_LFInst_0_U5  ( .A(AddRoundKeyOutput[25]), .ZN(
        SubCellInst_LFInst_6_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst_LFInst_6_LFInst_0_U4  ( .A(AddRoundKeyOutput[24]), .B(
        AddRoundKeyOutput[27]), .Z(SubCellInst_LFInst_6_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst_LFInst_6_LFInst_0_U3  ( .A(
        SubCellInst_LFInst_6_LFInst_0_n6 ), .B(
        SubCellInst_LFInst_6_LFInst_0_n5 ), .ZN(MCInst1_MC3_v2_3 [1]) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_3_U9  ( .A1(
        SubCellInst_LFInst_7_LFInst_3_n16 ), .A2(
        SubCellInst_LFInst_7_LFInst_3_n15 ), .ZN(MCInst1_MC2_v2_0 [0]) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_3_U8  ( .A1(AddRoundKeyOutput[29]), 
        .A2(SubCellInst_LFInst_7_LFInst_3_n14 ), .ZN(
        SubCellInst_LFInst_7_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst_LFInst_7_LFInst_3_U7  ( .A(AddRoundKeyOutput[31]), .B(
        AddRoundKeyOutput[30]), .Z(SubCellInst_LFInst_7_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_3_U6  ( .A1(
        SubCellInst_LFInst_7_LFInst_3_n13 ), .A2(
        SubCellInst_LFInst_7_LFInst_3_n12 ), .ZN(
        SubCellInst_LFInst_7_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_3_U5  ( .A1(AddRoundKeyOutput[28]), 
        .A2(AddRoundKeyOutput[30]), .ZN(SubCellInst_LFInst_7_LFInst_3_n12 )
         );
  XNOR2_X1 SubCellInst_LFInst_7_LFInst_3_U4  ( .A(AddRoundKeyOutput[28]), .B(
        SubCellInst_LFInst_7_LFInst_3_n11 ), .ZN(
        SubCellInst_LFInst_7_LFInst_3_n13 ) );
  OR2_X1 SubCellInst_LFInst_7_LFInst_3_U3  ( .A1(AddRoundKeyOutput[31]), .A2(
        AddRoundKeyOutput[29]), .ZN(SubCellInst_LFInst_7_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_2_U11  ( .A1(
        SubCellInst_LFInst_7_LFInst_2_n22 ), .A2(
        SubCellInst_LFInst_7_LFInst_2_n21 ), .ZN(MCInst1_MC2_v2_0 [3]) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_2_U10  ( .A1(AddRoundKeyOutput[30]), 
        .A2(SubCellInst_LFInst_7_LFInst_2_n20 ), .ZN(
        SubCellInst_LFInst_7_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst_LFInst_7_LFInst_2_U9  ( .A1(AddRoundKeyOutput[29]), 
        .A2(SubCellInst_LFInst_7_LFInst_2_n19 ), .ZN(
        SubCellInst_LFInst_7_LFInst_2_n20 ) );
  INV_X1 SubCellInst_LFInst_7_LFInst_2_U8  ( .A(AddRoundKeyOutput[31]), .ZN(
        SubCellInst_LFInst_7_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_2_U7  ( .A1(
        SubCellInst_LFInst_7_LFInst_2_n18 ), .A2(
        SubCellInst_LFInst_7_LFInst_2_n17 ), .ZN(
        SubCellInst_LFInst_7_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst_LFInst_7_LFInst_2_U6  ( .A(
        SubCellInst_LFInst_7_LFInst_2_n16 ), .B(AddRoundKeyOutput[30]), .Z(
        SubCellInst_LFInst_7_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_2_U5  ( .A1(AddRoundKeyOutput[28]), 
        .A2(AddRoundKeyOutput[29]), .ZN(SubCellInst_LFInst_7_LFInst_2_n16 )
         );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_2_U4  ( .A1(
        SubCellInst_LFInst_7_LFInst_2_n15 ), .A2(AddRoundKeyOutput[31]), .ZN(
        SubCellInst_LFInst_7_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst_LFInst_7_LFInst_2_U3  ( .A(AddRoundKeyOutput[28]), .B(
        AddRoundKeyOutput[29]), .ZN(SubCellInst_LFInst_7_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_1_U12  ( .A1(
        SubCellInst_LFInst_7_LFInst_1_n18 ), .A2(
        SubCellInst_LFInst_7_LFInst_1_n17 ), .ZN(MCInst1_MC2_v2_0 [2]) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_1_U11  ( .A1(AddRoundKeyOutput[29]), 
        .A2(SubCellInst_LFInst_7_LFInst_1_n16 ), .ZN(
        SubCellInst_LFInst_7_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst_LFInst_7_LFInst_1_U10  ( .A1(AddRoundKeyOutput[31]), 
        .A2(SubCellInst_LFInst_7_LFInst_1_n15 ), .ZN(
        SubCellInst_LFInst_7_LFInst_1_n16 ) );
  AND2_X1 SubCellInst_LFInst_7_LFInst_1_U9  ( .A1(AddRoundKeyOutput[28]), 
        .A2(AddRoundKeyOutput[30]), .ZN(SubCellInst_LFInst_7_LFInst_1_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_1_U8  ( .A1(AddRoundKeyOutput[31]), 
        .A2(SubCellInst_LFInst_7_LFInst_1_n14 ), .ZN(
        SubCellInst_LFInst_7_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_1_U7  ( .A1(
        SubCellInst_LFInst_7_LFInst_1_n13 ), .A2(
        SubCellInst_LFInst_7_LFInst_1_n12 ), .ZN(
        SubCellInst_LFInst_7_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_1_U6  ( .A1(AddRoundKeyOutput[28]), 
        .A2(AddRoundKeyOutput[30]), .ZN(SubCellInst_LFInst_7_LFInst_1_n12 )
         );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_1_U5  ( .A1(
        SubCellInst_LFInst_7_LFInst_1_n11 ), .A2(
        SubCellInst_LFInst_7_LFInst_1_n10 ), .ZN(
        SubCellInst_LFInst_7_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_1_U4  ( .A1(AddRoundKeyOutput[28]), 
        .A2(AddRoundKeyOutput[29]), .ZN(SubCellInst_LFInst_7_LFInst_1_n10 )
         );
  INV_X1 SubCellInst_LFInst_7_LFInst_1_U3  ( .A(AddRoundKeyOutput[30]), .ZN(
        SubCellInst_LFInst_7_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_0_U6  ( .A1(AddRoundKeyOutput[30]), 
        .A2(SubCellInst_LFInst_7_LFInst_0_n4 ), .ZN(
        SubCellInst_LFInst_7_LFInst_0_n5 ) );
  INV_X1 SubCellInst_LFInst_7_LFInst_0_U5  ( .A(AddRoundKeyOutput[29]), .ZN(
        SubCellInst_LFInst_7_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst_LFInst_7_LFInst_0_U4  ( .A(AddRoundKeyOutput[28]), .B(
        AddRoundKeyOutput[31]), .Z(SubCellInst_LFInst_7_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst_LFInst_7_LFInst_0_U3  ( .A(
        SubCellInst_LFInst_7_LFInst_0_n6 ), .B(
        SubCellInst_LFInst_7_LFInst_0_n5 ), .ZN(MCInst1_MC2_v2_3 [1]) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_3_U9  ( .A1(
        SubCellInst_LFInst_8_LFInst_3_n16 ), .A2(
        SubCellInst_LFInst_8_LFInst_3_n15 ), .ZN(MCInst1_MC2_v1_3 [0]) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_3_U8  ( .A1(AddRoundKeyOutput[33]), 
        .A2(SubCellInst_LFInst_8_LFInst_3_n14 ), .ZN(
        SubCellInst_LFInst_8_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst_LFInst_8_LFInst_3_U7  ( .A(AddRoundKeyOutput[35]), .B(
        AddRoundKeyOutput[34]), .Z(SubCellInst_LFInst_8_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_3_U6  ( .A1(
        SubCellInst_LFInst_8_LFInst_3_n13 ), .A2(
        SubCellInst_LFInst_8_LFInst_3_n12 ), .ZN(
        SubCellInst_LFInst_8_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_3_U5  ( .A1(AddRoundKeyOutput[32]), 
        .A2(AddRoundKeyOutput[34]), .ZN(SubCellInst_LFInst_8_LFInst_3_n12 )
         );
  XNOR2_X1 SubCellInst_LFInst_8_LFInst_3_U4  ( .A(AddRoundKeyOutput[32]), .B(
        SubCellInst_LFInst_8_LFInst_3_n11 ), .ZN(
        SubCellInst_LFInst_8_LFInst_3_n13 ) );
  OR2_X1 SubCellInst_LFInst_8_LFInst_3_U3  ( .A1(AddRoundKeyOutput[35]), .A2(
        AddRoundKeyOutput[33]), .ZN(SubCellInst_LFInst_8_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_2_U11  ( .A1(
        SubCellInst_LFInst_8_LFInst_2_n22 ), .A2(
        SubCellInst_LFInst_8_LFInst_2_n21 ), .ZN(MCInst1_MC2_v1_3 [3]) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_2_U10  ( .A1(AddRoundKeyOutput[34]), 
        .A2(SubCellInst_LFInst_8_LFInst_2_n20 ), .ZN(
        SubCellInst_LFInst_8_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst_LFInst_8_LFInst_2_U9  ( .A1(AddRoundKeyOutput[33]), 
        .A2(SubCellInst_LFInst_8_LFInst_2_n19 ), .ZN(
        SubCellInst_LFInst_8_LFInst_2_n20 ) );
  INV_X1 SubCellInst_LFInst_8_LFInst_2_U8  ( .A(AddRoundKeyOutput[35]), .ZN(
        SubCellInst_LFInst_8_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_2_U7  ( .A1(
        SubCellInst_LFInst_8_LFInst_2_n18 ), .A2(
        SubCellInst_LFInst_8_LFInst_2_n17 ), .ZN(
        SubCellInst_LFInst_8_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst_LFInst_8_LFInst_2_U6  ( .A(
        SubCellInst_LFInst_8_LFInst_2_n16 ), .B(AddRoundKeyOutput[34]), .Z(
        SubCellInst_LFInst_8_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_2_U5  ( .A1(AddRoundKeyOutput[32]), 
        .A2(AddRoundKeyOutput[33]), .ZN(SubCellInst_LFInst_8_LFInst_2_n16 )
         );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_2_U4  ( .A1(
        SubCellInst_LFInst_8_LFInst_2_n15 ), .A2(AddRoundKeyOutput[35]), .ZN(
        SubCellInst_LFInst_8_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst_LFInst_8_LFInst_2_U3  ( .A(AddRoundKeyOutput[32]), .B(
        AddRoundKeyOutput[33]), .ZN(SubCellInst_LFInst_8_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_1_U12  ( .A1(
        SubCellInst_LFInst_8_LFInst_1_n18 ), .A2(
        SubCellInst_LFInst_8_LFInst_1_n17 ), .ZN(MCInst1_MC2_v1_3 [2]) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_1_U11  ( .A1(AddRoundKeyOutput[33]), 
        .A2(SubCellInst_LFInst_8_LFInst_1_n16 ), .ZN(
        SubCellInst_LFInst_8_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst_LFInst_8_LFInst_1_U10  ( .A1(AddRoundKeyOutput[35]), 
        .A2(SubCellInst_LFInst_8_LFInst_1_n15 ), .ZN(
        SubCellInst_LFInst_8_LFInst_1_n16 ) );
  AND2_X1 SubCellInst_LFInst_8_LFInst_1_U9  ( .A1(AddRoundKeyOutput[32]), 
        .A2(AddRoundKeyOutput[34]), .ZN(SubCellInst_LFInst_8_LFInst_1_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_1_U8  ( .A1(AddRoundKeyOutput[35]), 
        .A2(SubCellInst_LFInst_8_LFInst_1_n14 ), .ZN(
        SubCellInst_LFInst_8_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_1_U7  ( .A1(
        SubCellInst_LFInst_8_LFInst_1_n13 ), .A2(
        SubCellInst_LFInst_8_LFInst_1_n12 ), .ZN(
        SubCellInst_LFInst_8_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_1_U6  ( .A1(AddRoundKeyOutput[32]), 
        .A2(AddRoundKeyOutput[34]), .ZN(SubCellInst_LFInst_8_LFInst_1_n12 )
         );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_1_U5  ( .A1(
        SubCellInst_LFInst_8_LFInst_1_n11 ), .A2(
        SubCellInst_LFInst_8_LFInst_1_n10 ), .ZN(
        SubCellInst_LFInst_8_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_1_U4  ( .A1(AddRoundKeyOutput[32]), 
        .A2(AddRoundKeyOutput[33]), .ZN(SubCellInst_LFInst_8_LFInst_1_n10 )
         );
  INV_X1 SubCellInst_LFInst_8_LFInst_1_U3  ( .A(AddRoundKeyOutput[34]), .ZN(
        SubCellInst_LFInst_8_LFInst_1_n11 ) );
  XNOR2_X1 SubCellInst_LFInst_8_LFInst_0_U6  ( .A(
        SubCellInst_LFInst_8_LFInst_0_n6 ), .B(
        SubCellInst_LFInst_8_LFInst_0_n5 ), .ZN(ShiftRowsOutput[36]) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_0_U5  ( .A1(AddRoundKeyOutput[34]), 
        .A2(SubCellInst_LFInst_8_LFInst_0_n4 ), .ZN(
        SubCellInst_LFInst_8_LFInst_0_n5 ) );
  INV_X1 SubCellInst_LFInst_8_LFInst_0_U4  ( .A(AddRoundKeyOutput[33]), .ZN(
        SubCellInst_LFInst_8_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst_LFInst_8_LFInst_0_U3  ( .A(AddRoundKeyOutput[32]), .B(
        AddRoundKeyOutput[35]), .Z(SubCellInst_LFInst_8_LFInst_0_n6 ) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_3_U9  ( .A1(
        SubCellInst_LFInst_9_LFInst_3_n16 ), .A2(
        SubCellInst_LFInst_9_LFInst_3_n15 ), .ZN(MCInst1_MC1_v1_3 [0]) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_3_U8  ( .A1(AddRoundKeyOutput[37]), 
        .A2(SubCellInst_LFInst_9_LFInst_3_n14 ), .ZN(
        SubCellInst_LFInst_9_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst_LFInst_9_LFInst_3_U7  ( .A(AddRoundKeyOutput[39]), .B(
        AddRoundKeyOutput[38]), .Z(SubCellInst_LFInst_9_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_3_U6  ( .A1(
        SubCellInst_LFInst_9_LFInst_3_n13 ), .A2(
        SubCellInst_LFInst_9_LFInst_3_n12 ), .ZN(
        SubCellInst_LFInst_9_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_3_U5  ( .A1(AddRoundKeyOutput[36]), 
        .A2(AddRoundKeyOutput[38]), .ZN(SubCellInst_LFInst_9_LFInst_3_n12 )
         );
  XNOR2_X1 SubCellInst_LFInst_9_LFInst_3_U4  ( .A(AddRoundKeyOutput[36]), .B(
        SubCellInst_LFInst_9_LFInst_3_n11 ), .ZN(
        SubCellInst_LFInst_9_LFInst_3_n13 ) );
  OR2_X1 SubCellInst_LFInst_9_LFInst_3_U3  ( .A1(AddRoundKeyOutput[39]), .A2(
        AddRoundKeyOutput[37]), .ZN(SubCellInst_LFInst_9_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_2_U11  ( .A1(
        SubCellInst_LFInst_9_LFInst_2_n22 ), .A2(
        SubCellInst_LFInst_9_LFInst_2_n21 ), .ZN(MCInst1_MC1_v1_3 [3]) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_2_U10  ( .A1(AddRoundKeyOutput[38]), 
        .A2(SubCellInst_LFInst_9_LFInst_2_n20 ), .ZN(
        SubCellInst_LFInst_9_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst_LFInst_9_LFInst_2_U9  ( .A1(AddRoundKeyOutput[37]), 
        .A2(SubCellInst_LFInst_9_LFInst_2_n19 ), .ZN(
        SubCellInst_LFInst_9_LFInst_2_n20 ) );
  INV_X1 SubCellInst_LFInst_9_LFInst_2_U8  ( .A(AddRoundKeyOutput[39]), .ZN(
        SubCellInst_LFInst_9_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_2_U7  ( .A1(
        SubCellInst_LFInst_9_LFInst_2_n18 ), .A2(
        SubCellInst_LFInst_9_LFInst_2_n17 ), .ZN(
        SubCellInst_LFInst_9_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst_LFInst_9_LFInst_2_U6  ( .A(
        SubCellInst_LFInst_9_LFInst_2_n16 ), .B(AddRoundKeyOutput[38]), .Z(
        SubCellInst_LFInst_9_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_2_U5  ( .A1(AddRoundKeyOutput[36]), 
        .A2(AddRoundKeyOutput[37]), .ZN(SubCellInst_LFInst_9_LFInst_2_n16 )
         );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_2_U4  ( .A1(
        SubCellInst_LFInst_9_LFInst_2_n15 ), .A2(AddRoundKeyOutput[39]), .ZN(
        SubCellInst_LFInst_9_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst_LFInst_9_LFInst_2_U3  ( .A(AddRoundKeyOutput[36]), .B(
        AddRoundKeyOutput[37]), .ZN(SubCellInst_LFInst_9_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_1_U12  ( .A1(
        SubCellInst_LFInst_9_LFInst_1_n18 ), .A2(
        SubCellInst_LFInst_9_LFInst_1_n17 ), .ZN(MCInst1_MC1_v1_3 [2]) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_1_U11  ( .A1(AddRoundKeyOutput[37]), 
        .A2(SubCellInst_LFInst_9_LFInst_1_n16 ), .ZN(
        SubCellInst_LFInst_9_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst_LFInst_9_LFInst_1_U10  ( .A1(AddRoundKeyOutput[39]), 
        .A2(SubCellInst_LFInst_9_LFInst_1_n15 ), .ZN(
        SubCellInst_LFInst_9_LFInst_1_n16 ) );
  AND2_X1 SubCellInst_LFInst_9_LFInst_1_U9  ( .A1(AddRoundKeyOutput[36]), 
        .A2(AddRoundKeyOutput[38]), .ZN(SubCellInst_LFInst_9_LFInst_1_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_1_U8  ( .A1(AddRoundKeyOutput[39]), 
        .A2(SubCellInst_LFInst_9_LFInst_1_n14 ), .ZN(
        SubCellInst_LFInst_9_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_1_U7  ( .A1(
        SubCellInst_LFInst_9_LFInst_1_n13 ), .A2(
        SubCellInst_LFInst_9_LFInst_1_n12 ), .ZN(
        SubCellInst_LFInst_9_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_1_U6  ( .A1(AddRoundKeyOutput[36]), 
        .A2(AddRoundKeyOutput[38]), .ZN(SubCellInst_LFInst_9_LFInst_1_n12 )
         );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_1_U5  ( .A1(
        SubCellInst_LFInst_9_LFInst_1_n11 ), .A2(
        SubCellInst_LFInst_9_LFInst_1_n10 ), .ZN(
        SubCellInst_LFInst_9_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_1_U4  ( .A1(AddRoundKeyOutput[36]), 
        .A2(AddRoundKeyOutput[37]), .ZN(SubCellInst_LFInst_9_LFInst_1_n10 )
         );
  INV_X1 SubCellInst_LFInst_9_LFInst_1_U3  ( .A(AddRoundKeyOutput[38]), .ZN(
        SubCellInst_LFInst_9_LFInst_1_n11 ) );
  XNOR2_X1 SubCellInst_LFInst_9_LFInst_0_U6  ( .A(
        SubCellInst_LFInst_9_LFInst_0_n6 ), .B(
        SubCellInst_LFInst_9_LFInst_0_n5 ), .ZN(ShiftRowsOutput[40]) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_0_U5  ( .A1(AddRoundKeyOutput[38]), 
        .A2(SubCellInst_LFInst_9_LFInst_0_n4 ), .ZN(
        SubCellInst_LFInst_9_LFInst_0_n5 ) );
  INV_X1 SubCellInst_LFInst_9_LFInst_0_U4  ( .A(AddRoundKeyOutput[37]), .ZN(
        SubCellInst_LFInst_9_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst_LFInst_9_LFInst_0_U3  ( .A(AddRoundKeyOutput[36]), .B(
        AddRoundKeyOutput[39]), .Z(SubCellInst_LFInst_9_LFInst_0_n6 ) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_3_U9  ( .A1(
        SubCellInst_LFInst_10_LFInst_3_n16 ), .A2(
        SubCellInst_LFInst_10_LFInst_3_n15 ), .ZN(MCInst1_MC0_v1_3 [0]) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_3_U8  ( .A1(AddRoundKeyOutput[41]), 
        .A2(SubCellInst_LFInst_10_LFInst_3_n14 ), .ZN(
        SubCellInst_LFInst_10_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst_LFInst_10_LFInst_3_U7  ( .A(AddRoundKeyOutput[43]), .B(
        AddRoundKeyOutput[42]), .Z(SubCellInst_LFInst_10_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_3_U6  ( .A1(
        SubCellInst_LFInst_10_LFInst_3_n13 ), .A2(
        SubCellInst_LFInst_10_LFInst_3_n12 ), .ZN(
        SubCellInst_LFInst_10_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_3_U5  ( .A1(AddRoundKeyOutput[40]), 
        .A2(AddRoundKeyOutput[42]), .ZN(SubCellInst_LFInst_10_LFInst_3_n12 )
         );
  XNOR2_X1 SubCellInst_LFInst_10_LFInst_3_U4  ( .A(AddRoundKeyOutput[40]), 
        .B(SubCellInst_LFInst_10_LFInst_3_n11 ), .ZN(
        SubCellInst_LFInst_10_LFInst_3_n13 ) );
  OR2_X1 SubCellInst_LFInst_10_LFInst_3_U3  ( .A1(AddRoundKeyOutput[43]), 
        .A2(AddRoundKeyOutput[41]), .ZN(SubCellInst_LFInst_10_LFInst_3_n11 )
         );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_2_U11  ( .A1(
        SubCellInst_LFInst_10_LFInst_2_n22 ), .A2(
        SubCellInst_LFInst_10_LFInst_2_n21 ), .ZN(MCInst1_MC0_v1_3 [3]) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_2_U10  ( .A1(AddRoundKeyOutput[42]), 
        .A2(SubCellInst_LFInst_10_LFInst_2_n20 ), .ZN(
        SubCellInst_LFInst_10_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst_LFInst_10_LFInst_2_U9  ( .A1(AddRoundKeyOutput[41]), 
        .A2(SubCellInst_LFInst_10_LFInst_2_n19 ), .ZN(
        SubCellInst_LFInst_10_LFInst_2_n20 ) );
  INV_X1 SubCellInst_LFInst_10_LFInst_2_U8  ( .A(AddRoundKeyOutput[43]), .ZN(
        SubCellInst_LFInst_10_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_2_U7  ( .A1(
        SubCellInst_LFInst_10_LFInst_2_n18 ), .A2(
        SubCellInst_LFInst_10_LFInst_2_n17 ), .ZN(
        SubCellInst_LFInst_10_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst_LFInst_10_LFInst_2_U6  ( .A(
        SubCellInst_LFInst_10_LFInst_2_n16 ), .B(AddRoundKeyOutput[42]), .Z(
        SubCellInst_LFInst_10_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_2_U5  ( .A1(AddRoundKeyOutput[40]), 
        .A2(AddRoundKeyOutput[41]), .ZN(SubCellInst_LFInst_10_LFInst_2_n16 )
         );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_2_U4  ( .A1(
        SubCellInst_LFInst_10_LFInst_2_n15 ), .A2(AddRoundKeyOutput[43]), 
        .ZN(SubCellInst_LFInst_10_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst_LFInst_10_LFInst_2_U3  ( .A(AddRoundKeyOutput[40]), 
        .B(AddRoundKeyOutput[41]), .ZN(SubCellInst_LFInst_10_LFInst_2_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_1_U12  ( .A1(
        SubCellInst_LFInst_10_LFInst_1_n18 ), .A2(
        SubCellInst_LFInst_10_LFInst_1_n17 ), .ZN(MCInst1_MC0_v1_3 [2]) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_1_U11  ( .A1(AddRoundKeyOutput[41]), 
        .A2(SubCellInst_LFInst_10_LFInst_1_n16 ), .ZN(
        SubCellInst_LFInst_10_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst_LFInst_10_LFInst_1_U10  ( .A1(AddRoundKeyOutput[43]), 
        .A2(SubCellInst_LFInst_10_LFInst_1_n15 ), .ZN(
        SubCellInst_LFInst_10_LFInst_1_n16 ) );
  AND2_X1 SubCellInst_LFInst_10_LFInst_1_U9  ( .A1(AddRoundKeyOutput[40]), 
        .A2(AddRoundKeyOutput[42]), .ZN(SubCellInst_LFInst_10_LFInst_1_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_1_U8  ( .A1(AddRoundKeyOutput[43]), 
        .A2(SubCellInst_LFInst_10_LFInst_1_n14 ), .ZN(
        SubCellInst_LFInst_10_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_1_U7  ( .A1(
        SubCellInst_LFInst_10_LFInst_1_n13 ), .A2(
        SubCellInst_LFInst_10_LFInst_1_n12 ), .ZN(
        SubCellInst_LFInst_10_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_1_U6  ( .A1(AddRoundKeyOutput[40]), 
        .A2(AddRoundKeyOutput[42]), .ZN(SubCellInst_LFInst_10_LFInst_1_n12 )
         );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_1_U5  ( .A1(
        SubCellInst_LFInst_10_LFInst_1_n11 ), .A2(
        SubCellInst_LFInst_10_LFInst_1_n10 ), .ZN(
        SubCellInst_LFInst_10_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_1_U4  ( .A1(AddRoundKeyOutput[40]), 
        .A2(AddRoundKeyOutput[41]), .ZN(SubCellInst_LFInst_10_LFInst_1_n10 )
         );
  INV_X1 SubCellInst_LFInst_10_LFInst_1_U3  ( .A(AddRoundKeyOutput[42]), .ZN(
        SubCellInst_LFInst_10_LFInst_1_n11 ) );
  XNOR2_X1 SubCellInst_LFInst_10_LFInst_0_U6  ( .A(
        SubCellInst_LFInst_10_LFInst_0_n6 ), .B(
        SubCellInst_LFInst_10_LFInst_0_n5 ), .ZN(ShiftRowsOutput[44]) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_0_U5  ( .A1(AddRoundKeyOutput[42]), 
        .A2(SubCellInst_LFInst_10_LFInst_0_n4 ), .ZN(
        SubCellInst_LFInst_10_LFInst_0_n5 ) );
  INV_X1 SubCellInst_LFInst_10_LFInst_0_U4  ( .A(AddRoundKeyOutput[41]), .ZN(
        SubCellInst_LFInst_10_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst_LFInst_10_LFInst_0_U3  ( .A(AddRoundKeyOutput[40]), .B(
        AddRoundKeyOutput[43]), .Z(SubCellInst_LFInst_10_LFInst_0_n6 ) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_3_U9  ( .A1(
        SubCellInst_LFInst_11_LFInst_3_n16 ), .A2(
        SubCellInst_LFInst_11_LFInst_3_n15 ), .ZN(MCInst1_MC3_v1_3 [0]) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_3_U8  ( .A1(AddRoundKeyOutput[45]), 
        .A2(SubCellInst_LFInst_11_LFInst_3_n14 ), .ZN(
        SubCellInst_LFInst_11_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst_LFInst_11_LFInst_3_U7  ( .A(AddRoundKeyOutput[47]), .B(
        AddRoundKeyOutput[46]), .Z(SubCellInst_LFInst_11_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_3_U6  ( .A1(
        SubCellInst_LFInst_11_LFInst_3_n13 ), .A2(
        SubCellInst_LFInst_11_LFInst_3_n12 ), .ZN(
        SubCellInst_LFInst_11_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_3_U5  ( .A1(AddRoundKeyOutput[44]), 
        .A2(AddRoundKeyOutput[46]), .ZN(SubCellInst_LFInst_11_LFInst_3_n12 )
         );
  XNOR2_X1 SubCellInst_LFInst_11_LFInst_3_U4  ( .A(AddRoundKeyOutput[44]), 
        .B(SubCellInst_LFInst_11_LFInst_3_n11 ), .ZN(
        SubCellInst_LFInst_11_LFInst_3_n13 ) );
  OR2_X1 SubCellInst_LFInst_11_LFInst_3_U3  ( .A1(AddRoundKeyOutput[47]), 
        .A2(AddRoundKeyOutput[45]), .ZN(SubCellInst_LFInst_11_LFInst_3_n11 )
         );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_2_U11  ( .A1(
        SubCellInst_LFInst_11_LFInst_2_n22 ), .A2(
        SubCellInst_LFInst_11_LFInst_2_n21 ), .ZN(MCInst1_MC3_v1_3 [3]) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_2_U10  ( .A1(AddRoundKeyOutput[46]), 
        .A2(SubCellInst_LFInst_11_LFInst_2_n20 ), .ZN(
        SubCellInst_LFInst_11_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst_LFInst_11_LFInst_2_U9  ( .A1(AddRoundKeyOutput[45]), 
        .A2(SubCellInst_LFInst_11_LFInst_2_n19 ), .ZN(
        SubCellInst_LFInst_11_LFInst_2_n20 ) );
  INV_X1 SubCellInst_LFInst_11_LFInst_2_U8  ( .A(AddRoundKeyOutput[47]), .ZN(
        SubCellInst_LFInst_11_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_2_U7  ( .A1(
        SubCellInst_LFInst_11_LFInst_2_n18 ), .A2(
        SubCellInst_LFInst_11_LFInst_2_n17 ), .ZN(
        SubCellInst_LFInst_11_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst_LFInst_11_LFInst_2_U6  ( .A(
        SubCellInst_LFInst_11_LFInst_2_n16 ), .B(AddRoundKeyOutput[46]), .Z(
        SubCellInst_LFInst_11_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_2_U5  ( .A1(AddRoundKeyOutput[44]), 
        .A2(AddRoundKeyOutput[45]), .ZN(SubCellInst_LFInst_11_LFInst_2_n16 )
         );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_2_U4  ( .A1(
        SubCellInst_LFInst_11_LFInst_2_n15 ), .A2(AddRoundKeyOutput[47]), 
        .ZN(SubCellInst_LFInst_11_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst_LFInst_11_LFInst_2_U3  ( .A(AddRoundKeyOutput[44]), 
        .B(AddRoundKeyOutput[45]), .ZN(SubCellInst_LFInst_11_LFInst_2_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_1_U12  ( .A1(
        SubCellInst_LFInst_11_LFInst_1_n18 ), .A2(
        SubCellInst_LFInst_11_LFInst_1_n17 ), .ZN(MCInst1_MC3_v1_3 [2]) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_1_U11  ( .A1(AddRoundKeyOutput[45]), 
        .A2(SubCellInst_LFInst_11_LFInst_1_n16 ), .ZN(
        SubCellInst_LFInst_11_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst_LFInst_11_LFInst_1_U10  ( .A1(AddRoundKeyOutput[47]), 
        .A2(SubCellInst_LFInst_11_LFInst_1_n15 ), .ZN(
        SubCellInst_LFInst_11_LFInst_1_n16 ) );
  AND2_X1 SubCellInst_LFInst_11_LFInst_1_U9  ( .A1(AddRoundKeyOutput[44]), 
        .A2(AddRoundKeyOutput[46]), .ZN(SubCellInst_LFInst_11_LFInst_1_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_1_U8  ( .A1(AddRoundKeyOutput[47]), 
        .A2(SubCellInst_LFInst_11_LFInst_1_n14 ), .ZN(
        SubCellInst_LFInst_11_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_1_U7  ( .A1(
        SubCellInst_LFInst_11_LFInst_1_n13 ), .A2(
        SubCellInst_LFInst_11_LFInst_1_n12 ), .ZN(
        SubCellInst_LFInst_11_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_1_U6  ( .A1(AddRoundKeyOutput[44]), 
        .A2(AddRoundKeyOutput[46]), .ZN(SubCellInst_LFInst_11_LFInst_1_n12 )
         );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_1_U5  ( .A1(
        SubCellInst_LFInst_11_LFInst_1_n11 ), .A2(
        SubCellInst_LFInst_11_LFInst_1_n10 ), .ZN(
        SubCellInst_LFInst_11_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_1_U4  ( .A1(AddRoundKeyOutput[44]), 
        .A2(AddRoundKeyOutput[45]), .ZN(SubCellInst_LFInst_11_LFInst_1_n10 )
         );
  INV_X1 SubCellInst_LFInst_11_LFInst_1_U3  ( .A(AddRoundKeyOutput[46]), .ZN(
        SubCellInst_LFInst_11_LFInst_1_n11 ) );
  XNOR2_X1 SubCellInst_LFInst_11_LFInst_0_U6  ( .A(
        SubCellInst_LFInst_11_LFInst_0_n6 ), .B(
        SubCellInst_LFInst_11_LFInst_0_n5 ), .ZN(ShiftRowsOutput[32]) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_0_U5  ( .A1(AddRoundKeyOutput[46]), 
        .A2(SubCellInst_LFInst_11_LFInst_0_n4 ), .ZN(
        SubCellInst_LFInst_11_LFInst_0_n5 ) );
  INV_X1 SubCellInst_LFInst_11_LFInst_0_U4  ( .A(AddRoundKeyOutput[45]), .ZN(
        SubCellInst_LFInst_11_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst_LFInst_11_LFInst_0_U3  ( .A(AddRoundKeyOutput[44]), .B(
        AddRoundKeyOutput[47]), .Z(SubCellInst_LFInst_11_LFInst_0_n6 ) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_3_U9  ( .A1(
        SubCellInst_LFInst_12_LFInst_3_n16 ), .A2(
        SubCellInst_LFInst_12_LFInst_3_n15 ), .ZN(MCInst1_MC3_v0_3 [0]) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_3_U8  ( .A1(AddRoundKeyOutput[49]), 
        .A2(SubCellInst_LFInst_12_LFInst_3_n14 ), .ZN(
        SubCellInst_LFInst_12_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst_LFInst_12_LFInst_3_U7  ( .A(AddRoundKeyOutput[51]), .B(
        AddRoundKeyOutput[50]), .Z(SubCellInst_LFInst_12_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_3_U6  ( .A1(
        SubCellInst_LFInst_12_LFInst_3_n13 ), .A2(
        SubCellInst_LFInst_12_LFInst_3_n12 ), .ZN(
        SubCellInst_LFInst_12_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_3_U5  ( .A1(AddRoundKeyOutput[48]), 
        .A2(AddRoundKeyOutput[50]), .ZN(SubCellInst_LFInst_12_LFInst_3_n12 )
         );
  XNOR2_X1 SubCellInst_LFInst_12_LFInst_3_U4  ( .A(AddRoundKeyOutput[48]), 
        .B(SubCellInst_LFInst_12_LFInst_3_n11 ), .ZN(
        SubCellInst_LFInst_12_LFInst_3_n13 ) );
  OR2_X1 SubCellInst_LFInst_12_LFInst_3_U3  ( .A1(AddRoundKeyOutput[51]), 
        .A2(AddRoundKeyOutput[49]), .ZN(SubCellInst_LFInst_12_LFInst_3_n11 )
         );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_2_U11  ( .A1(
        SubCellInst_LFInst_12_LFInst_2_n22 ), .A2(
        SubCellInst_LFInst_12_LFInst_2_n21 ), .ZN(MCInst1_MC3_v0_3 [3]) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_2_U10  ( .A1(AddRoundKeyOutput[50]), 
        .A2(SubCellInst_LFInst_12_LFInst_2_n20 ), .ZN(
        SubCellInst_LFInst_12_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst_LFInst_12_LFInst_2_U9  ( .A1(AddRoundKeyOutput[49]), 
        .A2(SubCellInst_LFInst_12_LFInst_2_n19 ), .ZN(
        SubCellInst_LFInst_12_LFInst_2_n20 ) );
  INV_X1 SubCellInst_LFInst_12_LFInst_2_U8  ( .A(AddRoundKeyOutput[51]), .ZN(
        SubCellInst_LFInst_12_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_2_U7  ( .A1(
        SubCellInst_LFInst_12_LFInst_2_n18 ), .A2(
        SubCellInst_LFInst_12_LFInst_2_n17 ), .ZN(
        SubCellInst_LFInst_12_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst_LFInst_12_LFInst_2_U6  ( .A(
        SubCellInst_LFInst_12_LFInst_2_n16 ), .B(AddRoundKeyOutput[50]), .Z(
        SubCellInst_LFInst_12_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_2_U5  ( .A1(AddRoundKeyOutput[48]), 
        .A2(AddRoundKeyOutput[49]), .ZN(SubCellInst_LFInst_12_LFInst_2_n16 )
         );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_2_U4  ( .A1(
        SubCellInst_LFInst_12_LFInst_2_n15 ), .A2(AddRoundKeyOutput[51]), 
        .ZN(SubCellInst_LFInst_12_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst_LFInst_12_LFInst_2_U3  ( .A(AddRoundKeyOutput[48]), 
        .B(AddRoundKeyOutput[49]), .ZN(SubCellInst_LFInst_12_LFInst_2_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_1_U12  ( .A1(
        SubCellInst_LFInst_12_LFInst_1_n18 ), .A2(
        SubCellInst_LFInst_12_LFInst_1_n17 ), .ZN(MCInst1_MC3_v0_0 [3]) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_1_U11  ( .A1(AddRoundKeyOutput[49]), 
        .A2(SubCellInst_LFInst_12_LFInst_1_n16 ), .ZN(
        SubCellInst_LFInst_12_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst_LFInst_12_LFInst_1_U10  ( .A1(AddRoundKeyOutput[51]), 
        .A2(SubCellInst_LFInst_12_LFInst_1_n15 ), .ZN(
        SubCellInst_LFInst_12_LFInst_1_n16 ) );
  AND2_X1 SubCellInst_LFInst_12_LFInst_1_U9  ( .A1(AddRoundKeyOutput[48]), 
        .A2(AddRoundKeyOutput[50]), .ZN(SubCellInst_LFInst_12_LFInst_1_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_1_U8  ( .A1(AddRoundKeyOutput[51]), 
        .A2(SubCellInst_LFInst_12_LFInst_1_n14 ), .ZN(
        SubCellInst_LFInst_12_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_1_U7  ( .A1(
        SubCellInst_LFInst_12_LFInst_1_n13 ), .A2(
        SubCellInst_LFInst_12_LFInst_1_n12 ), .ZN(
        SubCellInst_LFInst_12_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_1_U6  ( .A1(AddRoundKeyOutput[48]), 
        .A2(AddRoundKeyOutput[50]), .ZN(SubCellInst_LFInst_12_LFInst_1_n12 )
         );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_1_U5  ( .A1(
        SubCellInst_LFInst_12_LFInst_1_n11 ), .A2(
        SubCellInst_LFInst_12_LFInst_1_n10 ), .ZN(
        SubCellInst_LFInst_12_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_1_U4  ( .A1(AddRoundKeyOutput[48]), 
        .A2(AddRoundKeyOutput[49]), .ZN(SubCellInst_LFInst_12_LFInst_1_n10 )
         );
  INV_X1 SubCellInst_LFInst_12_LFInst_1_U3  ( .A(AddRoundKeyOutput[50]), .ZN(
        SubCellInst_LFInst_12_LFInst_1_n11 ) );
  XNOR2_X1 SubCellInst_LFInst_12_LFInst_0_U6  ( .A(
        SubCellInst_LFInst_12_LFInst_0_n6 ), .B(
        SubCellInst_LFInst_12_LFInst_0_n5 ), .ZN(ShiftRowsOutput[48]) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_0_U5  ( .A1(AddRoundKeyOutput[50]), 
        .A2(SubCellInst_LFInst_12_LFInst_0_n4 ), .ZN(
        SubCellInst_LFInst_12_LFInst_0_n5 ) );
  INV_X1 SubCellInst_LFInst_12_LFInst_0_U4  ( .A(AddRoundKeyOutput[49]), .ZN(
        SubCellInst_LFInst_12_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst_LFInst_12_LFInst_0_U3  ( .A(AddRoundKeyOutput[48]), .B(
        AddRoundKeyOutput[51]), .Z(SubCellInst_LFInst_12_LFInst_0_n6 ) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_3_U9  ( .A1(
        SubCellInst_LFInst_13_LFInst_3_n16 ), .A2(
        SubCellInst_LFInst_13_LFInst_3_n15 ), .ZN(MCInst1_MC2_v0_3 [0]) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_3_U8  ( .A1(AddRoundKeyOutput[53]), 
        .A2(SubCellInst_LFInst_13_LFInst_3_n14 ), .ZN(
        SubCellInst_LFInst_13_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst_LFInst_13_LFInst_3_U7  ( .A(AddRoundKeyOutput[55]), .B(
        AddRoundKeyOutput[54]), .Z(SubCellInst_LFInst_13_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_3_U6  ( .A1(
        SubCellInst_LFInst_13_LFInst_3_n13 ), .A2(
        SubCellInst_LFInst_13_LFInst_3_n12 ), .ZN(
        SubCellInst_LFInst_13_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_3_U5  ( .A1(AddRoundKeyOutput[52]), 
        .A2(AddRoundKeyOutput[54]), .ZN(SubCellInst_LFInst_13_LFInst_3_n12 )
         );
  XNOR2_X1 SubCellInst_LFInst_13_LFInst_3_U4  ( .A(AddRoundKeyOutput[52]), 
        .B(SubCellInst_LFInst_13_LFInst_3_n11 ), .ZN(
        SubCellInst_LFInst_13_LFInst_3_n13 ) );
  OR2_X1 SubCellInst_LFInst_13_LFInst_3_U3  ( .A1(AddRoundKeyOutput[55]), 
        .A2(AddRoundKeyOutput[53]), .ZN(SubCellInst_LFInst_13_LFInst_3_n11 )
         );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_2_U11  ( .A1(
        SubCellInst_LFInst_13_LFInst_2_n22 ), .A2(
        SubCellInst_LFInst_13_LFInst_2_n21 ), .ZN(MCInst1_MC2_v0_3 [3]) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_2_U10  ( .A1(AddRoundKeyOutput[54]), 
        .A2(SubCellInst_LFInst_13_LFInst_2_n20 ), .ZN(
        SubCellInst_LFInst_13_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst_LFInst_13_LFInst_2_U9  ( .A1(AddRoundKeyOutput[53]), 
        .A2(SubCellInst_LFInst_13_LFInst_2_n19 ), .ZN(
        SubCellInst_LFInst_13_LFInst_2_n20 ) );
  INV_X1 SubCellInst_LFInst_13_LFInst_2_U8  ( .A(AddRoundKeyOutput[55]), .ZN(
        SubCellInst_LFInst_13_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_2_U7  ( .A1(
        SubCellInst_LFInst_13_LFInst_2_n18 ), .A2(
        SubCellInst_LFInst_13_LFInst_2_n17 ), .ZN(
        SubCellInst_LFInst_13_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst_LFInst_13_LFInst_2_U6  ( .A(
        SubCellInst_LFInst_13_LFInst_2_n16 ), .B(AddRoundKeyOutput[54]), .Z(
        SubCellInst_LFInst_13_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_2_U5  ( .A1(AddRoundKeyOutput[52]), 
        .A2(AddRoundKeyOutput[53]), .ZN(SubCellInst_LFInst_13_LFInst_2_n16 )
         );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_2_U4  ( .A1(
        SubCellInst_LFInst_13_LFInst_2_n15 ), .A2(AddRoundKeyOutput[55]), 
        .ZN(SubCellInst_LFInst_13_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst_LFInst_13_LFInst_2_U3  ( .A(AddRoundKeyOutput[52]), 
        .B(AddRoundKeyOutput[53]), .ZN(SubCellInst_LFInst_13_LFInst_2_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_1_U12  ( .A1(
        SubCellInst_LFInst_13_LFInst_1_n18 ), .A2(
        SubCellInst_LFInst_13_LFInst_1_n17 ), .ZN(MCInst1_MC2_v0_0 [3]) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_1_U11  ( .A1(AddRoundKeyOutput[53]), 
        .A2(SubCellInst_LFInst_13_LFInst_1_n16 ), .ZN(
        SubCellInst_LFInst_13_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst_LFInst_13_LFInst_1_U10  ( .A1(AddRoundKeyOutput[55]), 
        .A2(SubCellInst_LFInst_13_LFInst_1_n15 ), .ZN(
        SubCellInst_LFInst_13_LFInst_1_n16 ) );
  AND2_X1 SubCellInst_LFInst_13_LFInst_1_U9  ( .A1(AddRoundKeyOutput[52]), 
        .A2(AddRoundKeyOutput[54]), .ZN(SubCellInst_LFInst_13_LFInst_1_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_1_U8  ( .A1(AddRoundKeyOutput[55]), 
        .A2(SubCellInst_LFInst_13_LFInst_1_n14 ), .ZN(
        SubCellInst_LFInst_13_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_1_U7  ( .A1(
        SubCellInst_LFInst_13_LFInst_1_n13 ), .A2(
        SubCellInst_LFInst_13_LFInst_1_n12 ), .ZN(
        SubCellInst_LFInst_13_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_1_U6  ( .A1(AddRoundKeyOutput[52]), 
        .A2(AddRoundKeyOutput[54]), .ZN(SubCellInst_LFInst_13_LFInst_1_n12 )
         );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_1_U5  ( .A1(
        SubCellInst_LFInst_13_LFInst_1_n11 ), .A2(
        SubCellInst_LFInst_13_LFInst_1_n10 ), .ZN(
        SubCellInst_LFInst_13_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_1_U4  ( .A1(AddRoundKeyOutput[52]), 
        .A2(AddRoundKeyOutput[53]), .ZN(SubCellInst_LFInst_13_LFInst_1_n10 )
         );
  INV_X1 SubCellInst_LFInst_13_LFInst_1_U3  ( .A(AddRoundKeyOutput[54]), .ZN(
        SubCellInst_LFInst_13_LFInst_1_n11 ) );
  XNOR2_X1 SubCellInst_LFInst_13_LFInst_0_U6  ( .A(
        SubCellInst_LFInst_13_LFInst_0_n6 ), .B(
        SubCellInst_LFInst_13_LFInst_0_n5 ), .ZN(ShiftRowsOutput[52]) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_0_U5  ( .A1(AddRoundKeyOutput[54]), 
        .A2(SubCellInst_LFInst_13_LFInst_0_n4 ), .ZN(
        SubCellInst_LFInst_13_LFInst_0_n5 ) );
  INV_X1 SubCellInst_LFInst_13_LFInst_0_U4  ( .A(AddRoundKeyOutput[53]), .ZN(
        SubCellInst_LFInst_13_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst_LFInst_13_LFInst_0_U3  ( .A(AddRoundKeyOutput[52]), .B(
        AddRoundKeyOutput[55]), .Z(SubCellInst_LFInst_13_LFInst_0_n6 ) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_3_U9  ( .A1(
        SubCellInst_LFInst_14_LFInst_3_n16 ), .A2(
        SubCellInst_LFInst_14_LFInst_3_n15 ), .ZN(MCInst1_MC1_v0_3 [0]) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_3_U8  ( .A1(AddRoundKeyOutput[57]), 
        .A2(SubCellInst_LFInst_14_LFInst_3_n14 ), .ZN(
        SubCellInst_LFInst_14_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst_LFInst_14_LFInst_3_U7  ( .A(AddRoundKeyOutput[59]), .B(
        AddRoundKeyOutput[58]), .Z(SubCellInst_LFInst_14_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_3_U6  ( .A1(
        SubCellInst_LFInst_14_LFInst_3_n13 ), .A2(
        SubCellInst_LFInst_14_LFInst_3_n12 ), .ZN(
        SubCellInst_LFInst_14_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_3_U5  ( .A1(AddRoundKeyOutput[56]), 
        .A2(AddRoundKeyOutput[58]), .ZN(SubCellInst_LFInst_14_LFInst_3_n12 )
         );
  XNOR2_X1 SubCellInst_LFInst_14_LFInst_3_U4  ( .A(AddRoundKeyOutput[56]), 
        .B(SubCellInst_LFInst_14_LFInst_3_n11 ), .ZN(
        SubCellInst_LFInst_14_LFInst_3_n13 ) );
  OR2_X1 SubCellInst_LFInst_14_LFInst_3_U3  ( .A1(AddRoundKeyOutput[59]), 
        .A2(AddRoundKeyOutput[57]), .ZN(SubCellInst_LFInst_14_LFInst_3_n11 )
         );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_2_U11  ( .A1(
        SubCellInst_LFInst_14_LFInst_2_n22 ), .A2(
        SubCellInst_LFInst_14_LFInst_2_n21 ), .ZN(MCInst1_MC1_v0_3 [3]) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_2_U10  ( .A1(AddRoundKeyOutput[58]), 
        .A2(SubCellInst_LFInst_14_LFInst_2_n20 ), .ZN(
        SubCellInst_LFInst_14_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst_LFInst_14_LFInst_2_U9  ( .A1(AddRoundKeyOutput[57]), 
        .A2(SubCellInst_LFInst_14_LFInst_2_n19 ), .ZN(
        SubCellInst_LFInst_14_LFInst_2_n20 ) );
  INV_X1 SubCellInst_LFInst_14_LFInst_2_U8  ( .A(AddRoundKeyOutput[59]), .ZN(
        SubCellInst_LFInst_14_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_2_U7  ( .A1(
        SubCellInst_LFInst_14_LFInst_2_n18 ), .A2(
        SubCellInst_LFInst_14_LFInst_2_n17 ), .ZN(
        SubCellInst_LFInst_14_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst_LFInst_14_LFInst_2_U6  ( .A(
        SubCellInst_LFInst_14_LFInst_2_n16 ), .B(AddRoundKeyOutput[58]), .Z(
        SubCellInst_LFInst_14_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_2_U5  ( .A1(AddRoundKeyOutput[56]), 
        .A2(AddRoundKeyOutput[57]), .ZN(SubCellInst_LFInst_14_LFInst_2_n16 )
         );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_2_U4  ( .A1(
        SubCellInst_LFInst_14_LFInst_2_n15 ), .A2(AddRoundKeyOutput[59]), 
        .ZN(SubCellInst_LFInst_14_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst_LFInst_14_LFInst_2_U3  ( .A(AddRoundKeyOutput[56]), 
        .B(AddRoundKeyOutput[57]), .ZN(SubCellInst_LFInst_14_LFInst_2_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_1_U12  ( .A1(
        SubCellInst_LFInst_14_LFInst_1_n18 ), .A2(
        SubCellInst_LFInst_14_LFInst_1_n17 ), .ZN(MCInst1_MC1_v0_0 [3]) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_1_U11  ( .A1(AddRoundKeyOutput[57]), 
        .A2(SubCellInst_LFInst_14_LFInst_1_n16 ), .ZN(
        SubCellInst_LFInst_14_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst_LFInst_14_LFInst_1_U10  ( .A1(AddRoundKeyOutput[59]), 
        .A2(SubCellInst_LFInst_14_LFInst_1_n15 ), .ZN(
        SubCellInst_LFInst_14_LFInst_1_n16 ) );
  AND2_X1 SubCellInst_LFInst_14_LFInst_1_U9  ( .A1(AddRoundKeyOutput[56]), 
        .A2(AddRoundKeyOutput[58]), .ZN(SubCellInst_LFInst_14_LFInst_1_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_1_U8  ( .A1(AddRoundKeyOutput[59]), 
        .A2(SubCellInst_LFInst_14_LFInst_1_n14 ), .ZN(
        SubCellInst_LFInst_14_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_1_U7  ( .A1(
        SubCellInst_LFInst_14_LFInst_1_n13 ), .A2(
        SubCellInst_LFInst_14_LFInst_1_n12 ), .ZN(
        SubCellInst_LFInst_14_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_1_U6  ( .A1(AddRoundKeyOutput[56]), 
        .A2(AddRoundKeyOutput[58]), .ZN(SubCellInst_LFInst_14_LFInst_1_n12 )
         );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_1_U5  ( .A1(
        SubCellInst_LFInst_14_LFInst_1_n11 ), .A2(
        SubCellInst_LFInst_14_LFInst_1_n10 ), .ZN(
        SubCellInst_LFInst_14_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_1_U4  ( .A1(AddRoundKeyOutput[56]), 
        .A2(AddRoundKeyOutput[57]), .ZN(SubCellInst_LFInst_14_LFInst_1_n10 )
         );
  INV_X1 SubCellInst_LFInst_14_LFInst_1_U3  ( .A(AddRoundKeyOutput[58]), .ZN(
        SubCellInst_LFInst_14_LFInst_1_n11 ) );
  XNOR2_X1 SubCellInst_LFInst_14_LFInst_0_U6  ( .A(
        SubCellInst_LFInst_14_LFInst_0_n6 ), .B(
        SubCellInst_LFInst_14_LFInst_0_n5 ), .ZN(ShiftRowsOutput[56]) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_0_U5  ( .A1(AddRoundKeyOutput[58]), 
        .A2(SubCellInst_LFInst_14_LFInst_0_n4 ), .ZN(
        SubCellInst_LFInst_14_LFInst_0_n5 ) );
  INV_X1 SubCellInst_LFInst_14_LFInst_0_U4  ( .A(AddRoundKeyOutput[57]), .ZN(
        SubCellInst_LFInst_14_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst_LFInst_14_LFInst_0_U3  ( .A(AddRoundKeyOutput[56]), .B(
        AddRoundKeyOutput[59]), .Z(SubCellInst_LFInst_14_LFInst_0_n6 ) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_3_U9  ( .A1(
        SubCellInst_LFInst_15_LFInst_3_n16 ), .A2(
        SubCellInst_LFInst_15_LFInst_3_n15 ), .ZN(MCInst1_MC0_v0_3 [0]) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_3_U8  ( .A1(AddRoundKeyOutput[61]), 
        .A2(SubCellInst_LFInst_15_LFInst_3_n14 ), .ZN(
        SubCellInst_LFInst_15_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst_LFInst_15_LFInst_3_U7  ( .A(AddRoundKeyOutput[63]), .B(
        AddRoundKeyOutput[62]), .Z(SubCellInst_LFInst_15_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_3_U6  ( .A1(
        SubCellInst_LFInst_15_LFInst_3_n13 ), .A2(
        SubCellInst_LFInst_15_LFInst_3_n12 ), .ZN(
        SubCellInst_LFInst_15_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_3_U5  ( .A1(AddRoundKeyOutput[60]), 
        .A2(AddRoundKeyOutput[62]), .ZN(SubCellInst_LFInst_15_LFInst_3_n12 )
         );
  XNOR2_X1 SubCellInst_LFInst_15_LFInst_3_U4  ( .A(AddRoundKeyOutput[60]), 
        .B(SubCellInst_LFInst_15_LFInst_3_n11 ), .ZN(
        SubCellInst_LFInst_15_LFInst_3_n13 ) );
  OR2_X1 SubCellInst_LFInst_15_LFInst_3_U3  ( .A1(AddRoundKeyOutput[63]), 
        .A2(AddRoundKeyOutput[61]), .ZN(SubCellInst_LFInst_15_LFInst_3_n11 )
         );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_2_U11  ( .A1(
        SubCellInst_LFInst_15_LFInst_2_n22 ), .A2(
        SubCellInst_LFInst_15_LFInst_2_n21 ), .ZN(MCInst1_MC0_v0_3 [3]) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_2_U10  ( .A1(AddRoundKeyOutput[62]), 
        .A2(SubCellInst_LFInst_15_LFInst_2_n20 ), .ZN(
        SubCellInst_LFInst_15_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst_LFInst_15_LFInst_2_U9  ( .A1(AddRoundKeyOutput[61]), 
        .A2(SubCellInst_LFInst_15_LFInst_2_n19 ), .ZN(
        SubCellInst_LFInst_15_LFInst_2_n20 ) );
  INV_X1 SubCellInst_LFInst_15_LFInst_2_U8  ( .A(AddRoundKeyOutput[63]), .ZN(
        SubCellInst_LFInst_15_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_2_U7  ( .A1(
        SubCellInst_LFInst_15_LFInst_2_n18 ), .A2(
        SubCellInst_LFInst_15_LFInst_2_n17 ), .ZN(
        SubCellInst_LFInst_15_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst_LFInst_15_LFInst_2_U6  ( .A(
        SubCellInst_LFInst_15_LFInst_2_n16 ), .B(AddRoundKeyOutput[62]), .Z(
        SubCellInst_LFInst_15_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_2_U5  ( .A1(AddRoundKeyOutput[60]), 
        .A2(AddRoundKeyOutput[61]), .ZN(SubCellInst_LFInst_15_LFInst_2_n16 )
         );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_2_U4  ( .A1(
        SubCellInst_LFInst_15_LFInst_2_n15 ), .A2(AddRoundKeyOutput[63]), 
        .ZN(SubCellInst_LFInst_15_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst_LFInst_15_LFInst_2_U3  ( .A(AddRoundKeyOutput[60]), 
        .B(AddRoundKeyOutput[61]), .ZN(SubCellInst_LFInst_15_LFInst_2_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_1_U12  ( .A1(
        SubCellInst_LFInst_15_LFInst_1_n18 ), .A2(
        SubCellInst_LFInst_15_LFInst_1_n17 ), .ZN(MCInst1_MC0_v0_0 [3]) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_1_U11  ( .A1(AddRoundKeyOutput[61]), 
        .A2(SubCellInst_LFInst_15_LFInst_1_n16 ), .ZN(
        SubCellInst_LFInst_15_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst_LFInst_15_LFInst_1_U10  ( .A1(AddRoundKeyOutput[63]), 
        .A2(SubCellInst_LFInst_15_LFInst_1_n15 ), .ZN(
        SubCellInst_LFInst_15_LFInst_1_n16 ) );
  AND2_X1 SubCellInst_LFInst_15_LFInst_1_U9  ( .A1(AddRoundKeyOutput[60]), 
        .A2(AddRoundKeyOutput[62]), .ZN(SubCellInst_LFInst_15_LFInst_1_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_1_U8  ( .A1(AddRoundKeyOutput[63]), 
        .A2(SubCellInst_LFInst_15_LFInst_1_n14 ), .ZN(
        SubCellInst_LFInst_15_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_1_U7  ( .A1(
        SubCellInst_LFInst_15_LFInst_1_n13 ), .A2(
        SubCellInst_LFInst_15_LFInst_1_n12 ), .ZN(
        SubCellInst_LFInst_15_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_1_U6  ( .A1(AddRoundKeyOutput[60]), 
        .A2(AddRoundKeyOutput[62]), .ZN(SubCellInst_LFInst_15_LFInst_1_n12 )
         );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_1_U5  ( .A1(
        SubCellInst_LFInst_15_LFInst_1_n11 ), .A2(
        SubCellInst_LFInst_15_LFInst_1_n10 ), .ZN(
        SubCellInst_LFInst_15_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_1_U4  ( .A1(AddRoundKeyOutput[60]), 
        .A2(AddRoundKeyOutput[61]), .ZN(SubCellInst_LFInst_15_LFInst_1_n10 )
         );
  INV_X1 SubCellInst_LFInst_15_LFInst_1_U3  ( .A(AddRoundKeyOutput[62]), .ZN(
        SubCellInst_LFInst_15_LFInst_1_n11 ) );
  XNOR2_X1 SubCellInst_LFInst_15_LFInst_0_U6  ( .A(
        SubCellInst_LFInst_15_LFInst_0_n6 ), .B(
        SubCellInst_LFInst_15_LFInst_0_n5 ), .ZN(ShiftRowsOutput[60]) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_0_U5  ( .A1(AddRoundKeyOutput[62]), 
        .A2(SubCellInst_LFInst_15_LFInst_0_n4 ), .ZN(
        SubCellInst_LFInst_15_LFInst_0_n5 ) );
  INV_X1 SubCellInst_LFInst_15_LFInst_0_U4  ( .A(AddRoundKeyOutput[61]), .ZN(
        SubCellInst_LFInst_15_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst_LFInst_15_LFInst_0_U3  ( .A(AddRoundKeyOutput[60]), .B(
        AddRoundKeyOutput[63]), .Z(SubCellInst_LFInst_15_LFInst_0_n6 ) );
  XNOR2_X1 MCInst1_MC0_v0_2Inst_0_U4  ( .A(MCInst1_MC0_v0_2Inst_0_n2 ), .B(
        MCInst1_MC0_v0_0 [3]), .ZN(MCInst1_MC0_v0_2 [0]) );
  XNOR2_X1 MCInst1_MC0_v0_2Inst_0_U3  ( .A(MCInst1_MC0_v0_3 [0]), .B(
        ShiftRowsOutput[60]), .ZN(MCInst1_MC0_v0_2Inst_0_n2 ) );
  XOR2_X1 MCInst1_MC0_v1_1Inst_0_U3  ( .A(MCInst1_MC0_v1_3 [3]), .B(
        MCInst1_MC0_v1_3 [0]), .Z(MCInst1_MC0_v1_1 [0]) );
  XNOR2_X1 MCInst1_MC0_v1_2Inst_0_U4  ( .A(MCInst1_MC0_v1_2Inst_0_n2 ), .B(
        MCInst1_MC0_v1_3 [3]), .ZN(MCInst1_MC0_v1_2 [0]) );
  XNOR2_X1 MCInst1_MC0_v1_2Inst_0_U3  ( .A(MCInst1_MC0_v1_3 [0]), .B(
        MCInst1_MC0_v1_3 [2]), .ZN(MCInst1_MC0_v1_2Inst_0_n2 ) );
  XOR2_X1 MCInst1_MC0_v2_1Inst_0_U3  ( .A(MCInst1_MC0_v2_3 [1]), .B(
        MCInst1_MC0_v2_0 [3]), .Z(MCInst1_MC0_v2_1 [0]) );
  XOR2_X1 MCInst1_MC0_v2_2Inst_0_U3  ( .A(MCInst1_MC0_v2_0 [2]), .B(
        MCInst1_MC0_v2_0 [0]), .Z(MCInst1_MC0_v2_2 [0]) );
  XNOR2_X1 MCInst1_MC0_v2_3Inst_0_U5  ( .A(MCInst1_MC0_v2_3Inst_0_n4 ), .B(
        MCInst1_MC0_v2_3Inst_0_n3 ), .ZN(MCInst1_MC0_v2_3 [0]) );
  XNOR2_X1 MCInst1_MC0_v2_3Inst_0_U4  ( .A(MCInst1_MC0_v2_0 [2]), .B(
        MCInst1_MC0_v2_3 [1]), .ZN(MCInst1_MC0_v2_3Inst_0_n3 ) );
  XOR2_X1 MCInst1_MC0_v2_3Inst_0_U3  ( .A(MCInst1_MC0_v2_0 [3]), .B(
        MCInst1_MC0_v2_0 [0]), .Z(MCInst1_MC0_v2_3Inst_0_n4 ) );
  XOR2_X1 MCInst1_MC0_v3_1Inst_0_U3  ( .A(MCInst1_MC0_v3_0 [3]), .B(
        MCInst1_MC0_v3_2 [2]), .Z(MCInst1_MC0_v3_1 [0]) );
  XOR2_X1 MCInst1_MC0_v3_2Inst_0_U3  ( .A(MCInst1_MC0_v3_2 [3]), .B(
        MCInst1_MC0_v3_0 [2]), .Z(MCInst1_MC0_v3_2 [0]) );
  XNOR2_X1 MCInst1_MC0_v3_3Inst_0_U4  ( .A(MCInst1_MC0_v3_3Inst_0_n2 ), .B(
        MCInst1_MC0_v3_0 [2]), .ZN(MCInst1_MC0_v3_3 [0]) );
  XNOR2_X1 MCInst1_MC0_v3_3Inst_0_U3  ( .A(MCInst1_MC0_v3_2 [2]), .B(
        MCInst1_MC0_v3_2 [3]), .ZN(MCInst1_MC0_v3_3Inst_0_n2 ) );
  XOR2_X1 MCInst1_MC0_v0_0Inst_1_U3  ( .A(MCInst1_MC0_v0_3 [3]), .B(
        MCInst1_MC0_v0_3 [0]), .Z(MCInst1_MC0_v0_0 [1]) );
  XOR2_X1 MCInst1_MC0_v0_1Inst_1_U3  ( .A(MCInst1_MC0_v0_0 [3]), .B(
        MCInst1_MC0_v0_3 [3]), .Z(MCInst1_MC0_v0_1 [1]) );
  XNOR2_X1 MCInst1_MC0_v0_2Inst_1_U4  ( .A(MCInst1_MC0_v0_2Inst_1_n2 ), .B(
        MCInst1_MC0_v0_3 [3]), .ZN(MCInst1_MC0_v0_2 [1]) );
  XNOR2_X1 MCInst1_MC0_v0_2Inst_1_U3  ( .A(MCInst1_MC0_v0_3 [0]), .B(
        ShiftRowsOutput[60]), .ZN(MCInst1_MC0_v0_2Inst_1_n2 ) );
  XOR2_X1 MCInst1_MC0_v0_3Inst_1_U3  ( .A(ShiftRowsOutput[60]), .B(
        MCInst1_MC0_v0_3 [0]), .Z(MCInst1_MC0_v0_3 [1]) );
  XOR2_X1 MCInst1_MC0_v1_1Inst_1_U3  ( .A(ShiftRowsOutput[44]), .B(
        MCInst1_MC0_v1_3 [3]), .Z(MCInst1_MC0_v1_1 [1]) );
  XOR2_X1 MCInst1_MC0_v1_2Inst_1_U3  ( .A(ShiftRowsOutput[44]), .B(
        MCInst1_MC0_v1_3 [2]), .Z(MCInst1_MC0_v1_2 [1]) );
  XOR2_X1 MCInst1_MC0_v1_3Inst_1_U3  ( .A(ShiftRowsOutput[44]), .B(
        MCInst1_MC0_v1_3 [0]), .Z(MCInst1_MC0_v1_3 [1]) );
  XOR2_X1 MCInst1_MC0_v2_0Inst_1_U3  ( .A(MCInst1_MC0_v2_3 [1]), .B(
        MCInst1_MC0_v2_0 [0]), .Z(MCInst1_MC0_v2_0 [1]) );
  XNOR2_X1 MCInst1_MC0_v2_1Inst_1_U4  ( .A(MCInst1_MC0_v2_1Inst_1_n2 ), .B(
        MCInst1_MC0_v2_0 [3]), .ZN(MCInst1_MC0_v2_1 [1]) );
  XNOR2_X1 MCInst1_MC0_v2_1Inst_1_U3  ( .A(MCInst1_MC0_v2_0 [0]), .B(
        MCInst1_MC0_v2_0 [2]), .ZN(MCInst1_MC0_v2_1Inst_1_n2 ) );
  XNOR2_X1 MCInst1_MC0_v2_2Inst_1_U5  ( .A(MCInst1_MC0_v2_2Inst_1_n4 ), .B(
        MCInst1_MC0_v2_2Inst_1_n3 ), .ZN(MCInst1_MC0_v2_2 [1]) );
  XNOR2_X1 MCInst1_MC0_v2_2Inst_1_U4  ( .A(MCInst1_MC0_v2_0 [2]), .B(
        MCInst1_MC0_v2_3 [1]), .ZN(MCInst1_MC0_v2_2Inst_1_n3 ) );
  XOR2_X1 MCInst1_MC0_v2_2Inst_1_U3  ( .A(MCInst1_MC0_v2_0 [3]), .B(
        MCInst1_MC0_v2_0 [0]), .Z(MCInst1_MC0_v2_2Inst_1_n4 ) );
  XOR2_X1 MCInst1_MC0_v3_0Inst_1_U3  ( .A(MCInst1_MC0_v3_2 [3]), .B(
        MCInst1_MC0_v3_2 [2]), .Z(MCInst1_MC0_v3_0 [1]) );
  XOR2_X1 MCInst1_MC0_v3_1Inst_1_U3  ( .A(MCInst1_MC0_v3_2 [3]), .B(
        MCInst1_MC0_v3_0 [3]), .Z(MCInst1_MC0_v3_1 [1]) );
  XNOR2_X1 MCInst1_MC0_v3_3Inst_1_U4  ( .A(MCInst1_MC0_v3_3Inst_1_n2 ), .B(
        MCInst1_MC0_v3_0 [3]), .ZN(MCInst1_MC0_v3_3 [1]) );
  XNOR2_X1 MCInst1_MC0_v3_3Inst_1_U3  ( .A(MCInst1_MC0_v3_2 [2]), .B(
        MCInst1_MC0_v3_2 [3]), .ZN(MCInst1_MC0_v3_3Inst_1_n2 ) );
  XOR2_X1 MCInst1_MC0_v0_0Inst_2_U3  ( .A(ShiftRowsOutput[60]), .B(
        MCInst1_MC0_v0_3 [0]), .Z(MCInst1_MC0_v0_0 [2]) );
  XOR2_X1 MCInst1_MC0_v0_1Inst_2_U3  ( .A(MCInst1_MC0_v0_3 [3]), .B(
        MCInst1_MC0_v0_3 [0]), .Z(MCInst1_MC0_v0_1 [2]) );
  XOR2_X1 MCInst1_MC0_v0_2Inst_2_U3  ( .A(MCInst1_MC0_v0_0 [3]), .B(
        MCInst1_MC0_v0_3 [0]), .Z(MCInst1_MC0_v0_2 [2]) );
  XNOR2_X1 MCInst1_MC0_v1_1Inst_2_U4  ( .A(MCInst1_MC0_v1_1Inst_2_n2 ), .B(
        MCInst1_MC0_v1_3 [2]), .ZN(MCInst1_MC0_v1_1 [2]) );
  XNOR2_X1 MCInst1_MC0_v1_1Inst_2_U3  ( .A(MCInst1_MC0_v1_3 [0]), .B(
        ShiftRowsOutput[44]), .ZN(MCInst1_MC0_v1_1Inst_2_n2 ) );
  XNOR2_X1 MCInst1_MC0_v1_2Inst_2_U4  ( .A(MCInst1_MC0_v1_2Inst_2_n2 ), .B(
        MCInst1_MC0_v1_3 [2]), .ZN(MCInst1_MC0_v1_2 [2]) );
  XNOR2_X1 MCInst1_MC0_v1_2Inst_2_U3  ( .A(MCInst1_MC0_v1_3 [3]), .B(
        ShiftRowsOutput[44]), .ZN(MCInst1_MC0_v1_2Inst_2_n2 ) );
  XNOR2_X1 MCInst1_MC0_v2_1Inst_2_U4  ( .A(MCInst1_MC0_v2_1Inst_2_n2 ), .B(
        MCInst1_MC0_v2_0 [3]), .ZN(MCInst1_MC0_v2_1 [2]) );
  XNOR2_X1 MCInst1_MC0_v2_1Inst_2_U3  ( .A(MCInst1_MC0_v2_0 [0]), .B(
        MCInst1_MC0_v2_3 [1]), .ZN(MCInst1_MC0_v2_1Inst_2_n2 ) );
  XNOR2_X1 MCInst1_MC0_v2_2Inst_2_U4  ( .A(MCInst1_MC0_v2_2Inst_2_n2 ), .B(
        MCInst1_MC0_v2_0 [3]), .ZN(MCInst1_MC0_v2_2 [2]) );
  XNOR2_X1 MCInst1_MC0_v2_2Inst_2_U3  ( .A(MCInst1_MC0_v2_0 [0]), .B(
        MCInst1_MC0_v2_0 [2]), .ZN(MCInst1_MC0_v2_2Inst_2_n2 ) );
  XOR2_X1 MCInst1_MC0_v2_3Inst_2_U3  ( .A(MCInst1_MC0_v2_3 [1]), .B(
        MCInst1_MC0_v2_0 [2]), .Z(MCInst1_MC0_v2_3 [2]) );
  XNOR2_X1 MCInst1_MC0_v3_1Inst_2_U4  ( .A(MCInst1_MC0_v3_1Inst_2_n2 ), .B(
        MCInst1_MC0_v3_0 [2]), .ZN(MCInst1_MC0_v3_1 [2]) );
  XNOR2_X1 MCInst1_MC0_v3_1Inst_2_U3  ( .A(MCInst1_MC0_v3_2 [2]), .B(
        MCInst1_MC0_v3_2 [3]), .ZN(MCInst1_MC0_v3_1Inst_2_n2 ) );
  XOR2_X1 MCInst1_MC0_v3_3Inst_2_U3  ( .A(MCInst1_MC0_v3_0 [2]), .B(
        MCInst1_MC0_v3_2 [2]), .Z(MCInst1_MC0_v3_3 [2]) );
  XOR2_X1 MCInst1_MC0_v0_1Inst_3_U3  ( .A(ShiftRowsOutput[60]), .B(
        MCInst1_MC0_v0_3 [0]), .Z(MCInst1_MC0_v0_1 [3]) );
  XOR2_X1 MCInst1_MC0_v0_2Inst_3_U3  ( .A(ShiftRowsOutput[60]), .B(
        MCInst1_MC0_v0_3 [3]), .Z(MCInst1_MC0_v0_2 [3]) );
  XOR2_X1 MCInst1_MC0_v1_1Inst_3_U3  ( .A(MCInst1_MC0_v1_3 [2]), .B(
        MCInst1_MC0_v1_3 [3]), .Z(MCInst1_MC0_v1_1 [3]) );
  XNOR2_X1 MCInst1_MC0_v1_2Inst_3_U5  ( .A(MCInst1_MC0_v1_2Inst_3_n4 ), .B(
        MCInst1_MC0_v1_2Inst_3_n3 ), .ZN(MCInst1_MC0_v1_2 [3]) );
  XNOR2_X1 MCInst1_MC0_v1_2Inst_3_U4  ( .A(MCInst1_MC0_v1_3 [2]), .B(
        ShiftRowsOutput[44]), .ZN(MCInst1_MC0_v1_2Inst_3_n3 ) );
  XOR2_X1 MCInst1_MC0_v1_2Inst_3_U3  ( .A(MCInst1_MC0_v1_3 [3]), .B(
        MCInst1_MC0_v1_3 [0]), .Z(MCInst1_MC0_v1_2Inst_3_n4 ) );
  XOR2_X1 MCInst1_MC0_v2_1Inst_3_U3  ( .A(MCInst1_MC0_v2_0 [2]), .B(
        MCInst1_MC0_v2_0 [0]), .Z(MCInst1_MC0_v2_1 [3]) );
  XNOR2_X1 MCInst1_MC0_v2_2Inst_3_U4  ( .A(MCInst1_MC0_v2_2Inst_3_n2 ), .B(
        MCInst1_MC0_v2_0 [3]), .ZN(MCInst1_MC0_v2_2 [3]) );
  XNOR2_X1 MCInst1_MC0_v2_2Inst_3_U3  ( .A(MCInst1_MC0_v2_0 [0]), .B(
        MCInst1_MC0_v2_3 [1]), .ZN(MCInst1_MC0_v2_2Inst_3_n2 ) );
  XNOR2_X1 MCInst1_MC0_v2_3Inst_3_U4  ( .A(MCInst1_MC0_v2_3Inst_3_n2 ), .B(
        MCInst1_MC0_v2_0 [2]), .ZN(MCInst1_MC0_v2_3 [3]) );
  XNOR2_X1 MCInst1_MC0_v2_3Inst_3_U3  ( .A(MCInst1_MC0_v2_0 [3]), .B(
        MCInst1_MC0_v2_3 [1]), .ZN(MCInst1_MC0_v2_3Inst_3_n2 ) );
  XOR2_X1 MCInst1_MC0_v3_1Inst_3_U3  ( .A(MCInst1_MC0_v3_0 [2]), .B(
        MCInst1_MC0_v3_0 [3]), .Z(MCInst1_MC0_v3_1 [3]) );
  XOR2_X1 MCInst1_MC0_v3_3Inst_3_U3  ( .A(MCInst1_MC0_v3_2 [3]), .B(
        MCInst1_MC0_v3_0 [3]), .Z(MCInst1_MC0_v3_3 [3]) );
  XNOR2_X1 MCInst1_MC0_r0Inst_XORInst_0_0_U3  ( .A(
        MCInst1_MC0_r0Inst_XORInst_0_0_n5 ), .B(
        MCInst1_MC0_r0Inst_XORInst_0_0_n4 ), .ZN(Feedback[60]) );
  XNOR2_X1 MCInst1_MC0_r0Inst_XORInst_0_0_U2  ( .A(MCInst1_MC0_v3_2 [2]), 
        .B(MCInst1_MC0_v2_0 [0]), .ZN(MCInst1_MC0_r0Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst1_MC0_r0Inst_XORInst_0_0_U1  ( .A(MCInst1_MC0_v0_3 [3]), .B(
        ShiftRowsOutput[44]), .Z(MCInst1_MC0_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst1_MC0_r0Inst_XORInst_0_1_U3  ( .A(
        MCInst1_MC0_r0Inst_XORInst_0_1_n5 ), .B(
        MCInst1_MC0_r0Inst_XORInst_0_1_n4 ), .ZN(Feedback[61]) );
  XNOR2_X1 MCInst1_MC0_r0Inst_XORInst_0_1_U2  ( .A(MCInst1_MC0_v3_0 [1]), 
        .B(MCInst1_MC0_v2_0 [1]), .ZN(MCInst1_MC0_r0Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst1_MC0_r0Inst_XORInst_0_1_U1  ( .A(MCInst1_MC0_v0_0 [1]), .B(
        MCInst1_MC0_v1_3 [2]), .Z(MCInst1_MC0_r0Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst1_MC0_r0Inst_XORInst_0_2_U3  ( .A(
        MCInst1_MC0_r0Inst_XORInst_0_2_n5 ), .B(
        MCInst1_MC0_r0Inst_XORInst_0_2_n4 ), .ZN(Feedback[62]) );
  XNOR2_X1 MCInst1_MC0_r0Inst_XORInst_0_2_U2  ( .A(MCInst1_MC0_v3_0 [2]), 
        .B(MCInst1_MC0_v2_0 [2]), .ZN(MCInst1_MC0_r0Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst1_MC0_r0Inst_XORInst_0_2_U1  ( .A(MCInst1_MC0_v0_0 [2]), .B(
        MCInst1_MC0_v1_3 [3]), .Z(MCInst1_MC0_r0Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst1_MC0_r0Inst_XORInst_0_3_U3  ( .A(
        MCInst1_MC0_r0Inst_XORInst_0_3_n5 ), .B(
        MCInst1_MC0_r0Inst_XORInst_0_3_n4 ), .ZN(Feedback[63]) );
  XNOR2_X1 MCInst1_MC0_r0Inst_XORInst_0_3_U2  ( .A(MCInst1_MC0_v3_0 [3]), 
        .B(MCInst1_MC0_v2_0 [3]), .ZN(MCInst1_MC0_r0Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst1_MC0_r0Inst_XORInst_0_3_U1  ( .A(MCInst1_MC0_v0_0 [3]), .B(
        MCInst1_MC0_v1_3 [0]), .Z(MCInst1_MC0_r0Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst1_MC0_r1Inst_XORInst_0_0_U3  ( .A(
        MCInst1_MC0_r1Inst_XORInst_0_0_n5 ), .B(
        MCInst1_MC0_r1Inst_XORInst_0_0_n4 ), .ZN(Feedback[44]) );
  XNOR2_X1 MCInst1_MC0_r1Inst_XORInst_0_0_U2  ( .A(MCInst1_MC0_v3_1 [0]), 
        .B(MCInst1_MC0_v2_1 [0]), .ZN(MCInst1_MC0_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst1_MC0_r1Inst_XORInst_0_0_U1  ( .A(MCInst1_MC0_v0_0 [3]), .B(
        MCInst1_MC0_v1_1 [0]), .Z(MCInst1_MC0_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst1_MC0_r1Inst_XORInst_0_1_U3  ( .A(
        MCInst1_MC0_r1Inst_XORInst_0_1_n5 ), .B(
        MCInst1_MC0_r1Inst_XORInst_0_1_n4 ), .ZN(Feedback[45]) );
  XNOR2_X1 MCInst1_MC0_r1Inst_XORInst_0_1_U2  ( .A(MCInst1_MC0_v3_1 [1]), 
        .B(MCInst1_MC0_v2_1 [1]), .ZN(MCInst1_MC0_r1Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst1_MC0_r1Inst_XORInst_0_1_U1  ( .A(MCInst1_MC0_v0_1 [1]), .B(
        MCInst1_MC0_v1_1 [1]), .Z(MCInst1_MC0_r1Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst1_MC0_r1Inst_XORInst_0_2_U3  ( .A(
        MCInst1_MC0_r1Inst_XORInst_0_2_n5 ), .B(
        MCInst1_MC0_r1Inst_XORInst_0_2_n4 ), .ZN(Feedback[46]) );
  XNOR2_X1 MCInst1_MC0_r1Inst_XORInst_0_2_U2  ( .A(MCInst1_MC0_v3_1 [2]), 
        .B(MCInst1_MC0_v2_1 [2]), .ZN(MCInst1_MC0_r1Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst1_MC0_r1Inst_XORInst_0_2_U1  ( .A(MCInst1_MC0_v0_1 [2]), .B(
        MCInst1_MC0_v1_1 [2]), .Z(MCInst1_MC0_r1Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst1_MC0_r1Inst_XORInst_0_3_U3  ( .A(
        MCInst1_MC0_r1Inst_XORInst_0_3_n5 ), .B(
        MCInst1_MC0_r1Inst_XORInst_0_3_n4 ), .ZN(Feedback[47]) );
  XNOR2_X1 MCInst1_MC0_r1Inst_XORInst_0_3_U2  ( .A(MCInst1_MC0_v3_1 [3]), 
        .B(MCInst1_MC0_v2_1 [3]), .ZN(MCInst1_MC0_r1Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst1_MC0_r1Inst_XORInst_0_3_U1  ( .A(MCInst1_MC0_v0_1 [3]), .B(
        MCInst1_MC0_v1_1 [3]), .Z(MCInst1_MC0_r1Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst1_MC0_r2Inst_XORInst_0_0_U3  ( .A(
        MCInst1_MC0_r2Inst_XORInst_0_0_n5 ), .B(
        MCInst1_MC0_r2Inst_XORInst_0_0_n4 ), .ZN(Feedback[28]) );
  XNOR2_X1 MCInst1_MC0_r2Inst_XORInst_0_0_U2  ( .A(MCInst1_MC0_v3_2 [0]), 
        .B(MCInst1_MC0_v2_2 [0]), .ZN(MCInst1_MC0_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst1_MC0_r2Inst_XORInst_0_0_U1  ( .A(MCInst1_MC0_v0_2 [0]), .B(
        MCInst1_MC0_v1_2 [0]), .Z(MCInst1_MC0_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst1_MC0_r2Inst_XORInst_0_1_U3  ( .A(
        MCInst1_MC0_r2Inst_XORInst_0_1_n5 ), .B(
        MCInst1_MC0_r2Inst_XORInst_0_1_n4 ), .ZN(Feedback[29]) );
  XNOR2_X1 MCInst1_MC0_r2Inst_XORInst_0_1_U2  ( .A(MCInst1_MC0_v3_0 [3]), 
        .B(MCInst1_MC0_v2_2 [1]), .ZN(MCInst1_MC0_r2Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst1_MC0_r2Inst_XORInst_0_1_U1  ( .A(MCInst1_MC0_v0_2 [1]), .B(
        MCInst1_MC0_v1_2 [1]), .Z(MCInst1_MC0_r2Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst1_MC0_r2Inst_XORInst_0_2_U3  ( .A(
        MCInst1_MC0_r2Inst_XORInst_0_2_n5 ), .B(
        MCInst1_MC0_r2Inst_XORInst_0_2_n4 ), .ZN(Feedback[30]) );
  XNOR2_X1 MCInst1_MC0_r2Inst_XORInst_0_2_U2  ( .A(MCInst1_MC0_v3_2 [2]), 
        .B(MCInst1_MC0_v2_2 [2]), .ZN(MCInst1_MC0_r2Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst1_MC0_r2Inst_XORInst_0_2_U1  ( .A(MCInst1_MC0_v0_2 [2]), .B(
        MCInst1_MC0_v1_2 [2]), .Z(MCInst1_MC0_r2Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst1_MC0_r2Inst_XORInst_0_3_U3  ( .A(
        MCInst1_MC0_r2Inst_XORInst_0_3_n5 ), .B(
        MCInst1_MC0_r2Inst_XORInst_0_3_n4 ), .ZN(Feedback[31]) );
  XNOR2_X1 MCInst1_MC0_r2Inst_XORInst_0_3_U2  ( .A(MCInst1_MC0_v3_2 [3]), 
        .B(MCInst1_MC0_v2_2 [3]), .ZN(MCInst1_MC0_r2Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst1_MC0_r2Inst_XORInst_0_3_U1  ( .A(MCInst1_MC0_v0_2 [3]), .B(
        MCInst1_MC0_v1_2 [3]), .Z(MCInst1_MC0_r2Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst1_MC0_r3Inst_XORInst_0_0_U3  ( .A(
        MCInst1_MC0_r3Inst_XORInst_0_0_n5 ), .B(
        MCInst1_MC0_r3Inst_XORInst_0_0_n4 ), .ZN(Feedback[12]) );
  XNOR2_X1 MCInst1_MC0_r3Inst_XORInst_0_0_U2  ( .A(MCInst1_MC0_v3_3 [0]), 
        .B(MCInst1_MC0_v2_3 [0]), .ZN(MCInst1_MC0_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst1_MC0_r3Inst_XORInst_0_0_U1  ( .A(MCInst1_MC0_v0_3 [0]), .B(
        MCInst1_MC0_v1_3 [0]), .Z(MCInst1_MC0_r3Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst1_MC0_r3Inst_XORInst_0_1_U3  ( .A(
        MCInst1_MC0_r3Inst_XORInst_0_1_n5 ), .B(
        MCInst1_MC0_r3Inst_XORInst_0_1_n4 ), .ZN(Feedback[13]) );
  XNOR2_X1 MCInst1_MC0_r3Inst_XORInst_0_1_U2  ( .A(MCInst1_MC0_v3_3 [1]), 
        .B(MCInst1_MC0_v2_3 [1]), .ZN(MCInst1_MC0_r3Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst1_MC0_r3Inst_XORInst_0_1_U1  ( .A(MCInst1_MC0_v0_3 [1]), .B(
        MCInst1_MC0_v1_3 [1]), .Z(MCInst1_MC0_r3Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst1_MC0_r3Inst_XORInst_0_2_U3  ( .A(
        MCInst1_MC0_r3Inst_XORInst_0_2_n5 ), .B(
        MCInst1_MC0_r3Inst_XORInst_0_2_n4 ), .ZN(Feedback[14]) );
  XNOR2_X1 MCInst1_MC0_r3Inst_XORInst_0_2_U2  ( .A(MCInst1_MC0_v3_3 [2]), 
        .B(MCInst1_MC0_v2_3 [2]), .ZN(MCInst1_MC0_r3Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst1_MC0_r3Inst_XORInst_0_2_U1  ( .A(MCInst1_MC0_v0_0 [3]), .B(
        MCInst1_MC0_v1_3 [2]), .Z(MCInst1_MC0_r3Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst1_MC0_r3Inst_XORInst_0_3_U3  ( .A(
        MCInst1_MC0_r3Inst_XORInst_0_3_n5 ), .B(
        MCInst1_MC0_r3Inst_XORInst_0_3_n4 ), .ZN(Feedback[15]) );
  XNOR2_X1 MCInst1_MC0_r3Inst_XORInst_0_3_U2  ( .A(MCInst1_MC0_v3_3 [3]), 
        .B(MCInst1_MC0_v2_3 [3]), .ZN(MCInst1_MC0_r3Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst1_MC0_r3Inst_XORInst_0_3_U1  ( .A(MCInst1_MC0_v0_3 [3]), .B(
        MCInst1_MC0_v1_3 [3]), .Z(MCInst1_MC0_r3Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst1_MC1_v0_2Inst_0_U4  ( .A(MCInst1_MC1_v0_2Inst_0_n2 ), .B(
        MCInst1_MC1_v0_0 [3]), .ZN(MCInst1_MC1_v0_2 [0]) );
  XNOR2_X1 MCInst1_MC1_v0_2Inst_0_U3  ( .A(MCInst1_MC1_v0_3 [0]), .B(
        ShiftRowsOutput[56]), .ZN(MCInst1_MC1_v0_2Inst_0_n2 ) );
  XOR2_X1 MCInst1_MC1_v1_1Inst_0_U3  ( .A(MCInst1_MC1_v1_3 [3]), .B(
        MCInst1_MC1_v1_3 [0]), .Z(MCInst1_MC1_v1_1 [0]) );
  XNOR2_X1 MCInst1_MC1_v1_2Inst_0_U4  ( .A(MCInst1_MC1_v1_2Inst_0_n2 ), .B(
        MCInst1_MC1_v1_3 [3]), .ZN(MCInst1_MC1_v1_2 [0]) );
  XNOR2_X1 MCInst1_MC1_v1_2Inst_0_U3  ( .A(MCInst1_MC1_v1_3 [0]), .B(
        MCInst1_MC1_v1_3 [2]), .ZN(MCInst1_MC1_v1_2Inst_0_n2 ) );
  XOR2_X1 MCInst1_MC1_v2_1Inst_0_U3  ( .A(MCInst1_MC1_v2_3 [1]), .B(
        MCInst1_MC1_v2_0 [3]), .Z(MCInst1_MC1_v2_1 [0]) );
  XOR2_X1 MCInst1_MC1_v2_2Inst_0_U3  ( .A(MCInst1_MC1_v2_0 [2]), .B(
        MCInst1_MC1_v2_0 [0]), .Z(MCInst1_MC1_v2_2 [0]) );
  XNOR2_X1 MCInst1_MC1_v2_3Inst_0_U5  ( .A(MCInst1_MC1_v2_3Inst_0_n4 ), .B(
        MCInst1_MC1_v2_3Inst_0_n3 ), .ZN(MCInst1_MC1_v2_3 [0]) );
  XNOR2_X1 MCInst1_MC1_v2_3Inst_0_U4  ( .A(MCInst1_MC1_v2_0 [2]), .B(
        MCInst1_MC1_v2_3 [1]), .ZN(MCInst1_MC1_v2_3Inst_0_n3 ) );
  XOR2_X1 MCInst1_MC1_v2_3Inst_0_U3  ( .A(MCInst1_MC1_v2_0 [3]), .B(
        MCInst1_MC1_v2_0 [0]), .Z(MCInst1_MC1_v2_3Inst_0_n4 ) );
  XOR2_X1 MCInst1_MC1_v3_1Inst_0_U3  ( .A(MCInst1_MC1_v3_0 [3]), .B(
        MCInst1_MC1_v3_2 [2]), .Z(MCInst1_MC1_v3_1 [0]) );
  XOR2_X1 MCInst1_MC1_v3_2Inst_0_U3  ( .A(MCInst1_MC1_v3_2 [3]), .B(
        MCInst1_MC1_v3_0 [2]), .Z(MCInst1_MC1_v3_2 [0]) );
  XNOR2_X1 MCInst1_MC1_v3_3Inst_0_U4  ( .A(MCInst1_MC1_v3_3Inst_0_n2 ), .B(
        MCInst1_MC1_v3_0 [2]), .ZN(MCInst1_MC1_v3_3 [0]) );
  XNOR2_X1 MCInst1_MC1_v3_3Inst_0_U3  ( .A(MCInst1_MC1_v3_2 [2]), .B(
        MCInst1_MC1_v3_2 [3]), .ZN(MCInst1_MC1_v3_3Inst_0_n2 ) );
  XOR2_X1 MCInst1_MC1_v0_0Inst_1_U3  ( .A(MCInst1_MC1_v0_3 [3]), .B(
        MCInst1_MC1_v0_3 [0]), .Z(MCInst1_MC1_v0_0 [1]) );
  XOR2_X1 MCInst1_MC1_v0_1Inst_1_U3  ( .A(MCInst1_MC1_v0_0 [3]), .B(
        MCInst1_MC1_v0_3 [3]), .Z(MCInst1_MC1_v0_1 [1]) );
  XNOR2_X1 MCInst1_MC1_v0_2Inst_1_U4  ( .A(MCInst1_MC1_v0_2Inst_1_n2 ), .B(
        MCInst1_MC1_v0_3 [3]), .ZN(MCInst1_MC1_v0_2 [1]) );
  XNOR2_X1 MCInst1_MC1_v0_2Inst_1_U3  ( .A(MCInst1_MC1_v0_3 [0]), .B(
        ShiftRowsOutput[56]), .ZN(MCInst1_MC1_v0_2Inst_1_n2 ) );
  XOR2_X1 MCInst1_MC1_v0_3Inst_1_U3  ( .A(ShiftRowsOutput[56]), .B(
        MCInst1_MC1_v0_3 [0]), .Z(MCInst1_MC1_v0_3 [1]) );
  XOR2_X1 MCInst1_MC1_v1_1Inst_1_U3  ( .A(ShiftRowsOutput[40]), .B(
        MCInst1_MC1_v1_3 [3]), .Z(MCInst1_MC1_v1_1 [1]) );
  XOR2_X1 MCInst1_MC1_v1_2Inst_1_U3  ( .A(ShiftRowsOutput[40]), .B(
        MCInst1_MC1_v1_3 [2]), .Z(MCInst1_MC1_v1_2 [1]) );
  XOR2_X1 MCInst1_MC1_v1_3Inst_1_U3  ( .A(ShiftRowsOutput[40]), .B(
        MCInst1_MC1_v1_3 [0]), .Z(MCInst1_MC1_v1_3 [1]) );
  XOR2_X1 MCInst1_MC1_v2_0Inst_1_U3  ( .A(MCInst1_MC1_v2_3 [1]), .B(
        MCInst1_MC1_v2_0 [0]), .Z(MCInst1_MC1_v2_0 [1]) );
  XNOR2_X1 MCInst1_MC1_v2_1Inst_1_U4  ( .A(MCInst1_MC1_v2_1Inst_1_n2 ), .B(
        MCInst1_MC1_v2_0 [3]), .ZN(MCInst1_MC1_v2_1 [1]) );
  XNOR2_X1 MCInst1_MC1_v2_1Inst_1_U3  ( .A(MCInst1_MC1_v2_0 [0]), .B(
        MCInst1_MC1_v2_0 [2]), .ZN(MCInst1_MC1_v2_1Inst_1_n2 ) );
  XNOR2_X1 MCInst1_MC1_v2_2Inst_1_U5  ( .A(MCInst1_MC1_v2_2Inst_1_n4 ), .B(
        MCInst1_MC1_v2_2Inst_1_n3 ), .ZN(MCInst1_MC1_v2_2 [1]) );
  XNOR2_X1 MCInst1_MC1_v2_2Inst_1_U4  ( .A(MCInst1_MC1_v2_0 [2]), .B(
        MCInst1_MC1_v2_3 [1]), .ZN(MCInst1_MC1_v2_2Inst_1_n3 ) );
  XOR2_X1 MCInst1_MC1_v2_2Inst_1_U3  ( .A(MCInst1_MC1_v2_0 [3]), .B(
        MCInst1_MC1_v2_0 [0]), .Z(MCInst1_MC1_v2_2Inst_1_n4 ) );
  XOR2_X1 MCInst1_MC1_v3_0Inst_1_U3  ( .A(MCInst1_MC1_v3_2 [3]), .B(
        MCInst1_MC1_v3_2 [2]), .Z(MCInst1_MC1_v3_0 [1]) );
  XOR2_X1 MCInst1_MC1_v3_1Inst_1_U3  ( .A(MCInst1_MC1_v3_2 [3]), .B(
        MCInst1_MC1_v3_0 [3]), .Z(MCInst1_MC1_v3_1 [1]) );
  XNOR2_X1 MCInst1_MC1_v3_3Inst_1_U4  ( .A(MCInst1_MC1_v3_3Inst_1_n2 ), .B(
        MCInst1_MC1_v3_0 [3]), .ZN(MCInst1_MC1_v3_3 [1]) );
  XNOR2_X1 MCInst1_MC1_v3_3Inst_1_U3  ( .A(MCInst1_MC1_v3_2 [2]), .B(
        MCInst1_MC1_v3_2 [3]), .ZN(MCInst1_MC1_v3_3Inst_1_n2 ) );
  XOR2_X1 MCInst1_MC1_v0_0Inst_2_U3  ( .A(ShiftRowsOutput[56]), .B(
        MCInst1_MC1_v0_3 [0]), .Z(MCInst1_MC1_v0_0 [2]) );
  XOR2_X1 MCInst1_MC1_v0_1Inst_2_U3  ( .A(MCInst1_MC1_v0_3 [3]), .B(
        MCInst1_MC1_v0_3 [0]), .Z(MCInst1_MC1_v0_1 [2]) );
  XOR2_X1 MCInst1_MC1_v0_2Inst_2_U3  ( .A(MCInst1_MC1_v0_0 [3]), .B(
        MCInst1_MC1_v0_3 [0]), .Z(MCInst1_MC1_v0_2 [2]) );
  XNOR2_X1 MCInst1_MC1_v1_1Inst_2_U4  ( .A(MCInst1_MC1_v1_1Inst_2_n2 ), .B(
        MCInst1_MC1_v1_3 [2]), .ZN(MCInst1_MC1_v1_1 [2]) );
  XNOR2_X1 MCInst1_MC1_v1_1Inst_2_U3  ( .A(MCInst1_MC1_v1_3 [0]), .B(
        ShiftRowsOutput[40]), .ZN(MCInst1_MC1_v1_1Inst_2_n2 ) );
  XNOR2_X1 MCInst1_MC1_v1_2Inst_2_U4  ( .A(MCInst1_MC1_v1_2Inst_2_n2 ), .B(
        MCInst1_MC1_v1_3 [2]), .ZN(MCInst1_MC1_v1_2 [2]) );
  XNOR2_X1 MCInst1_MC1_v1_2Inst_2_U3  ( .A(MCInst1_MC1_v1_3 [3]), .B(
        ShiftRowsOutput[40]), .ZN(MCInst1_MC1_v1_2Inst_2_n2 ) );
  XNOR2_X1 MCInst1_MC1_v2_1Inst_2_U4  ( .A(MCInst1_MC1_v2_1Inst_2_n2 ), .B(
        MCInst1_MC1_v2_0 [3]), .ZN(MCInst1_MC1_v2_1 [2]) );
  XNOR2_X1 MCInst1_MC1_v2_1Inst_2_U3  ( .A(MCInst1_MC1_v2_0 [0]), .B(
        MCInst1_MC1_v2_3 [1]), .ZN(MCInst1_MC1_v2_1Inst_2_n2 ) );
  XNOR2_X1 MCInst1_MC1_v2_2Inst_2_U4  ( .A(MCInst1_MC1_v2_2Inst_2_n2 ), .B(
        MCInst1_MC1_v2_0 [3]), .ZN(MCInst1_MC1_v2_2 [2]) );
  XNOR2_X1 MCInst1_MC1_v2_2Inst_2_U3  ( .A(MCInst1_MC1_v2_0 [0]), .B(
        MCInst1_MC1_v2_0 [2]), .ZN(MCInst1_MC1_v2_2Inst_2_n2 ) );
  XOR2_X1 MCInst1_MC1_v2_3Inst_2_U3  ( .A(MCInst1_MC1_v2_3 [1]), .B(
        MCInst1_MC1_v2_0 [2]), .Z(MCInst1_MC1_v2_3 [2]) );
  XNOR2_X1 MCInst1_MC1_v3_1Inst_2_U4  ( .A(MCInst1_MC1_v3_1Inst_2_n2 ), .B(
        MCInst1_MC1_v3_0 [2]), .ZN(MCInst1_MC1_v3_1 [2]) );
  XNOR2_X1 MCInst1_MC1_v3_1Inst_2_U3  ( .A(MCInst1_MC1_v3_2 [2]), .B(
        MCInst1_MC1_v3_2 [3]), .ZN(MCInst1_MC1_v3_1Inst_2_n2 ) );
  XOR2_X1 MCInst1_MC1_v3_3Inst_2_U3  ( .A(MCInst1_MC1_v3_0 [2]), .B(
        MCInst1_MC1_v3_2 [2]), .Z(MCInst1_MC1_v3_3 [2]) );
  XOR2_X1 MCInst1_MC1_v0_1Inst_3_U3  ( .A(ShiftRowsOutput[56]), .B(
        MCInst1_MC1_v0_3 [0]), .Z(MCInst1_MC1_v0_1 [3]) );
  XOR2_X1 MCInst1_MC1_v0_2Inst_3_U3  ( .A(ShiftRowsOutput[56]), .B(
        MCInst1_MC1_v0_3 [3]), .Z(MCInst1_MC1_v0_2 [3]) );
  XOR2_X1 MCInst1_MC1_v1_1Inst_3_U3  ( .A(MCInst1_MC1_v1_3 [2]), .B(
        MCInst1_MC1_v1_3 [3]), .Z(MCInst1_MC1_v1_1 [3]) );
  XNOR2_X1 MCInst1_MC1_v1_2Inst_3_U5  ( .A(MCInst1_MC1_v1_2Inst_3_n4 ), .B(
        MCInst1_MC1_v1_2Inst_3_n3 ), .ZN(MCInst1_MC1_v1_2 [3]) );
  XNOR2_X1 MCInst1_MC1_v1_2Inst_3_U4  ( .A(MCInst1_MC1_v1_3 [2]), .B(
        ShiftRowsOutput[40]), .ZN(MCInst1_MC1_v1_2Inst_3_n3 ) );
  XOR2_X1 MCInst1_MC1_v1_2Inst_3_U3  ( .A(MCInst1_MC1_v1_3 [3]), .B(
        MCInst1_MC1_v1_3 [0]), .Z(MCInst1_MC1_v1_2Inst_3_n4 ) );
  XOR2_X1 MCInst1_MC1_v2_1Inst_3_U3  ( .A(MCInst1_MC1_v2_0 [2]), .B(
        MCInst1_MC1_v2_0 [0]), .Z(MCInst1_MC1_v2_1 [3]) );
  XNOR2_X1 MCInst1_MC1_v2_2Inst_3_U4  ( .A(MCInst1_MC1_v2_2Inst_3_n2 ), .B(
        MCInst1_MC1_v2_0 [3]), .ZN(MCInst1_MC1_v2_2 [3]) );
  XNOR2_X1 MCInst1_MC1_v2_2Inst_3_U3  ( .A(MCInst1_MC1_v2_0 [0]), .B(
        MCInst1_MC1_v2_3 [1]), .ZN(MCInst1_MC1_v2_2Inst_3_n2 ) );
  XNOR2_X1 MCInst1_MC1_v2_3Inst_3_U4  ( .A(MCInst1_MC1_v2_3Inst_3_n2 ), .B(
        MCInst1_MC1_v2_0 [2]), .ZN(MCInst1_MC1_v2_3 [3]) );
  XNOR2_X1 MCInst1_MC1_v2_3Inst_3_U3  ( .A(MCInst1_MC1_v2_0 [3]), .B(
        MCInst1_MC1_v2_3 [1]), .ZN(MCInst1_MC1_v2_3Inst_3_n2 ) );
  XOR2_X1 MCInst1_MC1_v3_1Inst_3_U3  ( .A(MCInst1_MC1_v3_0 [2]), .B(
        MCInst1_MC1_v3_0 [3]), .Z(MCInst1_MC1_v3_1 [3]) );
  XOR2_X1 MCInst1_MC1_v3_3Inst_3_U3  ( .A(MCInst1_MC1_v3_2 [3]), .B(
        MCInst1_MC1_v3_0 [3]), .Z(MCInst1_MC1_v3_3 [3]) );
  XNOR2_X1 MCInst1_MC1_r0Inst_XORInst_0_0_U3  ( .A(
        MCInst1_MC1_r0Inst_XORInst_0_0_n5 ), .B(
        MCInst1_MC1_r0Inst_XORInst_0_0_n4 ), .ZN(Feedback[56]) );
  XNOR2_X1 MCInst1_MC1_r0Inst_XORInst_0_0_U2  ( .A(MCInst1_MC1_v3_2 [2]), 
        .B(MCInst1_MC1_v2_0 [0]), .ZN(MCInst1_MC1_r0Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst1_MC1_r0Inst_XORInst_0_0_U1  ( .A(MCInst1_MC1_v0_3 [3]), .B(
        ShiftRowsOutput[40]), .Z(MCInst1_MC1_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst1_MC1_r0Inst_XORInst_0_1_U3  ( .A(
        MCInst1_MC1_r0Inst_XORInst_0_1_n5 ), .B(
        MCInst1_MC1_r0Inst_XORInst_0_1_n4 ), .ZN(Feedback[57]) );
  XNOR2_X1 MCInst1_MC1_r0Inst_XORInst_0_1_U2  ( .A(MCInst1_MC1_v3_0 [1]), 
        .B(MCInst1_MC1_v2_0 [1]), .ZN(MCInst1_MC1_r0Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst1_MC1_r0Inst_XORInst_0_1_U1  ( .A(MCInst1_MC1_v0_0 [1]), .B(
        MCInst1_MC1_v1_3 [2]), .Z(MCInst1_MC1_r0Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst1_MC1_r0Inst_XORInst_0_2_U3  ( .A(
        MCInst1_MC1_r0Inst_XORInst_0_2_n5 ), .B(
        MCInst1_MC1_r0Inst_XORInst_0_2_n4 ), .ZN(Feedback[58]) );
  XNOR2_X1 MCInst1_MC1_r0Inst_XORInst_0_2_U2  ( .A(MCInst1_MC1_v3_0 [2]), 
        .B(MCInst1_MC1_v2_0 [2]), .ZN(MCInst1_MC1_r0Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst1_MC1_r0Inst_XORInst_0_2_U1  ( .A(MCInst1_MC1_v0_0 [2]), .B(
        MCInst1_MC1_v1_3 [3]), .Z(MCInst1_MC1_r0Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst1_MC1_r0Inst_XORInst_0_3_U3  ( .A(
        MCInst1_MC1_r0Inst_XORInst_0_3_n5 ), .B(
        MCInst1_MC1_r0Inst_XORInst_0_3_n4 ), .ZN(Feedback[59]) );
  XNOR2_X1 MCInst1_MC1_r0Inst_XORInst_0_3_U2  ( .A(MCInst1_MC1_v3_0 [3]), 
        .B(MCInst1_MC1_v2_0 [3]), .ZN(MCInst1_MC1_r0Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst1_MC1_r0Inst_XORInst_0_3_U1  ( .A(MCInst1_MC1_v0_0 [3]), .B(
        MCInst1_MC1_v1_3 [0]), .Z(MCInst1_MC1_r0Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst1_MC1_r1Inst_XORInst_0_0_U3  ( .A(
        MCInst1_MC1_r1Inst_XORInst_0_0_n5 ), .B(
        MCInst1_MC1_r1Inst_XORInst_0_0_n4 ), .ZN(Feedback[40]) );
  XNOR2_X1 MCInst1_MC1_r1Inst_XORInst_0_0_U2  ( .A(MCInst1_MC1_v3_1 [0]), 
        .B(MCInst1_MC1_v2_1 [0]), .ZN(MCInst1_MC1_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst1_MC1_r1Inst_XORInst_0_0_U1  ( .A(MCInst1_MC1_v0_0 [3]), .B(
        MCInst1_MC1_v1_1 [0]), .Z(MCInst1_MC1_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst1_MC1_r1Inst_XORInst_0_1_U3  ( .A(
        MCInst1_MC1_r1Inst_XORInst_0_1_n5 ), .B(
        MCInst1_MC1_r1Inst_XORInst_0_1_n4 ), .ZN(Feedback[41]) );
  XNOR2_X1 MCInst1_MC1_r1Inst_XORInst_0_1_U2  ( .A(MCInst1_MC1_v3_1 [1]), 
        .B(MCInst1_MC1_v2_1 [1]), .ZN(MCInst1_MC1_r1Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst1_MC1_r1Inst_XORInst_0_1_U1  ( .A(MCInst1_MC1_v0_1 [1]), .B(
        MCInst1_MC1_v1_1 [1]), .Z(MCInst1_MC1_r1Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst1_MC1_r1Inst_XORInst_0_2_U3  ( .A(
        MCInst1_MC1_r1Inst_XORInst_0_2_n5 ), .B(
        MCInst1_MC1_r1Inst_XORInst_0_2_n4 ), .ZN(Feedback[42]) );
  XNOR2_X1 MCInst1_MC1_r1Inst_XORInst_0_2_U2  ( .A(MCInst1_MC1_v3_1 [2]), 
        .B(MCInst1_MC1_v2_1 [2]), .ZN(MCInst1_MC1_r1Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst1_MC1_r1Inst_XORInst_0_2_U1  ( .A(MCInst1_MC1_v0_1 [2]), .B(
        MCInst1_MC1_v1_1 [2]), .Z(MCInst1_MC1_r1Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst1_MC1_r1Inst_XORInst_0_3_U3  ( .A(
        MCInst1_MC1_r1Inst_XORInst_0_3_n5 ), .B(
        MCInst1_MC1_r1Inst_XORInst_0_3_n4 ), .ZN(Feedback[43]) );
  XNOR2_X1 MCInst1_MC1_r1Inst_XORInst_0_3_U2  ( .A(MCInst1_MC1_v3_1 [3]), 
        .B(MCInst1_MC1_v2_1 [3]), .ZN(MCInst1_MC1_r1Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst1_MC1_r1Inst_XORInst_0_3_U1  ( .A(MCInst1_MC1_v0_1 [3]), .B(
        MCInst1_MC1_v1_1 [3]), .Z(MCInst1_MC1_r1Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst1_MC1_r2Inst_XORInst_0_0_U3  ( .A(
        MCInst1_MC1_r2Inst_XORInst_0_0_n5 ), .B(
        MCInst1_MC1_r2Inst_XORInst_0_0_n4 ), .ZN(Feedback[24]) );
  XNOR2_X1 MCInst1_MC1_r2Inst_XORInst_0_0_U2  ( .A(MCInst1_MC1_v3_2 [0]), 
        .B(MCInst1_MC1_v2_2 [0]), .ZN(MCInst1_MC1_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst1_MC1_r2Inst_XORInst_0_0_U1  ( .A(MCInst1_MC1_v0_2 [0]), .B(
        MCInst1_MC1_v1_2 [0]), .Z(MCInst1_MC1_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst1_MC1_r2Inst_XORInst_0_1_U3  ( .A(
        MCInst1_MC1_r2Inst_XORInst_0_1_n5 ), .B(
        MCInst1_MC1_r2Inst_XORInst_0_1_n4 ), .ZN(Feedback[25]) );
  XNOR2_X1 MCInst1_MC1_r2Inst_XORInst_0_1_U2  ( .A(MCInst1_MC1_v3_0 [3]), 
        .B(MCInst1_MC1_v2_2 [1]), .ZN(MCInst1_MC1_r2Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst1_MC1_r2Inst_XORInst_0_1_U1  ( .A(MCInst1_MC1_v0_2 [1]), .B(
        MCInst1_MC1_v1_2 [1]), .Z(MCInst1_MC1_r2Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst1_MC1_r2Inst_XORInst_0_2_U3  ( .A(
        MCInst1_MC1_r2Inst_XORInst_0_2_n5 ), .B(
        MCInst1_MC1_r2Inst_XORInst_0_2_n4 ), .ZN(Feedback[26]) );
  XNOR2_X1 MCInst1_MC1_r2Inst_XORInst_0_2_U2  ( .A(MCInst1_MC1_v3_2 [2]), 
        .B(MCInst1_MC1_v2_2 [2]), .ZN(MCInst1_MC1_r2Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst1_MC1_r2Inst_XORInst_0_2_U1  ( .A(MCInst1_MC1_v0_2 [2]), .B(
        MCInst1_MC1_v1_2 [2]), .Z(MCInst1_MC1_r2Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst1_MC1_r2Inst_XORInst_0_3_U3  ( .A(
        MCInst1_MC1_r2Inst_XORInst_0_3_n5 ), .B(
        MCInst1_MC1_r2Inst_XORInst_0_3_n4 ), .ZN(Feedback[27]) );
  XNOR2_X1 MCInst1_MC1_r2Inst_XORInst_0_3_U2  ( .A(MCInst1_MC1_v3_2 [3]), 
        .B(MCInst1_MC1_v2_2 [3]), .ZN(MCInst1_MC1_r2Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst1_MC1_r2Inst_XORInst_0_3_U1  ( .A(MCInst1_MC1_v0_2 [3]), .B(
        MCInst1_MC1_v1_2 [3]), .Z(MCInst1_MC1_r2Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst1_MC1_r3Inst_XORInst_0_0_U3  ( .A(
        MCInst1_MC1_r3Inst_XORInst_0_0_n5 ), .B(
        MCInst1_MC1_r3Inst_XORInst_0_0_n4 ), .ZN(Feedback[8]) );
  XNOR2_X1 MCInst1_MC1_r3Inst_XORInst_0_0_U2  ( .A(MCInst1_MC1_v3_3 [0]), 
        .B(MCInst1_MC1_v2_3 [0]), .ZN(MCInst1_MC1_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst1_MC1_r3Inst_XORInst_0_0_U1  ( .A(MCInst1_MC1_v0_3 [0]), .B(
        MCInst1_MC1_v1_3 [0]), .Z(MCInst1_MC1_r3Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst1_MC1_r3Inst_XORInst_0_1_U3  ( .A(
        MCInst1_MC1_r3Inst_XORInst_0_1_n5 ), .B(
        MCInst1_MC1_r3Inst_XORInst_0_1_n4 ), .ZN(Feedback[9]) );
  XNOR2_X1 MCInst1_MC1_r3Inst_XORInst_0_1_U2  ( .A(MCInst1_MC1_v3_3 [1]), 
        .B(MCInst1_MC1_v2_3 [1]), .ZN(MCInst1_MC1_r3Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst1_MC1_r3Inst_XORInst_0_1_U1  ( .A(MCInst1_MC1_v0_3 [1]), .B(
        MCInst1_MC1_v1_3 [1]), .Z(MCInst1_MC1_r3Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst1_MC1_r3Inst_XORInst_0_2_U3  ( .A(
        MCInst1_MC1_r3Inst_XORInst_0_2_n5 ), .B(
        MCInst1_MC1_r3Inst_XORInst_0_2_n4 ), .ZN(Feedback[10]) );
  XNOR2_X1 MCInst1_MC1_r3Inst_XORInst_0_2_U2  ( .A(MCInst1_MC1_v3_3 [2]), 
        .B(MCInst1_MC1_v2_3 [2]), .ZN(MCInst1_MC1_r3Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst1_MC1_r3Inst_XORInst_0_2_U1  ( .A(MCInst1_MC1_v0_0 [3]), .B(
        MCInst1_MC1_v1_3 [2]), .Z(MCInst1_MC1_r3Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst1_MC1_r3Inst_XORInst_0_3_U3  ( .A(
        MCInst1_MC1_r3Inst_XORInst_0_3_n5 ), .B(
        MCInst1_MC1_r3Inst_XORInst_0_3_n4 ), .ZN(Feedback[11]) );
  XNOR2_X1 MCInst1_MC1_r3Inst_XORInst_0_3_U2  ( .A(MCInst1_MC1_v3_3 [3]), 
        .B(MCInst1_MC1_v2_3 [3]), .ZN(MCInst1_MC1_r3Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst1_MC1_r3Inst_XORInst_0_3_U1  ( .A(MCInst1_MC1_v0_3 [3]), .B(
        MCInst1_MC1_v1_3 [3]), .Z(MCInst1_MC1_r3Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst1_MC2_v0_2Inst_0_U4  ( .A(MCInst1_MC2_v0_2Inst_0_n2 ), .B(
        MCInst1_MC2_v0_0 [3]), .ZN(MCInst1_MC2_v0_2 [0]) );
  XNOR2_X1 MCInst1_MC2_v0_2Inst_0_U3  ( .A(MCInst1_MC2_v0_3 [0]), .B(
        ShiftRowsOutput[52]), .ZN(MCInst1_MC2_v0_2Inst_0_n2 ) );
  XOR2_X1 MCInst1_MC2_v1_1Inst_0_U3  ( .A(MCInst1_MC2_v1_3 [3]), .B(
        MCInst1_MC2_v1_3 [0]), .Z(MCInst1_MC2_v1_1 [0]) );
  XNOR2_X1 MCInst1_MC2_v1_2Inst_0_U4  ( .A(MCInst1_MC2_v1_2Inst_0_n2 ), .B(
        MCInst1_MC2_v1_3 [3]), .ZN(MCInst1_MC2_v1_2 [0]) );
  XNOR2_X1 MCInst1_MC2_v1_2Inst_0_U3  ( .A(MCInst1_MC2_v1_3 [0]), .B(
        MCInst1_MC2_v1_3 [2]), .ZN(MCInst1_MC2_v1_2Inst_0_n2 ) );
  XOR2_X1 MCInst1_MC2_v2_1Inst_0_U3  ( .A(MCInst1_MC2_v2_3 [1]), .B(
        MCInst1_MC2_v2_0 [3]), .Z(MCInst1_MC2_v2_1 [0]) );
  XOR2_X1 MCInst1_MC2_v2_2Inst_0_U3  ( .A(MCInst1_MC2_v2_0 [2]), .B(
        MCInst1_MC2_v2_0 [0]), .Z(MCInst1_MC2_v2_2 [0]) );
  XNOR2_X1 MCInst1_MC2_v2_3Inst_0_U5  ( .A(MCInst1_MC2_v2_3Inst_0_n4 ), .B(
        MCInst1_MC2_v2_3Inst_0_n3 ), .ZN(MCInst1_MC2_v2_3 [0]) );
  XNOR2_X1 MCInst1_MC2_v2_3Inst_0_U4  ( .A(MCInst1_MC2_v2_0 [2]), .B(
        MCInst1_MC2_v2_3 [1]), .ZN(MCInst1_MC2_v2_3Inst_0_n3 ) );
  XOR2_X1 MCInst1_MC2_v2_3Inst_0_U3  ( .A(MCInst1_MC2_v2_0 [3]), .B(
        MCInst1_MC2_v2_0 [0]), .Z(MCInst1_MC2_v2_3Inst_0_n4 ) );
  XOR2_X1 MCInst1_MC2_v3_1Inst_0_U3  ( .A(MCInst1_MC2_v3_0 [3]), .B(
        MCInst1_MC2_v3_2 [2]), .Z(MCInst1_MC2_v3_1 [0]) );
  XOR2_X1 MCInst1_MC2_v3_2Inst_0_U3  ( .A(MCInst1_MC2_v3_2 [3]), .B(
        MCInst1_MC2_v3_0 [2]), .Z(MCInst1_MC2_v3_2 [0]) );
  XNOR2_X1 MCInst1_MC2_v3_3Inst_0_U4  ( .A(MCInst1_MC2_v3_3Inst_0_n2 ), .B(
        MCInst1_MC2_v3_0 [2]), .ZN(MCInst1_MC2_v3_3 [0]) );
  XNOR2_X1 MCInst1_MC2_v3_3Inst_0_U3  ( .A(MCInst1_MC2_v3_2 [2]), .B(
        MCInst1_MC2_v3_2 [3]), .ZN(MCInst1_MC2_v3_3Inst_0_n2 ) );
  XOR2_X1 MCInst1_MC2_v0_0Inst_1_U3  ( .A(MCInst1_MC2_v0_3 [3]), .B(
        MCInst1_MC2_v0_3 [0]), .Z(MCInst1_MC2_v0_0 [1]) );
  XOR2_X1 MCInst1_MC2_v0_1Inst_1_U3  ( .A(MCInst1_MC2_v0_0 [3]), .B(
        MCInst1_MC2_v0_3 [3]), .Z(MCInst1_MC2_v0_1 [1]) );
  XNOR2_X1 MCInst1_MC2_v0_2Inst_1_U4  ( .A(MCInst1_MC2_v0_2Inst_1_n2 ), .B(
        MCInst1_MC2_v0_3 [3]), .ZN(MCInst1_MC2_v0_2 [1]) );
  XNOR2_X1 MCInst1_MC2_v0_2Inst_1_U3  ( .A(MCInst1_MC2_v0_3 [0]), .B(
        ShiftRowsOutput[52]), .ZN(MCInst1_MC2_v0_2Inst_1_n2 ) );
  XOR2_X1 MCInst1_MC2_v0_3Inst_1_U3  ( .A(ShiftRowsOutput[52]), .B(
        MCInst1_MC2_v0_3 [0]), .Z(MCInst1_MC2_v0_3 [1]) );
  XOR2_X1 MCInst1_MC2_v1_1Inst_1_U3  ( .A(ShiftRowsOutput[36]), .B(
        MCInst1_MC2_v1_3 [3]), .Z(MCInst1_MC2_v1_1 [1]) );
  XOR2_X1 MCInst1_MC2_v1_2Inst_1_U3  ( .A(ShiftRowsOutput[36]), .B(
        MCInst1_MC2_v1_3 [2]), .Z(MCInst1_MC2_v1_2 [1]) );
  XOR2_X1 MCInst1_MC2_v1_3Inst_1_U3  ( .A(ShiftRowsOutput[36]), .B(
        MCInst1_MC2_v1_3 [0]), .Z(MCInst1_MC2_v1_3 [1]) );
  XOR2_X1 MCInst1_MC2_v2_0Inst_1_U3  ( .A(MCInst1_MC2_v2_3 [1]), .B(
        MCInst1_MC2_v2_0 [0]), .Z(MCInst1_MC2_v2_0 [1]) );
  XNOR2_X1 MCInst1_MC2_v2_1Inst_1_U4  ( .A(MCInst1_MC2_v2_1Inst_1_n2 ), .B(
        MCInst1_MC2_v2_0 [3]), .ZN(MCInst1_MC2_v2_1 [1]) );
  XNOR2_X1 MCInst1_MC2_v2_1Inst_1_U3  ( .A(MCInst1_MC2_v2_0 [0]), .B(
        MCInst1_MC2_v2_0 [2]), .ZN(MCInst1_MC2_v2_1Inst_1_n2 ) );
  XNOR2_X1 MCInst1_MC2_v2_2Inst_1_U5  ( .A(MCInst1_MC2_v2_2Inst_1_n4 ), .B(
        MCInst1_MC2_v2_2Inst_1_n3 ), .ZN(MCInst1_MC2_v2_2 [1]) );
  XNOR2_X1 MCInst1_MC2_v2_2Inst_1_U4  ( .A(MCInst1_MC2_v2_0 [2]), .B(
        MCInst1_MC2_v2_3 [1]), .ZN(MCInst1_MC2_v2_2Inst_1_n3 ) );
  XOR2_X1 MCInst1_MC2_v2_2Inst_1_U3  ( .A(MCInst1_MC2_v2_0 [3]), .B(
        MCInst1_MC2_v2_0 [0]), .Z(MCInst1_MC2_v2_2Inst_1_n4 ) );
  XOR2_X1 MCInst1_MC2_v3_0Inst_1_U3  ( .A(MCInst1_MC2_v3_2 [3]), .B(
        MCInst1_MC2_v3_2 [2]), .Z(MCInst1_MC2_v3_0 [1]) );
  XOR2_X1 MCInst1_MC2_v3_1Inst_1_U3  ( .A(MCInst1_MC2_v3_2 [3]), .B(
        MCInst1_MC2_v3_0 [3]), .Z(MCInst1_MC2_v3_1 [1]) );
  XNOR2_X1 MCInst1_MC2_v3_3Inst_1_U4  ( .A(MCInst1_MC2_v3_3Inst_1_n2 ), .B(
        MCInst1_MC2_v3_0 [3]), .ZN(MCInst1_MC2_v3_3 [1]) );
  XNOR2_X1 MCInst1_MC2_v3_3Inst_1_U3  ( .A(MCInst1_MC2_v3_2 [2]), .B(
        MCInst1_MC2_v3_2 [3]), .ZN(MCInst1_MC2_v3_3Inst_1_n2 ) );
  XOR2_X1 MCInst1_MC2_v0_0Inst_2_U3  ( .A(ShiftRowsOutput[52]), .B(
        MCInst1_MC2_v0_3 [0]), .Z(MCInst1_MC2_v0_0 [2]) );
  XOR2_X1 MCInst1_MC2_v0_1Inst_2_U3  ( .A(MCInst1_MC2_v0_3 [3]), .B(
        MCInst1_MC2_v0_3 [0]), .Z(MCInst1_MC2_v0_1 [2]) );
  XOR2_X1 MCInst1_MC2_v0_2Inst_2_U3  ( .A(MCInst1_MC2_v0_0 [3]), .B(
        MCInst1_MC2_v0_3 [0]), .Z(MCInst1_MC2_v0_2 [2]) );
  XNOR2_X1 MCInst1_MC2_v1_1Inst_2_U4  ( .A(MCInst1_MC2_v1_1Inst_2_n2 ), .B(
        MCInst1_MC2_v1_3 [2]), .ZN(MCInst1_MC2_v1_1 [2]) );
  XNOR2_X1 MCInst1_MC2_v1_1Inst_2_U3  ( .A(MCInst1_MC2_v1_3 [0]), .B(
        ShiftRowsOutput[36]), .ZN(MCInst1_MC2_v1_1Inst_2_n2 ) );
  XNOR2_X1 MCInst1_MC2_v1_2Inst_2_U4  ( .A(MCInst1_MC2_v1_2Inst_2_n2 ), .B(
        MCInst1_MC2_v1_3 [2]), .ZN(MCInst1_MC2_v1_2 [2]) );
  XNOR2_X1 MCInst1_MC2_v1_2Inst_2_U3  ( .A(MCInst1_MC2_v1_3 [3]), .B(
        ShiftRowsOutput[36]), .ZN(MCInst1_MC2_v1_2Inst_2_n2 ) );
  XNOR2_X1 MCInst1_MC2_v2_1Inst_2_U4  ( .A(MCInst1_MC2_v2_1Inst_2_n2 ), .B(
        MCInst1_MC2_v2_0 [3]), .ZN(MCInst1_MC2_v2_1 [2]) );
  XNOR2_X1 MCInst1_MC2_v2_1Inst_2_U3  ( .A(MCInst1_MC2_v2_0 [0]), .B(
        MCInst1_MC2_v2_3 [1]), .ZN(MCInst1_MC2_v2_1Inst_2_n2 ) );
  XNOR2_X1 MCInst1_MC2_v2_2Inst_2_U4  ( .A(MCInst1_MC2_v2_2Inst_2_n2 ), .B(
        MCInst1_MC2_v2_0 [3]), .ZN(MCInst1_MC2_v2_2 [2]) );
  XNOR2_X1 MCInst1_MC2_v2_2Inst_2_U3  ( .A(MCInst1_MC2_v2_0 [0]), .B(
        MCInst1_MC2_v2_0 [2]), .ZN(MCInst1_MC2_v2_2Inst_2_n2 ) );
  XOR2_X1 MCInst1_MC2_v2_3Inst_2_U3  ( .A(MCInst1_MC2_v2_3 [1]), .B(
        MCInst1_MC2_v2_0 [2]), .Z(MCInst1_MC2_v2_3 [2]) );
  XNOR2_X1 MCInst1_MC2_v3_1Inst_2_U4  ( .A(MCInst1_MC2_v3_1Inst_2_n2 ), .B(
        MCInst1_MC2_v3_0 [2]), .ZN(MCInst1_MC2_v3_1 [2]) );
  XNOR2_X1 MCInst1_MC2_v3_1Inst_2_U3  ( .A(MCInst1_MC2_v3_2 [2]), .B(
        MCInst1_MC2_v3_2 [3]), .ZN(MCInst1_MC2_v3_1Inst_2_n2 ) );
  XOR2_X1 MCInst1_MC2_v3_3Inst_2_U3  ( .A(MCInst1_MC2_v3_0 [2]), .B(
        MCInst1_MC2_v3_2 [2]), .Z(MCInst1_MC2_v3_3 [2]) );
  XOR2_X1 MCInst1_MC2_v0_1Inst_3_U3  ( .A(ShiftRowsOutput[52]), .B(
        MCInst1_MC2_v0_3 [0]), .Z(MCInst1_MC2_v0_1 [3]) );
  XOR2_X1 MCInst1_MC2_v0_2Inst_3_U3  ( .A(ShiftRowsOutput[52]), .B(
        MCInst1_MC2_v0_3 [3]), .Z(MCInst1_MC2_v0_2 [3]) );
  XOR2_X1 MCInst1_MC2_v1_1Inst_3_U3  ( .A(MCInst1_MC2_v1_3 [2]), .B(
        MCInst1_MC2_v1_3 [3]), .Z(MCInst1_MC2_v1_1 [3]) );
  XNOR2_X1 MCInst1_MC2_v1_2Inst_3_U5  ( .A(MCInst1_MC2_v1_2Inst_3_n4 ), .B(
        MCInst1_MC2_v1_2Inst_3_n3 ), .ZN(MCInst1_MC2_v1_2 [3]) );
  XNOR2_X1 MCInst1_MC2_v1_2Inst_3_U4  ( .A(MCInst1_MC2_v1_3 [2]), .B(
        ShiftRowsOutput[36]), .ZN(MCInst1_MC2_v1_2Inst_3_n3 ) );
  XOR2_X1 MCInst1_MC2_v1_2Inst_3_U3  ( .A(MCInst1_MC2_v1_3 [3]), .B(
        MCInst1_MC2_v1_3 [0]), .Z(MCInst1_MC2_v1_2Inst_3_n4 ) );
  XOR2_X1 MCInst1_MC2_v2_1Inst_3_U3  ( .A(MCInst1_MC2_v2_0 [2]), .B(
        MCInst1_MC2_v2_0 [0]), .Z(MCInst1_MC2_v2_1 [3]) );
  XNOR2_X1 MCInst1_MC2_v2_2Inst_3_U4  ( .A(MCInst1_MC2_v2_2Inst_3_n2 ), .B(
        MCInst1_MC2_v2_0 [3]), .ZN(MCInst1_MC2_v2_2 [3]) );
  XNOR2_X1 MCInst1_MC2_v2_2Inst_3_U3  ( .A(MCInst1_MC2_v2_0 [0]), .B(
        MCInst1_MC2_v2_3 [1]), .ZN(MCInst1_MC2_v2_2Inst_3_n2 ) );
  XNOR2_X1 MCInst1_MC2_v2_3Inst_3_U4  ( .A(MCInst1_MC2_v2_3Inst_3_n2 ), .B(
        MCInst1_MC2_v2_0 [2]), .ZN(MCInst1_MC2_v2_3 [3]) );
  XNOR2_X1 MCInst1_MC2_v2_3Inst_3_U3  ( .A(MCInst1_MC2_v2_0 [3]), .B(
        MCInst1_MC2_v2_3 [1]), .ZN(MCInst1_MC2_v2_3Inst_3_n2 ) );
  XOR2_X1 MCInst1_MC2_v3_1Inst_3_U3  ( .A(MCInst1_MC2_v3_0 [2]), .B(
        MCInst1_MC2_v3_0 [3]), .Z(MCInst1_MC2_v3_1 [3]) );
  XOR2_X1 MCInst1_MC2_v3_3Inst_3_U3  ( .A(MCInst1_MC2_v3_2 [3]), .B(
        MCInst1_MC2_v3_0 [3]), .Z(MCInst1_MC2_v3_3 [3]) );
  XNOR2_X1 MCInst1_MC2_r0Inst_XORInst_0_0_U3  ( .A(
        MCInst1_MC2_r0Inst_XORInst_0_0_n5 ), .B(
        MCInst1_MC2_r0Inst_XORInst_0_0_n4 ), .ZN(Feedback[52]) );
  XNOR2_X1 MCInst1_MC2_r0Inst_XORInst_0_0_U2  ( .A(MCInst1_MC2_v3_2 [2]), 
        .B(MCInst1_MC2_v2_0 [0]), .ZN(MCInst1_MC2_r0Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst1_MC2_r0Inst_XORInst_0_0_U1  ( .A(MCInst1_MC2_v0_3 [3]), .B(
        ShiftRowsOutput[36]), .Z(MCInst1_MC2_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst1_MC2_r0Inst_XORInst_0_1_U3  ( .A(
        MCInst1_MC2_r0Inst_XORInst_0_1_n5 ), .B(
        MCInst1_MC2_r0Inst_XORInst_0_1_n4 ), .ZN(Feedback[53]) );
  XNOR2_X1 MCInst1_MC2_r0Inst_XORInst_0_1_U2  ( .A(MCInst1_MC2_v3_0 [1]), 
        .B(MCInst1_MC2_v2_0 [1]), .ZN(MCInst1_MC2_r0Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst1_MC2_r0Inst_XORInst_0_1_U1  ( .A(MCInst1_MC2_v0_0 [1]), .B(
        MCInst1_MC2_v1_3 [2]), .Z(MCInst1_MC2_r0Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst1_MC2_r0Inst_XORInst_0_2_U3  ( .A(
        MCInst1_MC2_r0Inst_XORInst_0_2_n5 ), .B(
        MCInst1_MC2_r0Inst_XORInst_0_2_n4 ), .ZN(Feedback[54]) );
  XNOR2_X1 MCInst1_MC2_r0Inst_XORInst_0_2_U2  ( .A(MCInst1_MC2_v3_0 [2]), 
        .B(MCInst1_MC2_v2_0 [2]), .ZN(MCInst1_MC2_r0Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst1_MC2_r0Inst_XORInst_0_2_U1  ( .A(MCInst1_MC2_v0_0 [2]), .B(
        MCInst1_MC2_v1_3 [3]), .Z(MCInst1_MC2_r0Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst1_MC2_r0Inst_XORInst_0_3_U3  ( .A(
        MCInst1_MC2_r0Inst_XORInst_0_3_n5 ), .B(
        MCInst1_MC2_r0Inst_XORInst_0_3_n4 ), .ZN(Feedback[55]) );
  XNOR2_X1 MCInst1_MC2_r0Inst_XORInst_0_3_U2  ( .A(MCInst1_MC2_v3_0 [3]), 
        .B(MCInst1_MC2_v2_0 [3]), .ZN(MCInst1_MC2_r0Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst1_MC2_r0Inst_XORInst_0_3_U1  ( .A(MCInst1_MC2_v0_0 [3]), .B(
        MCInst1_MC2_v1_3 [0]), .Z(MCInst1_MC2_r0Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst1_MC2_r1Inst_XORInst_0_0_U3  ( .A(
        MCInst1_MC2_r1Inst_XORInst_0_0_n5 ), .B(
        MCInst1_MC2_r1Inst_XORInst_0_0_n4 ), .ZN(Feedback[36]) );
  XNOR2_X1 MCInst1_MC2_r1Inst_XORInst_0_0_U2  ( .A(MCInst1_MC2_v3_1 [0]), 
        .B(MCInst1_MC2_v2_1 [0]), .ZN(MCInst1_MC2_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst1_MC2_r1Inst_XORInst_0_0_U1  ( .A(MCInst1_MC2_v0_0 [3]), .B(
        MCInst1_MC2_v1_1 [0]), .Z(MCInst1_MC2_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst1_MC2_r1Inst_XORInst_0_1_U3  ( .A(
        MCInst1_MC2_r1Inst_XORInst_0_1_n5 ), .B(
        MCInst1_MC2_r1Inst_XORInst_0_1_n4 ), .ZN(Feedback[37]) );
  XNOR2_X1 MCInst1_MC2_r1Inst_XORInst_0_1_U2  ( .A(MCInst1_MC2_v3_1 [1]), 
        .B(MCInst1_MC2_v2_1 [1]), .ZN(MCInst1_MC2_r1Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst1_MC2_r1Inst_XORInst_0_1_U1  ( .A(MCInst1_MC2_v0_1 [1]), .B(
        MCInst1_MC2_v1_1 [1]), .Z(MCInst1_MC2_r1Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst1_MC2_r1Inst_XORInst_0_2_U3  ( .A(
        MCInst1_MC2_r1Inst_XORInst_0_2_n5 ), .B(
        MCInst1_MC2_r1Inst_XORInst_0_2_n4 ), .ZN(Feedback[38]) );
  XNOR2_X1 MCInst1_MC2_r1Inst_XORInst_0_2_U2  ( .A(MCInst1_MC2_v3_1 [2]), 
        .B(MCInst1_MC2_v2_1 [2]), .ZN(MCInst1_MC2_r1Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst1_MC2_r1Inst_XORInst_0_2_U1  ( .A(MCInst1_MC2_v0_1 [2]), .B(
        MCInst1_MC2_v1_1 [2]), .Z(MCInst1_MC2_r1Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst1_MC2_r1Inst_XORInst_0_3_U3  ( .A(
        MCInst1_MC2_r1Inst_XORInst_0_3_n5 ), .B(
        MCInst1_MC2_r1Inst_XORInst_0_3_n4 ), .ZN(Feedback[39]) );
  XNOR2_X1 MCInst1_MC2_r1Inst_XORInst_0_3_U2  ( .A(MCInst1_MC2_v3_1 [3]), 
        .B(MCInst1_MC2_v2_1 [3]), .ZN(MCInst1_MC2_r1Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst1_MC2_r1Inst_XORInst_0_3_U1  ( .A(MCInst1_MC2_v0_1 [3]), .B(
        MCInst1_MC2_v1_1 [3]), .Z(MCInst1_MC2_r1Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst1_MC2_r2Inst_XORInst_0_0_U3  ( .A(
        MCInst1_MC2_r2Inst_XORInst_0_0_n5 ), .B(
        MCInst1_MC2_r2Inst_XORInst_0_0_n4 ), .ZN(Feedback[20]) );
  XNOR2_X1 MCInst1_MC2_r2Inst_XORInst_0_0_U2  ( .A(MCInst1_MC2_v3_2 [0]), 
        .B(MCInst1_MC2_v2_2 [0]), .ZN(MCInst1_MC2_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst1_MC2_r2Inst_XORInst_0_0_U1  ( .A(MCInst1_MC2_v0_2 [0]), .B(
        MCInst1_MC2_v1_2 [0]), .Z(MCInst1_MC2_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst1_MC2_r2Inst_XORInst_0_1_U3  ( .A(
        MCInst1_MC2_r2Inst_XORInst_0_1_n5 ), .B(
        MCInst1_MC2_r2Inst_XORInst_0_1_n4 ), .ZN(Feedback[21]) );
  XNOR2_X1 MCInst1_MC2_r2Inst_XORInst_0_1_U2  ( .A(MCInst1_MC2_v3_0 [3]), 
        .B(MCInst1_MC2_v2_2 [1]), .ZN(MCInst1_MC2_r2Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst1_MC2_r2Inst_XORInst_0_1_U1  ( .A(MCInst1_MC2_v0_2 [1]), .B(
        MCInst1_MC2_v1_2 [1]), .Z(MCInst1_MC2_r2Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst1_MC2_r2Inst_XORInst_0_2_U3  ( .A(
        MCInst1_MC2_r2Inst_XORInst_0_2_n5 ), .B(
        MCInst1_MC2_r2Inst_XORInst_0_2_n4 ), .ZN(Feedback[22]) );
  XNOR2_X1 MCInst1_MC2_r2Inst_XORInst_0_2_U2  ( .A(MCInst1_MC2_v3_2 [2]), 
        .B(MCInst1_MC2_v2_2 [2]), .ZN(MCInst1_MC2_r2Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst1_MC2_r2Inst_XORInst_0_2_U1  ( .A(MCInst1_MC2_v0_2 [2]), .B(
        MCInst1_MC2_v1_2 [2]), .Z(MCInst1_MC2_r2Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst1_MC2_r2Inst_XORInst_0_3_U3  ( .A(
        MCInst1_MC2_r2Inst_XORInst_0_3_n5 ), .B(
        MCInst1_MC2_r2Inst_XORInst_0_3_n4 ), .ZN(Feedback[23]) );
  XNOR2_X1 MCInst1_MC2_r2Inst_XORInst_0_3_U2  ( .A(MCInst1_MC2_v3_2 [3]), 
        .B(MCInst1_MC2_v2_2 [3]), .ZN(MCInst1_MC2_r2Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst1_MC2_r2Inst_XORInst_0_3_U1  ( .A(MCInst1_MC2_v0_2 [3]), .B(
        MCInst1_MC2_v1_2 [3]), .Z(MCInst1_MC2_r2Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst1_MC2_r3Inst_XORInst_0_0_U3  ( .A(
        MCInst1_MC2_r3Inst_XORInst_0_0_n5 ), .B(
        MCInst1_MC2_r3Inst_XORInst_0_0_n4 ), .ZN(Feedback[4]) );
  XNOR2_X1 MCInst1_MC2_r3Inst_XORInst_0_0_U2  ( .A(MCInst1_MC2_v3_3 [0]), 
        .B(MCInst1_MC2_v2_3 [0]), .ZN(MCInst1_MC2_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst1_MC2_r3Inst_XORInst_0_0_U1  ( .A(MCInst1_MC2_v0_3 [0]), .B(
        MCInst1_MC2_v1_3 [0]), .Z(MCInst1_MC2_r3Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst1_MC2_r3Inst_XORInst_0_1_U3  ( .A(
        MCInst1_MC2_r3Inst_XORInst_0_1_n5 ), .B(
        MCInst1_MC2_r3Inst_XORInst_0_1_n4 ), .ZN(Feedback[5]) );
  XNOR2_X1 MCInst1_MC2_r3Inst_XORInst_0_1_U2  ( .A(MCInst1_MC2_v3_3 [1]), 
        .B(MCInst1_MC2_v2_3 [1]), .ZN(MCInst1_MC2_r3Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst1_MC2_r3Inst_XORInst_0_1_U1  ( .A(MCInst1_MC2_v0_3 [1]), .B(
        MCInst1_MC2_v1_3 [1]), .Z(MCInst1_MC2_r3Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst1_MC2_r3Inst_XORInst_0_2_U3  ( .A(
        MCInst1_MC2_r3Inst_XORInst_0_2_n5 ), .B(
        MCInst1_MC2_r3Inst_XORInst_0_2_n4 ), .ZN(Feedback[6]) );
  XNOR2_X1 MCInst1_MC2_r3Inst_XORInst_0_2_U2  ( .A(MCInst1_MC2_v3_3 [2]), 
        .B(MCInst1_MC2_v2_3 [2]), .ZN(MCInst1_MC2_r3Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst1_MC2_r3Inst_XORInst_0_2_U1  ( .A(MCInst1_MC2_v0_0 [3]), .B(
        MCInst1_MC2_v1_3 [2]), .Z(MCInst1_MC2_r3Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst1_MC2_r3Inst_XORInst_0_3_U3  ( .A(
        MCInst1_MC2_r3Inst_XORInst_0_3_n5 ), .B(
        MCInst1_MC2_r3Inst_XORInst_0_3_n4 ), .ZN(Feedback[7]) );
  XNOR2_X1 MCInst1_MC2_r3Inst_XORInst_0_3_U2  ( .A(MCInst1_MC2_v3_3 [3]), 
        .B(MCInst1_MC2_v2_3 [3]), .ZN(MCInst1_MC2_r3Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst1_MC2_r3Inst_XORInst_0_3_U1  ( .A(MCInst1_MC2_v0_3 [3]), .B(
        MCInst1_MC2_v1_3 [3]), .Z(MCInst1_MC2_r3Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst1_MC3_v0_2Inst_0_U4  ( .A(MCInst1_MC3_v0_2Inst_0_n2 ), .B(
        MCInst1_MC3_v0_0 [3]), .ZN(MCInst1_MC3_v0_2 [0]) );
  XNOR2_X1 MCInst1_MC3_v0_2Inst_0_U3  ( .A(MCInst1_MC3_v0_3 [0]), .B(
        ShiftRowsOutput[48]), .ZN(MCInst1_MC3_v0_2Inst_0_n2 ) );
  XOR2_X1 MCInst1_MC3_v1_1Inst_0_U3  ( .A(MCInst1_MC3_v1_3 [3]), .B(
        MCInst1_MC3_v1_3 [0]), .Z(MCInst1_MC3_v1_1 [0]) );
  XNOR2_X1 MCInst1_MC3_v1_2Inst_0_U4  ( .A(MCInst1_MC3_v1_2Inst_0_n2 ), .B(
        MCInst1_MC3_v1_3 [3]), .ZN(MCInst1_MC3_v1_2 [0]) );
  XNOR2_X1 MCInst1_MC3_v1_2Inst_0_U3  ( .A(MCInst1_MC3_v1_3 [0]), .B(
        MCInst1_MC3_v1_3 [2]), .ZN(MCInst1_MC3_v1_2Inst_0_n2 ) );
  XOR2_X1 MCInst1_MC3_v2_1Inst_0_U3  ( .A(MCInst1_MC3_v2_3 [1]), .B(
        MCInst1_MC3_v2_0 [3]), .Z(MCInst1_MC3_v2_1 [0]) );
  XOR2_X1 MCInst1_MC3_v2_2Inst_0_U3  ( .A(MCInst1_MC3_v2_0 [2]), .B(
        MCInst1_MC3_v2_0 [0]), .Z(MCInst1_MC3_v2_2 [0]) );
  XNOR2_X1 MCInst1_MC3_v2_3Inst_0_U5  ( .A(MCInst1_MC3_v2_3Inst_0_n4 ), .B(
        MCInst1_MC3_v2_3Inst_0_n3 ), .ZN(MCInst1_MC3_v2_3 [0]) );
  XNOR2_X1 MCInst1_MC3_v2_3Inst_0_U4  ( .A(MCInst1_MC3_v2_0 [2]), .B(
        MCInst1_MC3_v2_3 [1]), .ZN(MCInst1_MC3_v2_3Inst_0_n3 ) );
  XOR2_X1 MCInst1_MC3_v2_3Inst_0_U3  ( .A(MCInst1_MC3_v2_0 [3]), .B(
        MCInst1_MC3_v2_0 [0]), .Z(MCInst1_MC3_v2_3Inst_0_n4 ) );
  XOR2_X1 MCInst1_MC3_v3_1Inst_0_U3  ( .A(MCInst1_MC3_v3_0 [3]), .B(
        MCInst1_MC3_v3_2 [2]), .Z(MCInst1_MC3_v3_1 [0]) );
  XOR2_X1 MCInst1_MC3_v3_2Inst_0_U3  ( .A(MCInst1_MC3_v3_2 [3]), .B(
        MCInst1_MC3_v3_0 [2]), .Z(MCInst1_MC3_v3_2 [0]) );
  XNOR2_X1 MCInst1_MC3_v3_3Inst_0_U4  ( .A(MCInst1_MC3_v3_3Inst_0_n2 ), .B(
        MCInst1_MC3_v3_0 [2]), .ZN(MCInst1_MC3_v3_3 [0]) );
  XNOR2_X1 MCInst1_MC3_v3_3Inst_0_U3  ( .A(MCInst1_MC3_v3_2 [2]), .B(
        MCInst1_MC3_v3_2 [3]), .ZN(MCInst1_MC3_v3_3Inst_0_n2 ) );
  XOR2_X1 MCInst1_MC3_v0_0Inst_1_U3  ( .A(MCInst1_MC3_v0_3 [3]), .B(
        MCInst1_MC3_v0_3 [0]), .Z(MCInst1_MC3_v0_0 [1]) );
  XOR2_X1 MCInst1_MC3_v0_1Inst_1_U3  ( .A(MCInst1_MC3_v0_0 [3]), .B(
        MCInst1_MC3_v0_3 [3]), .Z(MCInst1_MC3_v0_1 [1]) );
  XNOR2_X1 MCInst1_MC3_v0_2Inst_1_U4  ( .A(MCInst1_MC3_v0_2Inst_1_n2 ), .B(
        MCInst1_MC3_v0_3 [3]), .ZN(MCInst1_MC3_v0_2 [1]) );
  XNOR2_X1 MCInst1_MC3_v0_2Inst_1_U3  ( .A(MCInst1_MC3_v0_3 [0]), .B(
        ShiftRowsOutput[48]), .ZN(MCInst1_MC3_v0_2Inst_1_n2 ) );
  XOR2_X1 MCInst1_MC3_v0_3Inst_1_U3  ( .A(ShiftRowsOutput[48]), .B(
        MCInst1_MC3_v0_3 [0]), .Z(MCInst1_MC3_v0_3 [1]) );
  XOR2_X1 MCInst1_MC3_v1_1Inst_1_U3  ( .A(ShiftRowsOutput[32]), .B(
        MCInst1_MC3_v1_3 [3]), .Z(MCInst1_MC3_v1_1 [1]) );
  XOR2_X1 MCInst1_MC3_v1_2Inst_1_U3  ( .A(ShiftRowsOutput[32]), .B(
        MCInst1_MC3_v1_3 [2]), .Z(MCInst1_MC3_v1_2 [1]) );
  XOR2_X1 MCInst1_MC3_v1_3Inst_1_U3  ( .A(ShiftRowsOutput[32]), .B(
        MCInst1_MC3_v1_3 [0]), .Z(MCInst1_MC3_v1_3 [1]) );
  XOR2_X1 MCInst1_MC3_v2_0Inst_1_U3  ( .A(MCInst1_MC3_v2_3 [1]), .B(
        MCInst1_MC3_v2_0 [0]), .Z(MCInst1_MC3_v2_0 [1]) );
  XNOR2_X1 MCInst1_MC3_v2_1Inst_1_U4  ( .A(MCInst1_MC3_v2_1Inst_1_n2 ), .B(
        MCInst1_MC3_v2_0 [3]), .ZN(MCInst1_MC3_v2_1 [1]) );
  XNOR2_X1 MCInst1_MC3_v2_1Inst_1_U3  ( .A(MCInst1_MC3_v2_0 [0]), .B(
        MCInst1_MC3_v2_0 [2]), .ZN(MCInst1_MC3_v2_1Inst_1_n2 ) );
  XNOR2_X1 MCInst1_MC3_v2_2Inst_1_U5  ( .A(MCInst1_MC3_v2_2Inst_1_n4 ), .B(
        MCInst1_MC3_v2_2Inst_1_n3 ), .ZN(MCInst1_MC3_v2_2 [1]) );
  XNOR2_X1 MCInst1_MC3_v2_2Inst_1_U4  ( .A(MCInst1_MC3_v2_0 [2]), .B(
        MCInst1_MC3_v2_3 [1]), .ZN(MCInst1_MC3_v2_2Inst_1_n3 ) );
  XOR2_X1 MCInst1_MC3_v2_2Inst_1_U3  ( .A(MCInst1_MC3_v2_0 [3]), .B(
        MCInst1_MC3_v2_0 [0]), .Z(MCInst1_MC3_v2_2Inst_1_n4 ) );
  XOR2_X1 MCInst1_MC3_v3_0Inst_1_U3  ( .A(MCInst1_MC3_v3_2 [3]), .B(
        MCInst1_MC3_v3_2 [2]), .Z(MCInst1_MC3_v3_0 [1]) );
  XOR2_X1 MCInst1_MC3_v3_1Inst_1_U3  ( .A(MCInst1_MC3_v3_2 [3]), .B(
        MCInst1_MC3_v3_0 [3]), .Z(MCInst1_MC3_v3_1 [1]) );
  XNOR2_X1 MCInst1_MC3_v3_3Inst_1_U4  ( .A(MCInst1_MC3_v3_3Inst_1_n2 ), .B(
        MCInst1_MC3_v3_0 [3]), .ZN(MCInst1_MC3_v3_3 [1]) );
  XNOR2_X1 MCInst1_MC3_v3_3Inst_1_U3  ( .A(MCInst1_MC3_v3_2 [2]), .B(
        MCInst1_MC3_v3_2 [3]), .ZN(MCInst1_MC3_v3_3Inst_1_n2 ) );
  XOR2_X1 MCInst1_MC3_v0_0Inst_2_U3  ( .A(ShiftRowsOutput[48]), .B(
        MCInst1_MC3_v0_3 [0]), .Z(MCInst1_MC3_v0_0 [2]) );
  XOR2_X1 MCInst1_MC3_v0_1Inst_2_U3  ( .A(MCInst1_MC3_v0_3 [3]), .B(
        MCInst1_MC3_v0_3 [0]), .Z(MCInst1_MC3_v0_1 [2]) );
  XOR2_X1 MCInst1_MC3_v0_2Inst_2_U3  ( .A(MCInst1_MC3_v0_0 [3]), .B(
        MCInst1_MC3_v0_3 [0]), .Z(MCInst1_MC3_v0_2 [2]) );
  XNOR2_X1 MCInst1_MC3_v1_1Inst_2_U4  ( .A(MCInst1_MC3_v1_1Inst_2_n2 ), .B(
        MCInst1_MC3_v1_3 [2]), .ZN(MCInst1_MC3_v1_1 [2]) );
  XNOR2_X1 MCInst1_MC3_v1_1Inst_2_U3  ( .A(MCInst1_MC3_v1_3 [0]), .B(
        ShiftRowsOutput[32]), .ZN(MCInst1_MC3_v1_1Inst_2_n2 ) );
  XNOR2_X1 MCInst1_MC3_v1_2Inst_2_U4  ( .A(MCInst1_MC3_v1_2Inst_2_n2 ), .B(
        MCInst1_MC3_v1_3 [2]), .ZN(MCInst1_MC3_v1_2 [2]) );
  XNOR2_X1 MCInst1_MC3_v1_2Inst_2_U3  ( .A(MCInst1_MC3_v1_3 [3]), .B(
        ShiftRowsOutput[32]), .ZN(MCInst1_MC3_v1_2Inst_2_n2 ) );
  XNOR2_X1 MCInst1_MC3_v2_1Inst_2_U4  ( .A(MCInst1_MC3_v2_1Inst_2_n2 ), .B(
        MCInst1_MC3_v2_0 [3]), .ZN(MCInst1_MC3_v2_1 [2]) );
  XNOR2_X1 MCInst1_MC3_v2_1Inst_2_U3  ( .A(MCInst1_MC3_v2_0 [0]), .B(
        MCInst1_MC3_v2_3 [1]), .ZN(MCInst1_MC3_v2_1Inst_2_n2 ) );
  XNOR2_X1 MCInst1_MC3_v2_2Inst_2_U4  ( .A(MCInst1_MC3_v2_2Inst_2_n2 ), .B(
        MCInst1_MC3_v2_0 [3]), .ZN(MCInst1_MC3_v2_2 [2]) );
  XNOR2_X1 MCInst1_MC3_v2_2Inst_2_U3  ( .A(MCInst1_MC3_v2_0 [0]), .B(
        MCInst1_MC3_v2_0 [2]), .ZN(MCInst1_MC3_v2_2Inst_2_n2 ) );
  XOR2_X1 MCInst1_MC3_v2_3Inst_2_U3  ( .A(MCInst1_MC3_v2_3 [1]), .B(
        MCInst1_MC3_v2_0 [2]), .Z(MCInst1_MC3_v2_3 [2]) );
  XNOR2_X1 MCInst1_MC3_v3_1Inst_2_U4  ( .A(MCInst1_MC3_v3_1Inst_2_n2 ), .B(
        MCInst1_MC3_v3_0 [2]), .ZN(MCInst1_MC3_v3_1 [2]) );
  XNOR2_X1 MCInst1_MC3_v3_1Inst_2_U3  ( .A(MCInst1_MC3_v3_2 [2]), .B(
        MCInst1_MC3_v3_2 [3]), .ZN(MCInst1_MC3_v3_1Inst_2_n2 ) );
  XOR2_X1 MCInst1_MC3_v3_3Inst_2_U3  ( .A(MCInst1_MC3_v3_0 [2]), .B(
        MCInst1_MC3_v3_2 [2]), .Z(MCInst1_MC3_v3_3 [2]) );
  XOR2_X1 MCInst1_MC3_v0_1Inst_3_U3  ( .A(ShiftRowsOutput[48]), .B(
        MCInst1_MC3_v0_3 [0]), .Z(MCInst1_MC3_v0_1 [3]) );
  XOR2_X1 MCInst1_MC3_v0_2Inst_3_U3  ( .A(ShiftRowsOutput[48]), .B(
        MCInst1_MC3_v0_3 [3]), .Z(MCInst1_MC3_v0_2 [3]) );
  XOR2_X1 MCInst1_MC3_v1_1Inst_3_U3  ( .A(MCInst1_MC3_v1_3 [2]), .B(
        MCInst1_MC3_v1_3 [3]), .Z(MCInst1_MC3_v1_1 [3]) );
  XNOR2_X1 MCInst1_MC3_v1_2Inst_3_U5  ( .A(MCInst1_MC3_v1_2Inst_3_n4 ), .B(
        MCInst1_MC3_v1_2Inst_3_n3 ), .ZN(MCInst1_MC3_v1_2 [3]) );
  XNOR2_X1 MCInst1_MC3_v1_2Inst_3_U4  ( .A(MCInst1_MC3_v1_3 [2]), .B(
        ShiftRowsOutput[32]), .ZN(MCInst1_MC3_v1_2Inst_3_n3 ) );
  XOR2_X1 MCInst1_MC3_v1_2Inst_3_U3  ( .A(MCInst1_MC3_v1_3 [3]), .B(
        MCInst1_MC3_v1_3 [0]), .Z(MCInst1_MC3_v1_2Inst_3_n4 ) );
  XOR2_X1 MCInst1_MC3_v2_1Inst_3_U3  ( .A(MCInst1_MC3_v2_0 [2]), .B(
        MCInst1_MC3_v2_0 [0]), .Z(MCInst1_MC3_v2_1 [3]) );
  XNOR2_X1 MCInst1_MC3_v2_2Inst_3_U4  ( .A(MCInst1_MC3_v2_2Inst_3_n2 ), .B(
        MCInst1_MC3_v2_0 [3]), .ZN(MCInst1_MC3_v2_2 [3]) );
  XNOR2_X1 MCInst1_MC3_v2_2Inst_3_U3  ( .A(MCInst1_MC3_v2_0 [0]), .B(
        MCInst1_MC3_v2_3 [1]), .ZN(MCInst1_MC3_v2_2Inst_3_n2 ) );
  XNOR2_X1 MCInst1_MC3_v2_3Inst_3_U4  ( .A(MCInst1_MC3_v2_3Inst_3_n2 ), .B(
        MCInst1_MC3_v2_0 [2]), .ZN(MCInst1_MC3_v2_3 [3]) );
  XNOR2_X1 MCInst1_MC3_v2_3Inst_3_U3  ( .A(MCInst1_MC3_v2_0 [3]), .B(
        MCInst1_MC3_v2_3 [1]), .ZN(MCInst1_MC3_v2_3Inst_3_n2 ) );
  XOR2_X1 MCInst1_MC3_v3_1Inst_3_U3  ( .A(MCInst1_MC3_v3_0 [2]), .B(
        MCInst1_MC3_v3_0 [3]), .Z(MCInst1_MC3_v3_1 [3]) );
  XOR2_X1 MCInst1_MC3_v3_3Inst_3_U3  ( .A(MCInst1_MC3_v3_2 [3]), .B(
        MCInst1_MC3_v3_0 [3]), .Z(MCInst1_MC3_v3_3 [3]) );
  XNOR2_X1 MCInst1_MC3_r0Inst_XORInst_0_0_U3  ( .A(
        MCInst1_MC3_r0Inst_XORInst_0_0_n5 ), .B(
        MCInst1_MC3_r0Inst_XORInst_0_0_n4 ), .ZN(Feedback[48]) );
  XNOR2_X1 MCInst1_MC3_r0Inst_XORInst_0_0_U2  ( .A(MCInst1_MC3_v3_2 [2]), 
        .B(MCInst1_MC3_v2_0 [0]), .ZN(MCInst1_MC3_r0Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst1_MC3_r0Inst_XORInst_0_0_U1  ( .A(MCInst1_MC3_v0_3 [3]), .B(
        ShiftRowsOutput[32]), .Z(MCInst1_MC3_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst1_MC3_r0Inst_XORInst_0_1_U3  ( .A(
        MCInst1_MC3_r0Inst_XORInst_0_1_n5 ), .B(
        MCInst1_MC3_r0Inst_XORInst_0_1_n4 ), .ZN(Feedback[49]) );
  XNOR2_X1 MCInst1_MC3_r0Inst_XORInst_0_1_U2  ( .A(MCInst1_MC3_v3_0 [1]), 
        .B(MCInst1_MC3_v2_0 [1]), .ZN(MCInst1_MC3_r0Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst1_MC3_r0Inst_XORInst_0_1_U1  ( .A(MCInst1_MC3_v0_0 [1]), .B(
        MCInst1_MC3_v1_3 [2]), .Z(MCInst1_MC3_r0Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst1_MC3_r0Inst_XORInst_0_2_U3  ( .A(
        MCInst1_MC3_r0Inst_XORInst_0_2_n5 ), .B(
        MCInst1_MC3_r0Inst_XORInst_0_2_n4 ), .ZN(Feedback[50]) );
  XNOR2_X1 MCInst1_MC3_r0Inst_XORInst_0_2_U2  ( .A(MCInst1_MC3_v3_0 [2]), 
        .B(MCInst1_MC3_v2_0 [2]), .ZN(MCInst1_MC3_r0Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst1_MC3_r0Inst_XORInst_0_2_U1  ( .A(MCInst1_MC3_v0_0 [2]), .B(
        MCInst1_MC3_v1_3 [3]), .Z(MCInst1_MC3_r0Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst1_MC3_r0Inst_XORInst_0_3_U3  ( .A(
        MCInst1_MC3_r0Inst_XORInst_0_3_n5 ), .B(
        MCInst1_MC3_r0Inst_XORInst_0_3_n4 ), .ZN(Feedback[51]) );
  XNOR2_X1 MCInst1_MC3_r0Inst_XORInst_0_3_U2  ( .A(MCInst1_MC3_v3_0 [3]), 
        .B(MCInst1_MC3_v2_0 [3]), .ZN(MCInst1_MC3_r0Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst1_MC3_r0Inst_XORInst_0_3_U1  ( .A(MCInst1_MC3_v0_0 [3]), .B(
        MCInst1_MC3_v1_3 [0]), .Z(MCInst1_MC3_r0Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst1_MC3_r1Inst_XORInst_0_0_U3  ( .A(
        MCInst1_MC3_r1Inst_XORInst_0_0_n5 ), .B(
        MCInst1_MC3_r1Inst_XORInst_0_0_n4 ), .ZN(Feedback[32]) );
  XNOR2_X1 MCInst1_MC3_r1Inst_XORInst_0_0_U2  ( .A(MCInst1_MC3_v3_1 [0]), 
        .B(MCInst1_MC3_v2_1 [0]), .ZN(MCInst1_MC3_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst1_MC3_r1Inst_XORInst_0_0_U1  ( .A(MCInst1_MC3_v0_0 [3]), .B(
        MCInst1_MC3_v1_1 [0]), .Z(MCInst1_MC3_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst1_MC3_r1Inst_XORInst_0_1_U3  ( .A(
        MCInst1_MC3_r1Inst_XORInst_0_1_n5 ), .B(
        MCInst1_MC3_r1Inst_XORInst_0_1_n4 ), .ZN(Feedback[33]) );
  XNOR2_X1 MCInst1_MC3_r1Inst_XORInst_0_1_U2  ( .A(MCInst1_MC3_v3_1 [1]), 
        .B(MCInst1_MC3_v2_1 [1]), .ZN(MCInst1_MC3_r1Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst1_MC3_r1Inst_XORInst_0_1_U1  ( .A(MCInst1_MC3_v0_1 [1]), .B(
        MCInst1_MC3_v1_1 [1]), .Z(MCInst1_MC3_r1Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst1_MC3_r1Inst_XORInst_0_2_U3  ( .A(
        MCInst1_MC3_r1Inst_XORInst_0_2_n5 ), .B(
        MCInst1_MC3_r1Inst_XORInst_0_2_n4 ), .ZN(Feedback[34]) );
  XNOR2_X1 MCInst1_MC3_r1Inst_XORInst_0_2_U2  ( .A(MCInst1_MC3_v3_1 [2]), 
        .B(MCInst1_MC3_v2_1 [2]), .ZN(MCInst1_MC3_r1Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst1_MC3_r1Inst_XORInst_0_2_U1  ( .A(MCInst1_MC3_v0_1 [2]), .B(
        MCInst1_MC3_v1_1 [2]), .Z(MCInst1_MC3_r1Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst1_MC3_r1Inst_XORInst_0_3_U3  ( .A(
        MCInst1_MC3_r1Inst_XORInst_0_3_n5 ), .B(
        MCInst1_MC3_r1Inst_XORInst_0_3_n4 ), .ZN(Feedback[35]) );
  XNOR2_X1 MCInst1_MC3_r1Inst_XORInst_0_3_U2  ( .A(MCInst1_MC3_v3_1 [3]), 
        .B(MCInst1_MC3_v2_1 [3]), .ZN(MCInst1_MC3_r1Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst1_MC3_r1Inst_XORInst_0_3_U1  ( .A(MCInst1_MC3_v0_1 [3]), .B(
        MCInst1_MC3_v1_1 [3]), .Z(MCInst1_MC3_r1Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst1_MC3_r2Inst_XORInst_0_0_U3  ( .A(
        MCInst1_MC3_r2Inst_XORInst_0_0_n5 ), .B(
        MCInst1_MC3_r2Inst_XORInst_0_0_n4 ), .ZN(Feedback[16]) );
  XNOR2_X1 MCInst1_MC3_r2Inst_XORInst_0_0_U2  ( .A(MCInst1_MC3_v3_2 [0]), 
        .B(MCInst1_MC3_v2_2 [0]), .ZN(MCInst1_MC3_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst1_MC3_r2Inst_XORInst_0_0_U1  ( .A(MCInst1_MC3_v0_2 [0]), .B(
        MCInst1_MC3_v1_2 [0]), .Z(MCInst1_MC3_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst1_MC3_r2Inst_XORInst_0_1_U3  ( .A(
        MCInst1_MC3_r2Inst_XORInst_0_1_n5 ), .B(
        MCInst1_MC3_r2Inst_XORInst_0_1_n4 ), .ZN(Feedback[17]) );
  XNOR2_X1 MCInst1_MC3_r2Inst_XORInst_0_1_U2  ( .A(MCInst1_MC3_v3_0 [3]), 
        .B(MCInst1_MC3_v2_2 [1]), .ZN(MCInst1_MC3_r2Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst1_MC3_r2Inst_XORInst_0_1_U1  ( .A(MCInst1_MC3_v0_2 [1]), .B(
        MCInst1_MC3_v1_2 [1]), .Z(MCInst1_MC3_r2Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst1_MC3_r2Inst_XORInst_0_2_U3  ( .A(
        MCInst1_MC3_r2Inst_XORInst_0_2_n5 ), .B(
        MCInst1_MC3_r2Inst_XORInst_0_2_n4 ), .ZN(Feedback[18]) );
  XNOR2_X1 MCInst1_MC3_r2Inst_XORInst_0_2_U2  ( .A(MCInst1_MC3_v3_2 [2]), 
        .B(MCInst1_MC3_v2_2 [2]), .ZN(MCInst1_MC3_r2Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst1_MC3_r2Inst_XORInst_0_2_U1  ( .A(MCInst1_MC3_v0_2 [2]), .B(
        MCInst1_MC3_v1_2 [2]), .Z(MCInst1_MC3_r2Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst1_MC3_r2Inst_XORInst_0_3_U3  ( .A(
        MCInst1_MC3_r2Inst_XORInst_0_3_n5 ), .B(
        MCInst1_MC3_r2Inst_XORInst_0_3_n4 ), .ZN(Feedback[19]) );
  XNOR2_X1 MCInst1_MC3_r2Inst_XORInst_0_3_U2  ( .A(MCInst1_MC3_v3_2 [3]), 
        .B(MCInst1_MC3_v2_2 [3]), .ZN(MCInst1_MC3_r2Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst1_MC3_r2Inst_XORInst_0_3_U1  ( .A(MCInst1_MC3_v0_2 [3]), .B(
        MCInst1_MC3_v1_2 [3]), .Z(MCInst1_MC3_r2Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst1_MC3_r3Inst_XORInst_0_0_U3  ( .A(
        MCInst1_MC3_r3Inst_XORInst_0_0_n5 ), .B(
        MCInst1_MC3_r3Inst_XORInst_0_0_n4 ), .ZN(Feedback[0]) );
  XNOR2_X1 MCInst1_MC3_r3Inst_XORInst_0_0_U2  ( .A(MCInst1_MC3_v3_3 [0]), 
        .B(MCInst1_MC3_v2_3 [0]), .ZN(MCInst1_MC3_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst1_MC3_r3Inst_XORInst_0_0_U1  ( .A(MCInst1_MC3_v0_3 [0]), .B(
        MCInst1_MC3_v1_3 [0]), .Z(MCInst1_MC3_r3Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst1_MC3_r3Inst_XORInst_0_1_U3  ( .A(
        MCInst1_MC3_r3Inst_XORInst_0_1_n5 ), .B(
        MCInst1_MC3_r3Inst_XORInst_0_1_n4 ), .ZN(Feedback[1]) );
  XNOR2_X1 MCInst1_MC3_r3Inst_XORInst_0_1_U2  ( .A(MCInst1_MC3_v3_3 [1]), 
        .B(MCInst1_MC3_v2_3 [1]), .ZN(MCInst1_MC3_r3Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst1_MC3_r3Inst_XORInst_0_1_U1  ( .A(MCInst1_MC3_v0_3 [1]), .B(
        MCInst1_MC3_v1_3 [1]), .Z(MCInst1_MC3_r3Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst1_MC3_r3Inst_XORInst_0_2_U3  ( .A(
        MCInst1_MC3_r3Inst_XORInst_0_2_n5 ), .B(
        MCInst1_MC3_r3Inst_XORInst_0_2_n4 ), .ZN(Feedback[2]) );
  XNOR2_X1 MCInst1_MC3_r3Inst_XORInst_0_2_U2  ( .A(MCInst1_MC3_v3_3 [2]), 
        .B(MCInst1_MC3_v2_3 [2]), .ZN(MCInst1_MC3_r3Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst1_MC3_r3Inst_XORInst_0_2_U1  ( .A(MCInst1_MC3_v0_0 [3]), .B(
        MCInst1_MC3_v1_3 [2]), .Z(MCInst1_MC3_r3Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst1_MC3_r3Inst_XORInst_0_3_U3  ( .A(
        MCInst1_MC3_r3Inst_XORInst_0_3_n5 ), .B(
        MCInst1_MC3_r3Inst_XORInst_0_3_n4 ), .ZN(Feedback[3]) );
  XNOR2_X1 MCInst1_MC3_r3Inst_XORInst_0_3_U2  ( .A(MCInst1_MC3_v3_3 [3]), 
        .B(MCInst1_MC3_v2_3 [3]), .ZN(MCInst1_MC3_r3Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst1_MC3_r3Inst_XORInst_0_3_U1  ( .A(MCInst1_MC3_v0_3 [3]), .B(
        MCInst1_MC3_v1_3 [3]), .Z(MCInst1_MC3_r3Inst_XORInst_0_3_n5 ) );
  DFF_X1 StateReg_s_current_state_reg[0]  ( .D(Feedback[0]), .CK(clk), .Q(
        SubCellInput[0]) );
  DFF_X1 StateReg_s_current_state_reg[1]  ( .D(Feedback[1]), .CK(clk), .Q(
        SubCellInput[1]) );
  DFF_X1 StateReg_s_current_state_reg[2]  ( .D(Feedback[2]), .CK(clk), .Q(
        SubCellInput[2]) );
  DFF_X1 StateReg_s_current_state_reg[3]  ( .D(Feedback[3]), .CK(clk), .Q(
        SubCellInput[3]) );
  DFF_X1 StateReg_s_current_state_reg[4]  ( .D(Feedback[4]), .CK(clk), .Q(
        SubCellInput[4]) );
  DFF_X1 StateReg_s_current_state_reg[5]  ( .D(Feedback[5]), .CK(clk), .Q(
        SubCellInput[5]) );
  DFF_X1 StateReg_s_current_state_reg[6]  ( .D(Feedback[6]), .CK(clk), .Q(
        SubCellInput[6]) );
  DFF_X1 StateReg_s_current_state_reg[7]  ( .D(Feedback[7]), .CK(clk), .Q(
        SubCellInput[7]) );
  DFF_X1 StateReg_s_current_state_reg[8]  ( .D(Feedback[8]), .CK(clk), .Q(
        SubCellInput[8]) );
  DFF_X1 StateReg_s_current_state_reg[9]  ( .D(Feedback[9]), .CK(clk), .Q(
        SubCellInput[9]) );
  DFF_X1 StateReg_s_current_state_reg[10]  ( .D(Feedback[10]), .CK(clk), .Q(
        SubCellInput[10]) );
  DFF_X1 StateReg_s_current_state_reg[11]  ( .D(Feedback[11]), .CK(clk), .Q(
        SubCellInput[11]) );
  DFF_X1 StateReg_s_current_state_reg[12]  ( .D(Feedback[12]), .CK(clk), .Q(
        SubCellInput[12]) );
  DFF_X1 StateReg_s_current_state_reg[13]  ( .D(Feedback[13]), .CK(clk), .Q(
        SubCellInput[13]) );
  DFF_X1 StateReg_s_current_state_reg[14]  ( .D(Feedback[14]), .CK(clk), .Q(
        SubCellInput[14]) );
  DFF_X1 StateReg_s_current_state_reg[15]  ( .D(Feedback[15]), .CK(clk), .Q(
        SubCellInput[15]) );
  DFF_X1 StateReg_s_current_state_reg[16]  ( .D(Feedback[16]), .CK(clk), .Q(
        SubCellInput[16]) );
  DFF_X1 StateReg_s_current_state_reg[17]  ( .D(Feedback[17]), .CK(clk), .Q(
        SubCellInput[17]) );
  DFF_X1 StateReg_s_current_state_reg[18]  ( .D(Feedback[18]), .CK(clk), .Q(
        SubCellInput[18]) );
  DFF_X1 StateReg_s_current_state_reg[19]  ( .D(Feedback[19]), .CK(clk), .Q(
        SubCellInput[19]) );
  DFF_X1 StateReg_s_current_state_reg[20]  ( .D(Feedback[20]), .CK(clk), .Q(
        SubCellInput[20]) );
  DFF_X1 StateReg_s_current_state_reg[21]  ( .D(Feedback[21]), .CK(clk), .Q(
        SubCellInput[21]) );
  DFF_X1 StateReg_s_current_state_reg[22]  ( .D(Feedback[22]), .CK(clk), .Q(
        SubCellInput[22]) );
  DFF_X1 StateReg_s_current_state_reg[23]  ( .D(Feedback[23]), .CK(clk), .Q(
        SubCellInput[23]) );
  DFF_X1 StateReg_s_current_state_reg[24]  ( .D(Feedback[24]), .CK(clk), .Q(
        SubCellInput[24]) );
  DFF_X1 StateReg_s_current_state_reg[25]  ( .D(Feedback[25]), .CK(clk), .Q(
        SubCellInput[25]) );
  DFF_X1 StateReg_s_current_state_reg[26]  ( .D(Feedback[26]), .CK(clk), .Q(
        SubCellInput[26]) );
  DFF_X1 StateReg_s_current_state_reg[27]  ( .D(Feedback[27]), .CK(clk), .Q(
        SubCellInput[27]) );
  DFF_X1 StateReg_s_current_state_reg[28]  ( .D(Feedback[28]), .CK(clk), .Q(
        SubCellInput[28]) );
  DFF_X1 StateReg_s_current_state_reg[29]  ( .D(Feedback[29]), .CK(clk), .Q(
        SubCellInput[29]) );
  DFF_X1 StateReg_s_current_state_reg[30]  ( .D(Feedback[30]), .CK(clk), .Q(
        SubCellInput[30]) );
  DFF_X1 StateReg_s_current_state_reg[31]  ( .D(Feedback[31]), .CK(clk), .Q(
        SubCellInput[31]) );
  DFF_X1 StateReg_s_current_state_reg[32]  ( .D(Feedback[32]), .CK(clk), .Q(
        SubCellInput[32]) );
  DFF_X1 StateReg_s_current_state_reg[33]  ( .D(Feedback[33]), .CK(clk), .Q(
        SubCellInput[33]) );
  DFF_X1 StateReg_s_current_state_reg[34]  ( .D(Feedback[34]), .CK(clk), .Q(
        SubCellInput[34]) );
  DFF_X1 StateReg_s_current_state_reg[35]  ( .D(Feedback[35]), .CK(clk), .Q(
        SubCellInput[35]) );
  DFF_X1 StateReg_s_current_state_reg[36]  ( .D(Feedback[36]), .CK(clk), .Q(
        SubCellInput[36]) );
  DFF_X1 StateReg_s_current_state_reg[37]  ( .D(Feedback[37]), .CK(clk), .Q(
        SubCellInput[37]) );
  DFF_X1 StateReg_s_current_state_reg[38]  ( .D(Feedback[38]), .CK(clk), .Q(
        SubCellInput[38]) );
  DFF_X1 StateReg_s_current_state_reg[39]  ( .D(Feedback[39]), .CK(clk), .Q(
        SubCellInput[39]) );
  DFF_X1 StateReg_s_current_state_reg[40]  ( .D(Feedback[40]), .CK(clk), .Q(
        SubCellInput[40]) );
  DFF_X1 StateReg_s_current_state_reg[41]  ( .D(Feedback[41]), .CK(clk), .Q(
        SubCellInput[41]) );
  DFF_X1 StateReg_s_current_state_reg[42]  ( .D(Feedback[42]), .CK(clk), .Q(
        SubCellInput[42]) );
  DFF_X1 StateReg_s_current_state_reg[43]  ( .D(Feedback[43]), .CK(clk), .Q(
        SubCellInput[43]) );
  DFF_X1 StateReg_s_current_state_reg[44]  ( .D(Feedback[44]), .CK(clk), .Q(
        SubCellInput[44]) );
  DFF_X1 StateReg_s_current_state_reg[45]  ( .D(Feedback[45]), .CK(clk), .Q(
        SubCellInput[45]) );
  DFF_X1 StateReg_s_current_state_reg[46]  ( .D(Feedback[46]), .CK(clk), .Q(
        SubCellInput[46]) );
  DFF_X1 StateReg_s_current_state_reg[47]  ( .D(Feedback[47]), .CK(clk), .Q(
        SubCellInput[47]) );
  DFF_X1 StateReg_s_current_state_reg[48]  ( .D(Feedback[48]), .CK(clk), .Q(
        SubCellInput[48]) );
  DFF_X1 StateReg_s_current_state_reg[49]  ( .D(Feedback[49]), .CK(clk), .Q(
        SubCellInput[49]) );
  DFF_X1 StateReg_s_current_state_reg[50]  ( .D(Feedback[50]), .CK(clk), .Q(
        SubCellInput[50]) );
  DFF_X1 StateReg_s_current_state_reg[51]  ( .D(Feedback[51]), .CK(clk), .Q(
        SubCellInput[51]) );
  DFF_X1 StateReg_s_current_state_reg[52]  ( .D(Feedback[52]), .CK(clk), .Q(
        SubCellInput[52]) );
  DFF_X1 StateReg_s_current_state_reg[53]  ( .D(Feedback[53]), .CK(clk), .Q(
        SubCellInput[53]) );
  DFF_X1 StateReg_s_current_state_reg[54]  ( .D(Feedback[54]), .CK(clk), .Q(
        SubCellInput[54]) );
  DFF_X1 StateReg_s_current_state_reg[55]  ( .D(Feedback[55]), .CK(clk), .Q(
        SubCellInput[55]) );
  DFF_X1 StateReg_s_current_state_reg[56]  ( .D(Feedback[56]), .CK(clk), .Q(
        SubCellInput[56]) );
  DFF_X1 StateReg_s_current_state_reg[57]  ( .D(Feedback[57]), .CK(clk), .Q(
        SubCellInput[57]) );
  DFF_X1 StateReg_s_current_state_reg[58]  ( .D(Feedback[58]), .CK(clk), .Q(
        SubCellInput[58]) );
  DFF_X1 StateReg_s_current_state_reg[59]  ( .D(Feedback[59]), .CK(clk), .Q(
        SubCellInput[59]) );
  DFF_X1 StateReg_s_current_state_reg[60]  ( .D(Feedback[60]), .CK(clk), .Q(
        SubCellInput[60]) );
  DFF_X1 StateReg_s_current_state_reg[61]  ( .D(Feedback[61]), .CK(clk), .Q(
        SubCellInput[61]) );
  DFF_X1 StateReg_s_current_state_reg[62]  ( .D(Feedback[62]), .CK(clk), .Q(
        SubCellInput[62]) );
  DFF_X1 StateReg_s_current_state_reg[63]  ( .D(Feedback[63]), .CK(clk), .Q(
        SubCellInput[63]) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_3_U9  ( .A1(
        SubCellInst2_LFInst_0_LFInst_3_n16 ), .A2(
        SubCellInst2_LFInst_0_LFInst_3_n15 ), .ZN(MCInst2_MC0_v3_2 [2]) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_3_U8  ( .A1(SubCellInput[1]), .A2(
        SubCellInst2_LFInst_0_LFInst_3_n14 ), .ZN(
        SubCellInst2_LFInst_0_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst2_LFInst_0_LFInst_3_U7  ( .A(SubCellInput[3]), .B(
        SubCellInput[2]), .Z(SubCellInst2_LFInst_0_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_3_U6  ( .A1(
        SubCellInst2_LFInst_0_LFInst_3_n13 ), .A2(
        SubCellInst2_LFInst_0_LFInst_3_n12 ), .ZN(
        SubCellInst2_LFInst_0_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_3_U5  ( .A1(SubCellInput[0]), .A2(
        SubCellInput[2]), .ZN(SubCellInst2_LFInst_0_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst2_LFInst_0_LFInst_3_U4  ( .A(SubCellInput[0]), .B(
        SubCellInst2_LFInst_0_LFInst_3_n11 ), .ZN(
        SubCellInst2_LFInst_0_LFInst_3_n13 ) );
  OR2_X1 SubCellInst2_LFInst_0_LFInst_3_U3  ( .A1(SubCellInput[3]), .A2(
        SubCellInput[1]), .ZN(SubCellInst2_LFInst_0_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_2_U11  ( .A1(
        SubCellInst2_LFInst_0_LFInst_2_n22 ), .A2(
        SubCellInst2_LFInst_0_LFInst_2_n21 ), .ZN(MCInst2_MC0_v3_0 [3]) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_2_U10  ( .A1(SubCellInput[2]), .A2(
        SubCellInst2_LFInst_0_LFInst_2_n20 ), .ZN(
        SubCellInst2_LFInst_0_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst2_LFInst_0_LFInst_2_U9  ( .A1(SubCellInput[1]), .A2(
        SubCellInst2_LFInst_0_LFInst_2_n19 ), .ZN(
        SubCellInst2_LFInst_0_LFInst_2_n20 ) );
  INV_X1 SubCellInst2_LFInst_0_LFInst_2_U8  ( .A(SubCellInput[3]), .ZN(
        SubCellInst2_LFInst_0_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_2_U7  ( .A1(
        SubCellInst2_LFInst_0_LFInst_2_n18 ), .A2(
        SubCellInst2_LFInst_0_LFInst_2_n17 ), .ZN(
        SubCellInst2_LFInst_0_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst2_LFInst_0_LFInst_2_U6  ( .A(
        SubCellInst2_LFInst_0_LFInst_2_n16 ), .B(SubCellInput[2]), .Z(
        SubCellInst2_LFInst_0_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_2_U5  ( .A1(SubCellInput[0]), .A2(
        SubCellInput[1]), .ZN(SubCellInst2_LFInst_0_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_2_U4  ( .A1(
        SubCellInst2_LFInst_0_LFInst_2_n15 ), .A2(SubCellInput[3]), .ZN(
        SubCellInst2_LFInst_0_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst2_LFInst_0_LFInst_2_U3  ( .A(SubCellInput[0]), .B(
        SubCellInput[1]), .ZN(SubCellInst2_LFInst_0_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_1_U12  ( .A1(
        SubCellInst2_LFInst_0_LFInst_1_n18 ), .A2(
        SubCellInst2_LFInst_0_LFInst_1_n17 ), .ZN(MCInst2_MC0_v3_0 [2]) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_1_U11  ( .A1(SubCellInput[1]), .A2(
        SubCellInst2_LFInst_0_LFInst_1_n16 ), .ZN(
        SubCellInst2_LFInst_0_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst2_LFInst_0_LFInst_1_U10  ( .A1(SubCellInput[3]), .A2(
        SubCellInst2_LFInst_0_LFInst_1_n15 ), .ZN(
        SubCellInst2_LFInst_0_LFInst_1_n16 ) );
  AND2_X1 SubCellInst2_LFInst_0_LFInst_1_U9  ( .A1(SubCellInput[0]), .A2(
        SubCellInput[2]), .ZN(SubCellInst2_LFInst_0_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_1_U8  ( .A1(SubCellInput[3]), .A2(
        SubCellInst2_LFInst_0_LFInst_1_n14 ), .ZN(
        SubCellInst2_LFInst_0_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_1_U7  ( .A1(
        SubCellInst2_LFInst_0_LFInst_1_n13 ), .A2(
        SubCellInst2_LFInst_0_LFInst_1_n12 ), .ZN(
        SubCellInst2_LFInst_0_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_1_U6  ( .A1(SubCellInput[0]), .A2(
        SubCellInput[2]), .ZN(SubCellInst2_LFInst_0_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_1_U5  ( .A1(
        SubCellInst2_LFInst_0_LFInst_1_n11 ), .A2(
        SubCellInst2_LFInst_0_LFInst_1_n10 ), .ZN(
        SubCellInst2_LFInst_0_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_1_U4  ( .A1(SubCellInput[0]), .A2(
        SubCellInput[1]), .ZN(SubCellInst2_LFInst_0_LFInst_1_n10 ) );
  INV_X1 SubCellInst2_LFInst_0_LFInst_1_U3  ( .A(SubCellInput[2]), .ZN(
        SubCellInst2_LFInst_0_LFInst_1_n11 ) );
  XNOR2_X1 SubCellInst2_LFInst_0_LFInst_0_U6  ( .A(
        SubCellInst2_LFInst_0_LFInst_0_n6 ), .B(
        SubCellInst2_LFInst_0_LFInst_0_n5 ), .ZN(MCInst2_MC0_v3_2 [3]) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_0_U5  ( .A1(SubCellInput[2]), .A2(
        SubCellInst2_LFInst_0_LFInst_0_n4 ), .ZN(
        SubCellInst2_LFInst_0_LFInst_0_n5 ) );
  INV_X1 SubCellInst2_LFInst_0_LFInst_0_U4  ( .A(SubCellInput[1]), .ZN(
        SubCellInst2_LFInst_0_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst2_LFInst_0_LFInst_0_U3  ( .A(SubCellInput[0]), .B(
        SubCellInput[3]), .Z(SubCellInst2_LFInst_0_LFInst_0_n6 ) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_3_U9  ( .A1(
        SubCellInst2_LFInst_1_LFInst_3_n16 ), .A2(
        SubCellInst2_LFInst_1_LFInst_3_n15 ), .ZN(MCInst2_MC3_v3_2 [2]) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_3_U8  ( .A1(SubCellInput[5]), .A2(
        SubCellInst2_LFInst_1_LFInst_3_n14 ), .ZN(
        SubCellInst2_LFInst_1_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst2_LFInst_1_LFInst_3_U7  ( .A(SubCellInput[7]), .B(
        SubCellInput[6]), .Z(SubCellInst2_LFInst_1_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_3_U6  ( .A1(
        SubCellInst2_LFInst_1_LFInst_3_n13 ), .A2(
        SubCellInst2_LFInst_1_LFInst_3_n12 ), .ZN(
        SubCellInst2_LFInst_1_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_3_U5  ( .A1(SubCellInput[4]), .A2(
        SubCellInput[6]), .ZN(SubCellInst2_LFInst_1_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst2_LFInst_1_LFInst_3_U4  ( .A(SubCellInput[4]), .B(
        SubCellInst2_LFInst_1_LFInst_3_n11 ), .ZN(
        SubCellInst2_LFInst_1_LFInst_3_n13 ) );
  OR2_X1 SubCellInst2_LFInst_1_LFInst_3_U3  ( .A1(SubCellInput[7]), .A2(
        SubCellInput[5]), .ZN(SubCellInst2_LFInst_1_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_2_U11  ( .A1(
        SubCellInst2_LFInst_1_LFInst_2_n22 ), .A2(
        SubCellInst2_LFInst_1_LFInst_2_n21 ), .ZN(MCInst2_MC3_v3_0 [3]) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_2_U10  ( .A1(SubCellInput[6]), .A2(
        SubCellInst2_LFInst_1_LFInst_2_n20 ), .ZN(
        SubCellInst2_LFInst_1_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst2_LFInst_1_LFInst_2_U9  ( .A1(SubCellInput[5]), .A2(
        SubCellInst2_LFInst_1_LFInst_2_n19 ), .ZN(
        SubCellInst2_LFInst_1_LFInst_2_n20 ) );
  INV_X1 SubCellInst2_LFInst_1_LFInst_2_U8  ( .A(SubCellInput[7]), .ZN(
        SubCellInst2_LFInst_1_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_2_U7  ( .A1(
        SubCellInst2_LFInst_1_LFInst_2_n18 ), .A2(
        SubCellInst2_LFInst_1_LFInst_2_n17 ), .ZN(
        SubCellInst2_LFInst_1_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst2_LFInst_1_LFInst_2_U6  ( .A(
        SubCellInst2_LFInst_1_LFInst_2_n16 ), .B(SubCellInput[6]), .Z(
        SubCellInst2_LFInst_1_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_2_U5  ( .A1(SubCellInput[4]), .A2(
        SubCellInput[5]), .ZN(SubCellInst2_LFInst_1_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_2_U4  ( .A1(
        SubCellInst2_LFInst_1_LFInst_2_n15 ), .A2(SubCellInput[7]), .ZN(
        SubCellInst2_LFInst_1_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst2_LFInst_1_LFInst_2_U3  ( .A(SubCellInput[4]), .B(
        SubCellInput[5]), .ZN(SubCellInst2_LFInst_1_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_1_U12  ( .A1(
        SubCellInst2_LFInst_1_LFInst_1_n18 ), .A2(
        SubCellInst2_LFInst_1_LFInst_1_n17 ), .ZN(MCInst2_MC3_v3_0 [2]) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_1_U11  ( .A1(SubCellInput[5]), .A2(
        SubCellInst2_LFInst_1_LFInst_1_n16 ), .ZN(
        SubCellInst2_LFInst_1_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst2_LFInst_1_LFInst_1_U10  ( .A1(SubCellInput[7]), .A2(
        SubCellInst2_LFInst_1_LFInst_1_n15 ), .ZN(
        SubCellInst2_LFInst_1_LFInst_1_n16 ) );
  AND2_X1 SubCellInst2_LFInst_1_LFInst_1_U9  ( .A1(SubCellInput[4]), .A2(
        SubCellInput[6]), .ZN(SubCellInst2_LFInst_1_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_1_U8  ( .A1(SubCellInput[7]), .A2(
        SubCellInst2_LFInst_1_LFInst_1_n14 ), .ZN(
        SubCellInst2_LFInst_1_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_1_U7  ( .A1(
        SubCellInst2_LFInst_1_LFInst_1_n13 ), .A2(
        SubCellInst2_LFInst_1_LFInst_1_n12 ), .ZN(
        SubCellInst2_LFInst_1_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_1_U6  ( .A1(SubCellInput[4]), .A2(
        SubCellInput[6]), .ZN(SubCellInst2_LFInst_1_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_1_U5  ( .A1(
        SubCellInst2_LFInst_1_LFInst_1_n11 ), .A2(
        SubCellInst2_LFInst_1_LFInst_1_n10 ), .ZN(
        SubCellInst2_LFInst_1_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_1_U4  ( .A1(SubCellInput[4]), .A2(
        SubCellInput[5]), .ZN(SubCellInst2_LFInst_1_LFInst_1_n10 ) );
  INV_X1 SubCellInst2_LFInst_1_LFInst_1_U3  ( .A(SubCellInput[6]), .ZN(
        SubCellInst2_LFInst_1_LFInst_1_n11 ) );
  XNOR2_X1 SubCellInst2_LFInst_1_LFInst_0_U6  ( .A(
        SubCellInst2_LFInst_1_LFInst_0_n6 ), .B(
        SubCellInst2_LFInst_1_LFInst_0_n5 ), .ZN(MCInst2_MC3_v3_2 [3]) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_0_U5  ( .A1(SubCellInput[6]), .A2(
        SubCellInst2_LFInst_1_LFInst_0_n4 ), .ZN(
        SubCellInst2_LFInst_1_LFInst_0_n5 ) );
  INV_X1 SubCellInst2_LFInst_1_LFInst_0_U4  ( .A(SubCellInput[5]), .ZN(
        SubCellInst2_LFInst_1_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst2_LFInst_1_LFInst_0_U3  ( .A(SubCellInput[4]), .B(
        SubCellInput[7]), .Z(SubCellInst2_LFInst_1_LFInst_0_n6 ) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_3_U9  ( .A1(
        SubCellInst2_LFInst_2_LFInst_3_n16 ), .A2(
        SubCellInst2_LFInst_2_LFInst_3_n15 ), .ZN(MCInst2_MC2_v3_2 [2]) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_3_U8  ( .A1(SubCellInput[9]), .A2(
        SubCellInst2_LFInst_2_LFInst_3_n14 ), .ZN(
        SubCellInst2_LFInst_2_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst2_LFInst_2_LFInst_3_U7  ( .A(SubCellInput[11]), .B(
        SubCellInput[10]), .Z(SubCellInst2_LFInst_2_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_3_U6  ( .A1(
        SubCellInst2_LFInst_2_LFInst_3_n13 ), .A2(
        SubCellInst2_LFInst_2_LFInst_3_n12 ), .ZN(
        SubCellInst2_LFInst_2_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_3_U5  ( .A1(SubCellInput[8]), .A2(
        SubCellInput[10]), .ZN(SubCellInst2_LFInst_2_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst2_LFInst_2_LFInst_3_U4  ( .A(SubCellInput[8]), .B(
        SubCellInst2_LFInst_2_LFInst_3_n11 ), .ZN(
        SubCellInst2_LFInst_2_LFInst_3_n13 ) );
  OR2_X1 SubCellInst2_LFInst_2_LFInst_3_U3  ( .A1(SubCellInput[11]), .A2(
        SubCellInput[9]), .ZN(SubCellInst2_LFInst_2_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_2_U11  ( .A1(
        SubCellInst2_LFInst_2_LFInst_2_n22 ), .A2(
        SubCellInst2_LFInst_2_LFInst_2_n21 ), .ZN(MCInst2_MC2_v3_0 [3]) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_2_U10  ( .A1(SubCellInput[10]), .A2(
        SubCellInst2_LFInst_2_LFInst_2_n20 ), .ZN(
        SubCellInst2_LFInst_2_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst2_LFInst_2_LFInst_2_U9  ( .A1(SubCellInput[9]), .A2(
        SubCellInst2_LFInst_2_LFInst_2_n19 ), .ZN(
        SubCellInst2_LFInst_2_LFInst_2_n20 ) );
  INV_X1 SubCellInst2_LFInst_2_LFInst_2_U8  ( .A(SubCellInput[11]), .ZN(
        SubCellInst2_LFInst_2_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_2_U7  ( .A1(
        SubCellInst2_LFInst_2_LFInst_2_n18 ), .A2(
        SubCellInst2_LFInst_2_LFInst_2_n17 ), .ZN(
        SubCellInst2_LFInst_2_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst2_LFInst_2_LFInst_2_U6  ( .A(
        SubCellInst2_LFInst_2_LFInst_2_n16 ), .B(SubCellInput[10]), .Z(
        SubCellInst2_LFInst_2_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_2_U5  ( .A1(SubCellInput[8]), .A2(
        SubCellInput[9]), .ZN(SubCellInst2_LFInst_2_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_2_U4  ( .A1(
        SubCellInst2_LFInst_2_LFInst_2_n15 ), .A2(SubCellInput[11]), .ZN(
        SubCellInst2_LFInst_2_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst2_LFInst_2_LFInst_2_U3  ( .A(SubCellInput[8]), .B(
        SubCellInput[9]), .ZN(SubCellInst2_LFInst_2_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_1_U12  ( .A1(
        SubCellInst2_LFInst_2_LFInst_1_n18 ), .A2(
        SubCellInst2_LFInst_2_LFInst_1_n17 ), .ZN(MCInst2_MC2_v3_0 [2]) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_1_U11  ( .A1(SubCellInput[9]), .A2(
        SubCellInst2_LFInst_2_LFInst_1_n16 ), .ZN(
        SubCellInst2_LFInst_2_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst2_LFInst_2_LFInst_1_U10  ( .A1(SubCellInput[11]), .A2(
        SubCellInst2_LFInst_2_LFInst_1_n15 ), .ZN(
        SubCellInst2_LFInst_2_LFInst_1_n16 ) );
  AND2_X1 SubCellInst2_LFInst_2_LFInst_1_U9  ( .A1(SubCellInput[8]), .A2(
        SubCellInput[10]), .ZN(SubCellInst2_LFInst_2_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_1_U8  ( .A1(SubCellInput[11]), .A2(
        SubCellInst2_LFInst_2_LFInst_1_n14 ), .ZN(
        SubCellInst2_LFInst_2_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_1_U7  ( .A1(
        SubCellInst2_LFInst_2_LFInst_1_n13 ), .A2(
        SubCellInst2_LFInst_2_LFInst_1_n12 ), .ZN(
        SubCellInst2_LFInst_2_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_1_U6  ( .A1(SubCellInput[8]), .A2(
        SubCellInput[10]), .ZN(SubCellInst2_LFInst_2_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_1_U5  ( .A1(
        SubCellInst2_LFInst_2_LFInst_1_n11 ), .A2(
        SubCellInst2_LFInst_2_LFInst_1_n10 ), .ZN(
        SubCellInst2_LFInst_2_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_1_U4  ( .A1(SubCellInput[8]), .A2(
        SubCellInput[9]), .ZN(SubCellInst2_LFInst_2_LFInst_1_n10 ) );
  INV_X1 SubCellInst2_LFInst_2_LFInst_1_U3  ( .A(SubCellInput[10]), .ZN(
        SubCellInst2_LFInst_2_LFInst_1_n11 ) );
  XNOR2_X1 SubCellInst2_LFInst_2_LFInst_0_U6  ( .A(
        SubCellInst2_LFInst_2_LFInst_0_n6 ), .B(
        SubCellInst2_LFInst_2_LFInst_0_n5 ), .ZN(MCInst2_MC2_v3_2 [3]) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_0_U5  ( .A1(SubCellInput[10]), .A2(
        SubCellInst2_LFInst_2_LFInst_0_n4 ), .ZN(
        SubCellInst2_LFInst_2_LFInst_0_n5 ) );
  INV_X1 SubCellInst2_LFInst_2_LFInst_0_U4  ( .A(SubCellInput[9]), .ZN(
        SubCellInst2_LFInst_2_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst2_LFInst_2_LFInst_0_U3  ( .A(SubCellInput[8]), .B(
        SubCellInput[11]), .Z(SubCellInst2_LFInst_2_LFInst_0_n6 ) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_3_U9  ( .A1(
        SubCellInst2_LFInst_3_LFInst_3_n16 ), .A2(
        SubCellInst2_LFInst_3_LFInst_3_n15 ), .ZN(MCInst2_MC1_v3_2 [2]) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_3_U8  ( .A1(SubCellInput[13]), .A2(
        SubCellInst2_LFInst_3_LFInst_3_n14 ), .ZN(
        SubCellInst2_LFInst_3_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst2_LFInst_3_LFInst_3_U7  ( .A(SubCellInput[15]), .B(
        SubCellInput[14]), .Z(SubCellInst2_LFInst_3_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_3_U6  ( .A1(
        SubCellInst2_LFInst_3_LFInst_3_n13 ), .A2(
        SubCellInst2_LFInst_3_LFInst_3_n12 ), .ZN(
        SubCellInst2_LFInst_3_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_3_U5  ( .A1(SubCellInput[12]), .A2(
        SubCellInput[14]), .ZN(SubCellInst2_LFInst_3_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst2_LFInst_3_LFInst_3_U4  ( .A(SubCellInput[12]), .B(
        SubCellInst2_LFInst_3_LFInst_3_n11 ), .ZN(
        SubCellInst2_LFInst_3_LFInst_3_n13 ) );
  OR2_X1 SubCellInst2_LFInst_3_LFInst_3_U3  ( .A1(SubCellInput[15]), .A2(
        SubCellInput[13]), .ZN(SubCellInst2_LFInst_3_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_2_U11  ( .A1(
        SubCellInst2_LFInst_3_LFInst_2_n22 ), .A2(
        SubCellInst2_LFInst_3_LFInst_2_n21 ), .ZN(MCInst2_MC1_v3_0 [3]) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_2_U10  ( .A1(SubCellInput[14]), .A2(
        SubCellInst2_LFInst_3_LFInst_2_n20 ), .ZN(
        SubCellInst2_LFInst_3_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst2_LFInst_3_LFInst_2_U9  ( .A1(SubCellInput[13]), .A2(
        SubCellInst2_LFInst_3_LFInst_2_n19 ), .ZN(
        SubCellInst2_LFInst_3_LFInst_2_n20 ) );
  INV_X1 SubCellInst2_LFInst_3_LFInst_2_U8  ( .A(SubCellInput[15]), .ZN(
        SubCellInst2_LFInst_3_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_2_U7  ( .A1(
        SubCellInst2_LFInst_3_LFInst_2_n18 ), .A2(
        SubCellInst2_LFInst_3_LFInst_2_n17 ), .ZN(
        SubCellInst2_LFInst_3_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst2_LFInst_3_LFInst_2_U6  ( .A(
        SubCellInst2_LFInst_3_LFInst_2_n16 ), .B(SubCellInput[14]), .Z(
        SubCellInst2_LFInst_3_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_2_U5  ( .A1(SubCellInput[12]), .A2(
        SubCellInput[13]), .ZN(SubCellInst2_LFInst_3_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_2_U4  ( .A1(
        SubCellInst2_LFInst_3_LFInst_2_n15 ), .A2(SubCellInput[15]), .ZN(
        SubCellInst2_LFInst_3_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst2_LFInst_3_LFInst_2_U3  ( .A(SubCellInput[12]), .B(
        SubCellInput[13]), .ZN(SubCellInst2_LFInst_3_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_1_U12  ( .A1(
        SubCellInst2_LFInst_3_LFInst_1_n18 ), .A2(
        SubCellInst2_LFInst_3_LFInst_1_n17 ), .ZN(MCInst2_MC1_v3_0 [2]) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_1_U11  ( .A1(SubCellInput[13]), .A2(
        SubCellInst2_LFInst_3_LFInst_1_n16 ), .ZN(
        SubCellInst2_LFInst_3_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst2_LFInst_3_LFInst_1_U10  ( .A1(SubCellInput[15]), .A2(
        SubCellInst2_LFInst_3_LFInst_1_n15 ), .ZN(
        SubCellInst2_LFInst_3_LFInst_1_n16 ) );
  AND2_X1 SubCellInst2_LFInst_3_LFInst_1_U9  ( .A1(SubCellInput[12]), .A2(
        SubCellInput[14]), .ZN(SubCellInst2_LFInst_3_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_1_U8  ( .A1(SubCellInput[15]), .A2(
        SubCellInst2_LFInst_3_LFInst_1_n14 ), .ZN(
        SubCellInst2_LFInst_3_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_1_U7  ( .A1(
        SubCellInst2_LFInst_3_LFInst_1_n13 ), .A2(
        SubCellInst2_LFInst_3_LFInst_1_n12 ), .ZN(
        SubCellInst2_LFInst_3_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_1_U6  ( .A1(SubCellInput[12]), .A2(
        SubCellInput[14]), .ZN(SubCellInst2_LFInst_3_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_1_U5  ( .A1(
        SubCellInst2_LFInst_3_LFInst_1_n11 ), .A2(
        SubCellInst2_LFInst_3_LFInst_1_n10 ), .ZN(
        SubCellInst2_LFInst_3_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_1_U4  ( .A1(SubCellInput[12]), .A2(
        SubCellInput[13]), .ZN(SubCellInst2_LFInst_3_LFInst_1_n10 ) );
  INV_X1 SubCellInst2_LFInst_3_LFInst_1_U3  ( .A(SubCellInput[14]), .ZN(
        SubCellInst2_LFInst_3_LFInst_1_n11 ) );
  XNOR2_X1 SubCellInst2_LFInst_3_LFInst_0_U6  ( .A(
        SubCellInst2_LFInst_3_LFInst_0_n6 ), .B(
        SubCellInst2_LFInst_3_LFInst_0_n5 ), .ZN(MCInst2_MC1_v3_2 [3]) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_0_U5  ( .A1(SubCellInput[14]), .A2(
        SubCellInst2_LFInst_3_LFInst_0_n4 ), .ZN(
        SubCellInst2_LFInst_3_LFInst_0_n5 ) );
  INV_X1 SubCellInst2_LFInst_3_LFInst_0_U4  ( .A(SubCellInput[13]), .ZN(
        SubCellInst2_LFInst_3_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst2_LFInst_3_LFInst_0_U3  ( .A(SubCellInput[12]), .B(
        SubCellInput[15]), .Z(SubCellInst2_LFInst_3_LFInst_0_n6 ) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_3_U9  ( .A1(
        SubCellInst2_LFInst_4_LFInst_3_n16 ), .A2(
        SubCellInst2_LFInst_4_LFInst_3_n15 ), .ZN(MCInst2_MC1_v2_0 [0]) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_3_U8  ( .A1(SubCellInput[17]), .A2(
        SubCellInst2_LFInst_4_LFInst_3_n14 ), .ZN(
        SubCellInst2_LFInst_4_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst2_LFInst_4_LFInst_3_U7  ( .A(SubCellInput[19]), .B(
        SubCellInput[18]), .Z(SubCellInst2_LFInst_4_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_3_U6  ( .A1(
        SubCellInst2_LFInst_4_LFInst_3_n13 ), .A2(
        SubCellInst2_LFInst_4_LFInst_3_n12 ), .ZN(
        SubCellInst2_LFInst_4_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_3_U5  ( .A1(SubCellInput[16]), .A2(
        SubCellInput[18]), .ZN(SubCellInst2_LFInst_4_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst2_LFInst_4_LFInst_3_U4  ( .A(SubCellInput[16]), .B(
        SubCellInst2_LFInst_4_LFInst_3_n11 ), .ZN(
        SubCellInst2_LFInst_4_LFInst_3_n13 ) );
  OR2_X1 SubCellInst2_LFInst_4_LFInst_3_U3  ( .A1(SubCellInput[19]), .A2(
        SubCellInput[17]), .ZN(SubCellInst2_LFInst_4_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_2_U11  ( .A1(
        SubCellInst2_LFInst_4_LFInst_2_n22 ), .A2(
        SubCellInst2_LFInst_4_LFInst_2_n21 ), .ZN(MCInst2_MC1_v2_0 [3]) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_2_U10  ( .A1(SubCellInput[18]), .A2(
        SubCellInst2_LFInst_4_LFInst_2_n20 ), .ZN(
        SubCellInst2_LFInst_4_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst2_LFInst_4_LFInst_2_U9  ( .A1(SubCellInput[17]), .A2(
        SubCellInst2_LFInst_4_LFInst_2_n19 ), .ZN(
        SubCellInst2_LFInst_4_LFInst_2_n20 ) );
  INV_X1 SubCellInst2_LFInst_4_LFInst_2_U8  ( .A(SubCellInput[19]), .ZN(
        SubCellInst2_LFInst_4_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_2_U7  ( .A1(
        SubCellInst2_LFInst_4_LFInst_2_n18 ), .A2(
        SubCellInst2_LFInst_4_LFInst_2_n17 ), .ZN(
        SubCellInst2_LFInst_4_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst2_LFInst_4_LFInst_2_U6  ( .A(
        SubCellInst2_LFInst_4_LFInst_2_n16 ), .B(SubCellInput[18]), .Z(
        SubCellInst2_LFInst_4_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_2_U5  ( .A1(SubCellInput[16]), .A2(
        SubCellInput[17]), .ZN(SubCellInst2_LFInst_4_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_2_U4  ( .A1(
        SubCellInst2_LFInst_4_LFInst_2_n15 ), .A2(SubCellInput[19]), .ZN(
        SubCellInst2_LFInst_4_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst2_LFInst_4_LFInst_2_U3  ( .A(SubCellInput[16]), .B(
        SubCellInput[17]), .ZN(SubCellInst2_LFInst_4_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_1_U12  ( .A1(
        SubCellInst2_LFInst_4_LFInst_1_n18 ), .A2(
        SubCellInst2_LFInst_4_LFInst_1_n17 ), .ZN(MCInst2_MC1_v2_0 [2]) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_1_U11  ( .A1(SubCellInput[17]), .A2(
        SubCellInst2_LFInst_4_LFInst_1_n16 ), .ZN(
        SubCellInst2_LFInst_4_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst2_LFInst_4_LFInst_1_U10  ( .A1(SubCellInput[19]), .A2(
        SubCellInst2_LFInst_4_LFInst_1_n15 ), .ZN(
        SubCellInst2_LFInst_4_LFInst_1_n16 ) );
  AND2_X1 SubCellInst2_LFInst_4_LFInst_1_U9  ( .A1(SubCellInput[16]), .A2(
        SubCellInput[18]), .ZN(SubCellInst2_LFInst_4_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_1_U8  ( .A1(SubCellInput[19]), .A2(
        SubCellInst2_LFInst_4_LFInst_1_n14 ), .ZN(
        SubCellInst2_LFInst_4_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_1_U7  ( .A1(
        SubCellInst2_LFInst_4_LFInst_1_n13 ), .A2(
        SubCellInst2_LFInst_4_LFInst_1_n12 ), .ZN(
        SubCellInst2_LFInst_4_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_1_U6  ( .A1(SubCellInput[16]), .A2(
        SubCellInput[18]), .ZN(SubCellInst2_LFInst_4_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_1_U5  ( .A1(
        SubCellInst2_LFInst_4_LFInst_1_n11 ), .A2(
        SubCellInst2_LFInst_4_LFInst_1_n10 ), .ZN(
        SubCellInst2_LFInst_4_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_1_U4  ( .A1(SubCellInput[16]), .A2(
        SubCellInput[17]), .ZN(SubCellInst2_LFInst_4_LFInst_1_n10 ) );
  INV_X1 SubCellInst2_LFInst_4_LFInst_1_U3  ( .A(SubCellInput[18]), .ZN(
        SubCellInst2_LFInst_4_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_0_U6  ( .A1(SubCellInput[18]), .A2(
        SubCellInst2_LFInst_4_LFInst_0_n4 ), .ZN(
        SubCellInst2_LFInst_4_LFInst_0_n5 ) );
  INV_X1 SubCellInst2_LFInst_4_LFInst_0_U5  ( .A(SubCellInput[17]), .ZN(
        SubCellInst2_LFInst_4_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst2_LFInst_4_LFInst_0_U4  ( .A(SubCellInput[16]), .B(
        SubCellInput[19]), .Z(SubCellInst2_LFInst_4_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst2_LFInst_4_LFInst_0_U3  ( .A(
        SubCellInst2_LFInst_4_LFInst_0_n6 ), .B(
        SubCellInst2_LFInst_4_LFInst_0_n5 ), .ZN(MCInst2_MC1_v2_3 [1]) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_3_U9  ( .A1(
        SubCellInst2_LFInst_5_LFInst_3_n16 ), .A2(
        SubCellInst2_LFInst_5_LFInst_3_n15 ), .ZN(MCInst2_MC0_v2_0 [0]) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_3_U8  ( .A1(SubCellInput[21]), .A2(
        SubCellInst2_LFInst_5_LFInst_3_n14 ), .ZN(
        SubCellInst2_LFInst_5_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst2_LFInst_5_LFInst_3_U7  ( .A(SubCellInput[23]), .B(
        SubCellInput[22]), .Z(SubCellInst2_LFInst_5_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_3_U6  ( .A1(
        SubCellInst2_LFInst_5_LFInst_3_n13 ), .A2(
        SubCellInst2_LFInst_5_LFInst_3_n12 ), .ZN(
        SubCellInst2_LFInst_5_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_3_U5  ( .A1(SubCellInput[20]), .A2(
        SubCellInput[22]), .ZN(SubCellInst2_LFInst_5_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst2_LFInst_5_LFInst_3_U4  ( .A(SubCellInput[20]), .B(
        SubCellInst2_LFInst_5_LFInst_3_n11 ), .ZN(
        SubCellInst2_LFInst_5_LFInst_3_n13 ) );
  OR2_X1 SubCellInst2_LFInst_5_LFInst_3_U3  ( .A1(SubCellInput[23]), .A2(
        SubCellInput[21]), .ZN(SubCellInst2_LFInst_5_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_2_U11  ( .A1(
        SubCellInst2_LFInst_5_LFInst_2_n22 ), .A2(
        SubCellInst2_LFInst_5_LFInst_2_n21 ), .ZN(MCInst2_MC0_v2_0 [3]) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_2_U10  ( .A1(SubCellInput[22]), .A2(
        SubCellInst2_LFInst_5_LFInst_2_n20 ), .ZN(
        SubCellInst2_LFInst_5_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst2_LFInst_5_LFInst_2_U9  ( .A1(SubCellInput[21]), .A2(
        SubCellInst2_LFInst_5_LFInst_2_n19 ), .ZN(
        SubCellInst2_LFInst_5_LFInst_2_n20 ) );
  INV_X1 SubCellInst2_LFInst_5_LFInst_2_U8  ( .A(SubCellInput[23]), .ZN(
        SubCellInst2_LFInst_5_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_2_U7  ( .A1(
        SubCellInst2_LFInst_5_LFInst_2_n18 ), .A2(
        SubCellInst2_LFInst_5_LFInst_2_n17 ), .ZN(
        SubCellInst2_LFInst_5_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst2_LFInst_5_LFInst_2_U6  ( .A(
        SubCellInst2_LFInst_5_LFInst_2_n16 ), .B(SubCellInput[22]), .Z(
        SubCellInst2_LFInst_5_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_2_U5  ( .A1(SubCellInput[20]), .A2(
        SubCellInput[21]), .ZN(SubCellInst2_LFInst_5_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_2_U4  ( .A1(
        SubCellInst2_LFInst_5_LFInst_2_n15 ), .A2(SubCellInput[23]), .ZN(
        SubCellInst2_LFInst_5_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst2_LFInst_5_LFInst_2_U3  ( .A(SubCellInput[20]), .B(
        SubCellInput[21]), .ZN(SubCellInst2_LFInst_5_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_1_U12  ( .A1(
        SubCellInst2_LFInst_5_LFInst_1_n18 ), .A2(
        SubCellInst2_LFInst_5_LFInst_1_n17 ), .ZN(MCInst2_MC0_v2_0 [2]) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_1_U11  ( .A1(SubCellInput[21]), .A2(
        SubCellInst2_LFInst_5_LFInst_1_n16 ), .ZN(
        SubCellInst2_LFInst_5_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst2_LFInst_5_LFInst_1_U10  ( .A1(SubCellInput[23]), .A2(
        SubCellInst2_LFInst_5_LFInst_1_n15 ), .ZN(
        SubCellInst2_LFInst_5_LFInst_1_n16 ) );
  AND2_X1 SubCellInst2_LFInst_5_LFInst_1_U9  ( .A1(SubCellInput[20]), .A2(
        SubCellInput[22]), .ZN(SubCellInst2_LFInst_5_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_1_U8  ( .A1(SubCellInput[23]), .A2(
        SubCellInst2_LFInst_5_LFInst_1_n14 ), .ZN(
        SubCellInst2_LFInst_5_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_1_U7  ( .A1(
        SubCellInst2_LFInst_5_LFInst_1_n13 ), .A2(
        SubCellInst2_LFInst_5_LFInst_1_n12 ), .ZN(
        SubCellInst2_LFInst_5_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_1_U6  ( .A1(SubCellInput[20]), .A2(
        SubCellInput[22]), .ZN(SubCellInst2_LFInst_5_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_1_U5  ( .A1(
        SubCellInst2_LFInst_5_LFInst_1_n11 ), .A2(
        SubCellInst2_LFInst_5_LFInst_1_n10 ), .ZN(
        SubCellInst2_LFInst_5_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_1_U4  ( .A1(SubCellInput[20]), .A2(
        SubCellInput[21]), .ZN(SubCellInst2_LFInst_5_LFInst_1_n10 ) );
  INV_X1 SubCellInst2_LFInst_5_LFInst_1_U3  ( .A(SubCellInput[22]), .ZN(
        SubCellInst2_LFInst_5_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_0_U6  ( .A1(SubCellInput[22]), .A2(
        SubCellInst2_LFInst_5_LFInst_0_n4 ), .ZN(
        SubCellInst2_LFInst_5_LFInst_0_n5 ) );
  INV_X1 SubCellInst2_LFInst_5_LFInst_0_U5  ( .A(SubCellInput[21]), .ZN(
        SubCellInst2_LFInst_5_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst2_LFInst_5_LFInst_0_U4  ( .A(SubCellInput[20]), .B(
        SubCellInput[23]), .Z(SubCellInst2_LFInst_5_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst2_LFInst_5_LFInst_0_U3  ( .A(
        SubCellInst2_LFInst_5_LFInst_0_n6 ), .B(
        SubCellInst2_LFInst_5_LFInst_0_n5 ), .ZN(MCInst2_MC0_v2_3 [1]) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_3_U9  ( .A1(
        SubCellInst2_LFInst_6_LFInst_3_n16 ), .A2(
        SubCellInst2_LFInst_6_LFInst_3_n15 ), .ZN(MCInst2_MC3_v2_0 [0]) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_3_U8  ( .A1(SubCellInput[25]), .A2(
        SubCellInst2_LFInst_6_LFInst_3_n14 ), .ZN(
        SubCellInst2_LFInst_6_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst2_LFInst_6_LFInst_3_U7  ( .A(SubCellInput[27]), .B(
        SubCellInput[26]), .Z(SubCellInst2_LFInst_6_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_3_U6  ( .A1(
        SubCellInst2_LFInst_6_LFInst_3_n13 ), .A2(
        SubCellInst2_LFInst_6_LFInst_3_n12 ), .ZN(
        SubCellInst2_LFInst_6_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_3_U5  ( .A1(SubCellInput[24]), .A2(
        SubCellInput[26]), .ZN(SubCellInst2_LFInst_6_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst2_LFInst_6_LFInst_3_U4  ( .A(SubCellInput[24]), .B(
        SubCellInst2_LFInst_6_LFInst_3_n11 ), .ZN(
        SubCellInst2_LFInst_6_LFInst_3_n13 ) );
  OR2_X1 SubCellInst2_LFInst_6_LFInst_3_U3  ( .A1(SubCellInput[27]), .A2(
        SubCellInput[25]), .ZN(SubCellInst2_LFInst_6_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_2_U11  ( .A1(
        SubCellInst2_LFInst_6_LFInst_2_n22 ), .A2(
        SubCellInst2_LFInst_6_LFInst_2_n21 ), .ZN(MCInst2_MC3_v2_0 [3]) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_2_U10  ( .A1(SubCellInput[26]), .A2(
        SubCellInst2_LFInst_6_LFInst_2_n20 ), .ZN(
        SubCellInst2_LFInst_6_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst2_LFInst_6_LFInst_2_U9  ( .A1(SubCellInput[25]), .A2(
        SubCellInst2_LFInst_6_LFInst_2_n19 ), .ZN(
        SubCellInst2_LFInst_6_LFInst_2_n20 ) );
  INV_X1 SubCellInst2_LFInst_6_LFInst_2_U8  ( .A(SubCellInput[27]), .ZN(
        SubCellInst2_LFInst_6_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_2_U7  ( .A1(
        SubCellInst2_LFInst_6_LFInst_2_n18 ), .A2(
        SubCellInst2_LFInst_6_LFInst_2_n17 ), .ZN(
        SubCellInst2_LFInst_6_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst2_LFInst_6_LFInst_2_U6  ( .A(
        SubCellInst2_LFInst_6_LFInst_2_n16 ), .B(SubCellInput[26]), .Z(
        SubCellInst2_LFInst_6_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_2_U5  ( .A1(SubCellInput[24]), .A2(
        SubCellInput[25]), .ZN(SubCellInst2_LFInst_6_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_2_U4  ( .A1(
        SubCellInst2_LFInst_6_LFInst_2_n15 ), .A2(SubCellInput[27]), .ZN(
        SubCellInst2_LFInst_6_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst2_LFInst_6_LFInst_2_U3  ( .A(SubCellInput[24]), .B(
        SubCellInput[25]), .ZN(SubCellInst2_LFInst_6_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_1_U12  ( .A1(
        SubCellInst2_LFInst_6_LFInst_1_n18 ), .A2(
        SubCellInst2_LFInst_6_LFInst_1_n17 ), .ZN(MCInst2_MC3_v2_0 [2]) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_1_U11  ( .A1(SubCellInput[25]), .A2(
        SubCellInst2_LFInst_6_LFInst_1_n16 ), .ZN(
        SubCellInst2_LFInst_6_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst2_LFInst_6_LFInst_1_U10  ( .A1(SubCellInput[27]), .A2(
        SubCellInst2_LFInst_6_LFInst_1_n15 ), .ZN(
        SubCellInst2_LFInst_6_LFInst_1_n16 ) );
  AND2_X1 SubCellInst2_LFInst_6_LFInst_1_U9  ( .A1(SubCellInput[24]), .A2(
        SubCellInput[26]), .ZN(SubCellInst2_LFInst_6_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_1_U8  ( .A1(SubCellInput[27]), .A2(
        SubCellInst2_LFInst_6_LFInst_1_n14 ), .ZN(
        SubCellInst2_LFInst_6_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_1_U7  ( .A1(
        SubCellInst2_LFInst_6_LFInst_1_n13 ), .A2(
        SubCellInst2_LFInst_6_LFInst_1_n12 ), .ZN(
        SubCellInst2_LFInst_6_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_1_U6  ( .A1(SubCellInput[24]), .A2(
        SubCellInput[26]), .ZN(SubCellInst2_LFInst_6_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_1_U5  ( .A1(
        SubCellInst2_LFInst_6_LFInst_1_n11 ), .A2(
        SubCellInst2_LFInst_6_LFInst_1_n10 ), .ZN(
        SubCellInst2_LFInst_6_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_1_U4  ( .A1(SubCellInput[24]), .A2(
        SubCellInput[25]), .ZN(SubCellInst2_LFInst_6_LFInst_1_n10 ) );
  INV_X1 SubCellInst2_LFInst_6_LFInst_1_U3  ( .A(SubCellInput[26]), .ZN(
        SubCellInst2_LFInst_6_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_0_U6  ( .A1(SubCellInput[26]), .A2(
        SubCellInst2_LFInst_6_LFInst_0_n4 ), .ZN(
        SubCellInst2_LFInst_6_LFInst_0_n5 ) );
  INV_X1 SubCellInst2_LFInst_6_LFInst_0_U5  ( .A(SubCellInput[25]), .ZN(
        SubCellInst2_LFInst_6_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst2_LFInst_6_LFInst_0_U4  ( .A(SubCellInput[24]), .B(
        SubCellInput[27]), .Z(SubCellInst2_LFInst_6_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst2_LFInst_6_LFInst_0_U3  ( .A(
        SubCellInst2_LFInst_6_LFInst_0_n6 ), .B(
        SubCellInst2_LFInst_6_LFInst_0_n5 ), .ZN(MCInst2_MC3_v2_3 [1]) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_3_U9  ( .A1(
        SubCellInst2_LFInst_7_LFInst_3_n16 ), .A2(
        SubCellInst2_LFInst_7_LFInst_3_n15 ), .ZN(MCInst2_MC2_v2_0 [0]) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_3_U8  ( .A1(SubCellInput[29]), .A2(
        SubCellInst2_LFInst_7_LFInst_3_n14 ), .ZN(
        SubCellInst2_LFInst_7_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst2_LFInst_7_LFInst_3_U7  ( .A(SubCellInput[31]), .B(
        SubCellInput[30]), .Z(SubCellInst2_LFInst_7_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_3_U6  ( .A1(
        SubCellInst2_LFInst_7_LFInst_3_n13 ), .A2(
        SubCellInst2_LFInst_7_LFInst_3_n12 ), .ZN(
        SubCellInst2_LFInst_7_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_3_U5  ( .A1(SubCellInput[28]), .A2(
        SubCellInput[30]), .ZN(SubCellInst2_LFInst_7_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst2_LFInst_7_LFInst_3_U4  ( .A(SubCellInput[28]), .B(
        SubCellInst2_LFInst_7_LFInst_3_n11 ), .ZN(
        SubCellInst2_LFInst_7_LFInst_3_n13 ) );
  OR2_X1 SubCellInst2_LFInst_7_LFInst_3_U3  ( .A1(SubCellInput[31]), .A2(
        SubCellInput[29]), .ZN(SubCellInst2_LFInst_7_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_2_U11  ( .A1(
        SubCellInst2_LFInst_7_LFInst_2_n22 ), .A2(
        SubCellInst2_LFInst_7_LFInst_2_n21 ), .ZN(MCInst2_MC2_v2_0 [3]) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_2_U10  ( .A1(SubCellInput[30]), .A2(
        SubCellInst2_LFInst_7_LFInst_2_n20 ), .ZN(
        SubCellInst2_LFInst_7_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst2_LFInst_7_LFInst_2_U9  ( .A1(SubCellInput[29]), .A2(
        SubCellInst2_LFInst_7_LFInst_2_n19 ), .ZN(
        SubCellInst2_LFInst_7_LFInst_2_n20 ) );
  INV_X1 SubCellInst2_LFInst_7_LFInst_2_U8  ( .A(SubCellInput[31]), .ZN(
        SubCellInst2_LFInst_7_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_2_U7  ( .A1(
        SubCellInst2_LFInst_7_LFInst_2_n18 ), .A2(
        SubCellInst2_LFInst_7_LFInst_2_n17 ), .ZN(
        SubCellInst2_LFInst_7_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst2_LFInst_7_LFInst_2_U6  ( .A(
        SubCellInst2_LFInst_7_LFInst_2_n16 ), .B(SubCellInput[30]), .Z(
        SubCellInst2_LFInst_7_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_2_U5  ( .A1(SubCellInput[28]), .A2(
        SubCellInput[29]), .ZN(SubCellInst2_LFInst_7_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_2_U4  ( .A1(
        SubCellInst2_LFInst_7_LFInst_2_n15 ), .A2(SubCellInput[31]), .ZN(
        SubCellInst2_LFInst_7_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst2_LFInst_7_LFInst_2_U3  ( .A(SubCellInput[28]), .B(
        SubCellInput[29]), .ZN(SubCellInst2_LFInst_7_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_1_U12  ( .A1(
        SubCellInst2_LFInst_7_LFInst_1_n18 ), .A2(
        SubCellInst2_LFInst_7_LFInst_1_n17 ), .ZN(MCInst2_MC2_v2_0 [2]) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_1_U11  ( .A1(SubCellInput[29]), .A2(
        SubCellInst2_LFInst_7_LFInst_1_n16 ), .ZN(
        SubCellInst2_LFInst_7_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst2_LFInst_7_LFInst_1_U10  ( .A1(SubCellInput[31]), .A2(
        SubCellInst2_LFInst_7_LFInst_1_n15 ), .ZN(
        SubCellInst2_LFInst_7_LFInst_1_n16 ) );
  AND2_X1 SubCellInst2_LFInst_7_LFInst_1_U9  ( .A1(SubCellInput[28]), .A2(
        SubCellInput[30]), .ZN(SubCellInst2_LFInst_7_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_1_U8  ( .A1(SubCellInput[31]), .A2(
        SubCellInst2_LFInst_7_LFInst_1_n14 ), .ZN(
        SubCellInst2_LFInst_7_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_1_U7  ( .A1(
        SubCellInst2_LFInst_7_LFInst_1_n13 ), .A2(
        SubCellInst2_LFInst_7_LFInst_1_n12 ), .ZN(
        SubCellInst2_LFInst_7_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_1_U6  ( .A1(SubCellInput[28]), .A2(
        SubCellInput[30]), .ZN(SubCellInst2_LFInst_7_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_1_U5  ( .A1(
        SubCellInst2_LFInst_7_LFInst_1_n11 ), .A2(
        SubCellInst2_LFInst_7_LFInst_1_n10 ), .ZN(
        SubCellInst2_LFInst_7_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_1_U4  ( .A1(SubCellInput[28]), .A2(
        SubCellInput[29]), .ZN(SubCellInst2_LFInst_7_LFInst_1_n10 ) );
  INV_X1 SubCellInst2_LFInst_7_LFInst_1_U3  ( .A(SubCellInput[30]), .ZN(
        SubCellInst2_LFInst_7_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_0_U6  ( .A1(SubCellInput[30]), .A2(
        SubCellInst2_LFInst_7_LFInst_0_n4 ), .ZN(
        SubCellInst2_LFInst_7_LFInst_0_n5 ) );
  INV_X1 SubCellInst2_LFInst_7_LFInst_0_U5  ( .A(SubCellInput[29]), .ZN(
        SubCellInst2_LFInst_7_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst2_LFInst_7_LFInst_0_U4  ( .A(SubCellInput[28]), .B(
        SubCellInput[31]), .Z(SubCellInst2_LFInst_7_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst2_LFInst_7_LFInst_0_U3  ( .A(
        SubCellInst2_LFInst_7_LFInst_0_n6 ), .B(
        SubCellInst2_LFInst_7_LFInst_0_n5 ), .ZN(MCInst2_MC2_v2_3 [1]) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_3_U9  ( .A1(
        SubCellInst2_LFInst_8_LFInst_3_n16 ), .A2(
        SubCellInst2_LFInst_8_LFInst_3_n15 ), .ZN(MCInst2_MC2_v1_3 [0]) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_3_U8  ( .A1(SubCellInput[33]), .A2(
        SubCellInst2_LFInst_8_LFInst_3_n14 ), .ZN(
        SubCellInst2_LFInst_8_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst2_LFInst_8_LFInst_3_U7  ( .A(SubCellInput[35]), .B(
        SubCellInput[34]), .Z(SubCellInst2_LFInst_8_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_3_U6  ( .A1(
        SubCellInst2_LFInst_8_LFInst_3_n13 ), .A2(
        SubCellInst2_LFInst_8_LFInst_3_n12 ), .ZN(
        SubCellInst2_LFInst_8_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_3_U5  ( .A1(SubCellInput[32]), .A2(
        SubCellInput[34]), .ZN(SubCellInst2_LFInst_8_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst2_LFInst_8_LFInst_3_U4  ( .A(SubCellInput[32]), .B(
        SubCellInst2_LFInst_8_LFInst_3_n11 ), .ZN(
        SubCellInst2_LFInst_8_LFInst_3_n13 ) );
  OR2_X1 SubCellInst2_LFInst_8_LFInst_3_U3  ( .A1(SubCellInput[35]), .A2(
        SubCellInput[33]), .ZN(SubCellInst2_LFInst_8_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_2_U11  ( .A1(
        SubCellInst2_LFInst_8_LFInst_2_n22 ), .A2(
        SubCellInst2_LFInst_8_LFInst_2_n21 ), .ZN(MCInst2_MC2_v1_3 [3]) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_2_U10  ( .A1(SubCellInput[34]), .A2(
        SubCellInst2_LFInst_8_LFInst_2_n20 ), .ZN(
        SubCellInst2_LFInst_8_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst2_LFInst_8_LFInst_2_U9  ( .A1(SubCellInput[33]), .A2(
        SubCellInst2_LFInst_8_LFInst_2_n19 ), .ZN(
        SubCellInst2_LFInst_8_LFInst_2_n20 ) );
  INV_X1 SubCellInst2_LFInst_8_LFInst_2_U8  ( .A(SubCellInput[35]), .ZN(
        SubCellInst2_LFInst_8_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_2_U7  ( .A1(
        SubCellInst2_LFInst_8_LFInst_2_n18 ), .A2(
        SubCellInst2_LFInst_8_LFInst_2_n17 ), .ZN(
        SubCellInst2_LFInst_8_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst2_LFInst_8_LFInst_2_U6  ( .A(
        SubCellInst2_LFInst_8_LFInst_2_n16 ), .B(SubCellInput[34]), .Z(
        SubCellInst2_LFInst_8_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_2_U5  ( .A1(SubCellInput[32]), .A2(
        SubCellInput[33]), .ZN(SubCellInst2_LFInst_8_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_2_U4  ( .A1(
        SubCellInst2_LFInst_8_LFInst_2_n15 ), .A2(SubCellInput[35]), .ZN(
        SubCellInst2_LFInst_8_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst2_LFInst_8_LFInst_2_U3  ( .A(SubCellInput[32]), .B(
        SubCellInput[33]), .ZN(SubCellInst2_LFInst_8_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_1_U12  ( .A1(
        SubCellInst2_LFInst_8_LFInst_1_n18 ), .A2(
        SubCellInst2_LFInst_8_LFInst_1_n17 ), .ZN(MCInst2_MC2_v1_3 [2]) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_1_U11  ( .A1(SubCellInput[33]), .A2(
        SubCellInst2_LFInst_8_LFInst_1_n16 ), .ZN(
        SubCellInst2_LFInst_8_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst2_LFInst_8_LFInst_1_U10  ( .A1(SubCellInput[35]), .A2(
        SubCellInst2_LFInst_8_LFInst_1_n15 ), .ZN(
        SubCellInst2_LFInst_8_LFInst_1_n16 ) );
  AND2_X1 SubCellInst2_LFInst_8_LFInst_1_U9  ( .A1(SubCellInput[32]), .A2(
        SubCellInput[34]), .ZN(SubCellInst2_LFInst_8_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_1_U8  ( .A1(SubCellInput[35]), .A2(
        SubCellInst2_LFInst_8_LFInst_1_n14 ), .ZN(
        SubCellInst2_LFInst_8_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_1_U7  ( .A1(
        SubCellInst2_LFInst_8_LFInst_1_n13 ), .A2(
        SubCellInst2_LFInst_8_LFInst_1_n12 ), .ZN(
        SubCellInst2_LFInst_8_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_1_U6  ( .A1(SubCellInput[32]), .A2(
        SubCellInput[34]), .ZN(SubCellInst2_LFInst_8_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_1_U5  ( .A1(
        SubCellInst2_LFInst_8_LFInst_1_n11 ), .A2(
        SubCellInst2_LFInst_8_LFInst_1_n10 ), .ZN(
        SubCellInst2_LFInst_8_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_1_U4  ( .A1(SubCellInput[32]), .A2(
        SubCellInput[33]), .ZN(SubCellInst2_LFInst_8_LFInst_1_n10 ) );
  INV_X1 SubCellInst2_LFInst_8_LFInst_1_U3  ( .A(SubCellInput[34]), .ZN(
        SubCellInst2_LFInst_8_LFInst_1_n11 ) );
  XNOR2_X1 SubCellInst2_LFInst_8_LFInst_0_U6  ( .A(
        SubCellInst2_LFInst_8_LFInst_0_n6 ), .B(
        SubCellInst2_LFInst_8_LFInst_0_n5 ), .ZN(ShiftRowsOutput2[36]) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_0_U5  ( .A1(SubCellInput[34]), .A2(
        SubCellInst2_LFInst_8_LFInst_0_n4 ), .ZN(
        SubCellInst2_LFInst_8_LFInst_0_n5 ) );
  INV_X1 SubCellInst2_LFInst_8_LFInst_0_U4  ( .A(SubCellInput[33]), .ZN(
        SubCellInst2_LFInst_8_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst2_LFInst_8_LFInst_0_U3  ( .A(SubCellInput[32]), .B(
        SubCellInput[35]), .Z(SubCellInst2_LFInst_8_LFInst_0_n6 ) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_3_U9  ( .A1(
        SubCellInst2_LFInst_9_LFInst_3_n16 ), .A2(
        SubCellInst2_LFInst_9_LFInst_3_n15 ), .ZN(MCInst2_MC1_v1_3 [0]) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_3_U8  ( .A1(SubCellInput[37]), .A2(
        SubCellInst2_LFInst_9_LFInst_3_n14 ), .ZN(
        SubCellInst2_LFInst_9_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst2_LFInst_9_LFInst_3_U7  ( .A(SubCellInput[39]), .B(
        SubCellInput[38]), .Z(SubCellInst2_LFInst_9_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_3_U6  ( .A1(
        SubCellInst2_LFInst_9_LFInst_3_n13 ), .A2(
        SubCellInst2_LFInst_9_LFInst_3_n12 ), .ZN(
        SubCellInst2_LFInst_9_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_3_U5  ( .A1(SubCellInput[36]), .A2(
        SubCellInput[38]), .ZN(SubCellInst2_LFInst_9_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst2_LFInst_9_LFInst_3_U4  ( .A(SubCellInput[36]), .B(
        SubCellInst2_LFInst_9_LFInst_3_n11 ), .ZN(
        SubCellInst2_LFInst_9_LFInst_3_n13 ) );
  OR2_X1 SubCellInst2_LFInst_9_LFInst_3_U3  ( .A1(SubCellInput[39]), .A2(
        SubCellInput[37]), .ZN(SubCellInst2_LFInst_9_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_2_U11  ( .A1(
        SubCellInst2_LFInst_9_LFInst_2_n22 ), .A2(
        SubCellInst2_LFInst_9_LFInst_2_n21 ), .ZN(MCInst2_MC1_v1_3 [3]) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_2_U10  ( .A1(SubCellInput[38]), .A2(
        SubCellInst2_LFInst_9_LFInst_2_n20 ), .ZN(
        SubCellInst2_LFInst_9_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst2_LFInst_9_LFInst_2_U9  ( .A1(SubCellInput[37]), .A2(
        SubCellInst2_LFInst_9_LFInst_2_n19 ), .ZN(
        SubCellInst2_LFInst_9_LFInst_2_n20 ) );
  INV_X1 SubCellInst2_LFInst_9_LFInst_2_U8  ( .A(SubCellInput[39]), .ZN(
        SubCellInst2_LFInst_9_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_2_U7  ( .A1(
        SubCellInst2_LFInst_9_LFInst_2_n18 ), .A2(
        SubCellInst2_LFInst_9_LFInst_2_n17 ), .ZN(
        SubCellInst2_LFInst_9_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst2_LFInst_9_LFInst_2_U6  ( .A(
        SubCellInst2_LFInst_9_LFInst_2_n16 ), .B(SubCellInput[38]), .Z(
        SubCellInst2_LFInst_9_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_2_U5  ( .A1(SubCellInput[36]), .A2(
        SubCellInput[37]), .ZN(SubCellInst2_LFInst_9_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_2_U4  ( .A1(
        SubCellInst2_LFInst_9_LFInst_2_n15 ), .A2(SubCellInput[39]), .ZN(
        SubCellInst2_LFInst_9_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst2_LFInst_9_LFInst_2_U3  ( .A(SubCellInput[36]), .B(
        SubCellInput[37]), .ZN(SubCellInst2_LFInst_9_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_1_U12  ( .A1(
        SubCellInst2_LFInst_9_LFInst_1_n18 ), .A2(
        SubCellInst2_LFInst_9_LFInst_1_n17 ), .ZN(MCInst2_MC1_v1_3 [2]) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_1_U11  ( .A1(SubCellInput[37]), .A2(
        SubCellInst2_LFInst_9_LFInst_1_n16 ), .ZN(
        SubCellInst2_LFInst_9_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst2_LFInst_9_LFInst_1_U10  ( .A1(SubCellInput[39]), .A2(
        SubCellInst2_LFInst_9_LFInst_1_n15 ), .ZN(
        SubCellInst2_LFInst_9_LFInst_1_n16 ) );
  AND2_X1 SubCellInst2_LFInst_9_LFInst_1_U9  ( .A1(SubCellInput[36]), .A2(
        SubCellInput[38]), .ZN(SubCellInst2_LFInst_9_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_1_U8  ( .A1(SubCellInput[39]), .A2(
        SubCellInst2_LFInst_9_LFInst_1_n14 ), .ZN(
        SubCellInst2_LFInst_9_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_1_U7  ( .A1(
        SubCellInst2_LFInst_9_LFInst_1_n13 ), .A2(
        SubCellInst2_LFInst_9_LFInst_1_n12 ), .ZN(
        SubCellInst2_LFInst_9_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_1_U6  ( .A1(SubCellInput[36]), .A2(
        SubCellInput[38]), .ZN(SubCellInst2_LFInst_9_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_1_U5  ( .A1(
        SubCellInst2_LFInst_9_LFInst_1_n11 ), .A2(
        SubCellInst2_LFInst_9_LFInst_1_n10 ), .ZN(
        SubCellInst2_LFInst_9_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_1_U4  ( .A1(SubCellInput[36]), .A2(
        SubCellInput[37]), .ZN(SubCellInst2_LFInst_9_LFInst_1_n10 ) );
  INV_X1 SubCellInst2_LFInst_9_LFInst_1_U3  ( .A(SubCellInput[38]), .ZN(
        SubCellInst2_LFInst_9_LFInst_1_n11 ) );
  XNOR2_X1 SubCellInst2_LFInst_9_LFInst_0_U6  ( .A(
        SubCellInst2_LFInst_9_LFInst_0_n6 ), .B(
        SubCellInst2_LFInst_9_LFInst_0_n5 ), .ZN(ShiftRowsOutput2[40]) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_0_U5  ( .A1(SubCellInput[38]), .A2(
        SubCellInst2_LFInst_9_LFInst_0_n4 ), .ZN(
        SubCellInst2_LFInst_9_LFInst_0_n5 ) );
  INV_X1 SubCellInst2_LFInst_9_LFInst_0_U4  ( .A(SubCellInput[37]), .ZN(
        SubCellInst2_LFInst_9_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst2_LFInst_9_LFInst_0_U3  ( .A(SubCellInput[36]), .B(
        SubCellInput[39]), .Z(SubCellInst2_LFInst_9_LFInst_0_n6 ) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_3_U9  ( .A1(
        SubCellInst2_LFInst_10_LFInst_3_n16 ), .A2(
        SubCellInst2_LFInst_10_LFInst_3_n15 ), .ZN(MCInst2_MC0_v1_3 [0]) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_3_U8  ( .A1(SubCellInput[41]), .A2(
        SubCellInst2_LFInst_10_LFInst_3_n14 ), .ZN(
        SubCellInst2_LFInst_10_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst2_LFInst_10_LFInst_3_U7  ( .A(SubCellInput[43]), .B(
        SubCellInput[42]), .Z(SubCellInst2_LFInst_10_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_3_U6  ( .A1(
        SubCellInst2_LFInst_10_LFInst_3_n13 ), .A2(
        SubCellInst2_LFInst_10_LFInst_3_n12 ), .ZN(
        SubCellInst2_LFInst_10_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_3_U5  ( .A1(SubCellInput[40]), .A2(
        SubCellInput[42]), .ZN(SubCellInst2_LFInst_10_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst2_LFInst_10_LFInst_3_U4  ( .A(SubCellInput[40]), .B(
        SubCellInst2_LFInst_10_LFInst_3_n11 ), .ZN(
        SubCellInst2_LFInst_10_LFInst_3_n13 ) );
  OR2_X1 SubCellInst2_LFInst_10_LFInst_3_U3  ( .A1(SubCellInput[43]), .A2(
        SubCellInput[41]), .ZN(SubCellInst2_LFInst_10_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_2_U11  ( .A1(
        SubCellInst2_LFInst_10_LFInst_2_n22 ), .A2(
        SubCellInst2_LFInst_10_LFInst_2_n21 ), .ZN(MCInst2_MC0_v1_3 [3]) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_2_U10  ( .A1(SubCellInput[42]), .A2(
        SubCellInst2_LFInst_10_LFInst_2_n20 ), .ZN(
        SubCellInst2_LFInst_10_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst2_LFInst_10_LFInst_2_U9  ( .A1(SubCellInput[41]), .A2(
        SubCellInst2_LFInst_10_LFInst_2_n19 ), .ZN(
        SubCellInst2_LFInst_10_LFInst_2_n20 ) );
  INV_X1 SubCellInst2_LFInst_10_LFInst_2_U8  ( .A(SubCellInput[43]), .ZN(
        SubCellInst2_LFInst_10_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_2_U7  ( .A1(
        SubCellInst2_LFInst_10_LFInst_2_n18 ), .A2(
        SubCellInst2_LFInst_10_LFInst_2_n17 ), .ZN(
        SubCellInst2_LFInst_10_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst2_LFInst_10_LFInst_2_U6  ( .A(
        SubCellInst2_LFInst_10_LFInst_2_n16 ), .B(SubCellInput[42]), .Z(
        SubCellInst2_LFInst_10_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_2_U5  ( .A1(SubCellInput[40]), .A2(
        SubCellInput[41]), .ZN(SubCellInst2_LFInst_10_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_2_U4  ( .A1(
        SubCellInst2_LFInst_10_LFInst_2_n15 ), .A2(SubCellInput[43]), .ZN(
        SubCellInst2_LFInst_10_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst2_LFInst_10_LFInst_2_U3  ( .A(SubCellInput[40]), .B(
        SubCellInput[41]), .ZN(SubCellInst2_LFInst_10_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_1_U12  ( .A1(
        SubCellInst2_LFInst_10_LFInst_1_n18 ), .A2(
        SubCellInst2_LFInst_10_LFInst_1_n17 ), .ZN(MCInst2_MC0_v1_3 [2]) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_1_U11  ( .A1(SubCellInput[41]), .A2(
        SubCellInst2_LFInst_10_LFInst_1_n16 ), .ZN(
        SubCellInst2_LFInst_10_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst2_LFInst_10_LFInst_1_U10  ( .A1(SubCellInput[43]), .A2(
        SubCellInst2_LFInst_10_LFInst_1_n15 ), .ZN(
        SubCellInst2_LFInst_10_LFInst_1_n16 ) );
  AND2_X1 SubCellInst2_LFInst_10_LFInst_1_U9  ( .A1(SubCellInput[40]), .A2(
        SubCellInput[42]), .ZN(SubCellInst2_LFInst_10_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_1_U8  ( .A1(SubCellInput[43]), .A2(
        SubCellInst2_LFInst_10_LFInst_1_n14 ), .ZN(
        SubCellInst2_LFInst_10_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_1_U7  ( .A1(
        SubCellInst2_LFInst_10_LFInst_1_n13 ), .A2(
        SubCellInst2_LFInst_10_LFInst_1_n12 ), .ZN(
        SubCellInst2_LFInst_10_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_1_U6  ( .A1(SubCellInput[40]), .A2(
        SubCellInput[42]), .ZN(SubCellInst2_LFInst_10_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_1_U5  ( .A1(
        SubCellInst2_LFInst_10_LFInst_1_n11 ), .A2(
        SubCellInst2_LFInst_10_LFInst_1_n10 ), .ZN(
        SubCellInst2_LFInst_10_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_1_U4  ( .A1(SubCellInput[40]), .A2(
        SubCellInput[41]), .ZN(SubCellInst2_LFInst_10_LFInst_1_n10 ) );
  INV_X1 SubCellInst2_LFInst_10_LFInst_1_U3  ( .A(SubCellInput[42]), .ZN(
        SubCellInst2_LFInst_10_LFInst_1_n11 ) );
  XNOR2_X1 SubCellInst2_LFInst_10_LFInst_0_U6  ( .A(
        SubCellInst2_LFInst_10_LFInst_0_n6 ), .B(
        SubCellInst2_LFInst_10_LFInst_0_n5 ), .ZN(ShiftRowsOutput2[44]) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_0_U5  ( .A1(SubCellInput[42]), .A2(
        SubCellInst2_LFInst_10_LFInst_0_n4 ), .ZN(
        SubCellInst2_LFInst_10_LFInst_0_n5 ) );
  INV_X1 SubCellInst2_LFInst_10_LFInst_0_U4  ( .A(SubCellInput[41]), .ZN(
        SubCellInst2_LFInst_10_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst2_LFInst_10_LFInst_0_U3  ( .A(SubCellInput[40]), .B(
        SubCellInput[43]), .Z(SubCellInst2_LFInst_10_LFInst_0_n6 ) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_3_U9  ( .A1(
        SubCellInst2_LFInst_11_LFInst_3_n16 ), .A2(
        SubCellInst2_LFInst_11_LFInst_3_n15 ), .ZN(MCInst2_MC3_v1_3 [0]) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_3_U8  ( .A1(SubCellInput[45]), .A2(
        SubCellInst2_LFInst_11_LFInst_3_n14 ), .ZN(
        SubCellInst2_LFInst_11_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst2_LFInst_11_LFInst_3_U7  ( .A(SubCellInput[47]), .B(
        SubCellInput[46]), .Z(SubCellInst2_LFInst_11_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_3_U6  ( .A1(
        SubCellInst2_LFInst_11_LFInst_3_n13 ), .A2(
        SubCellInst2_LFInst_11_LFInst_3_n12 ), .ZN(
        SubCellInst2_LFInst_11_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_3_U5  ( .A1(SubCellInput[44]), .A2(
        SubCellInput[46]), .ZN(SubCellInst2_LFInst_11_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst2_LFInst_11_LFInst_3_U4  ( .A(SubCellInput[44]), .B(
        SubCellInst2_LFInst_11_LFInst_3_n11 ), .ZN(
        SubCellInst2_LFInst_11_LFInst_3_n13 ) );
  OR2_X1 SubCellInst2_LFInst_11_LFInst_3_U3  ( .A1(SubCellInput[47]), .A2(
        SubCellInput[45]), .ZN(SubCellInst2_LFInst_11_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_2_U11  ( .A1(
        SubCellInst2_LFInst_11_LFInst_2_n22 ), .A2(
        SubCellInst2_LFInst_11_LFInst_2_n21 ), .ZN(MCInst2_MC3_v1_3 [3]) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_2_U10  ( .A1(SubCellInput[46]), .A2(
        SubCellInst2_LFInst_11_LFInst_2_n20 ), .ZN(
        SubCellInst2_LFInst_11_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst2_LFInst_11_LFInst_2_U9  ( .A1(SubCellInput[45]), .A2(
        SubCellInst2_LFInst_11_LFInst_2_n19 ), .ZN(
        SubCellInst2_LFInst_11_LFInst_2_n20 ) );
  INV_X1 SubCellInst2_LFInst_11_LFInst_2_U8  ( .A(SubCellInput[47]), .ZN(
        SubCellInst2_LFInst_11_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_2_U7  ( .A1(
        SubCellInst2_LFInst_11_LFInst_2_n18 ), .A2(
        SubCellInst2_LFInst_11_LFInst_2_n17 ), .ZN(
        SubCellInst2_LFInst_11_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst2_LFInst_11_LFInst_2_U6  ( .A(
        SubCellInst2_LFInst_11_LFInst_2_n16 ), .B(SubCellInput[46]), .Z(
        SubCellInst2_LFInst_11_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_2_U5  ( .A1(SubCellInput[44]), .A2(
        SubCellInput[45]), .ZN(SubCellInst2_LFInst_11_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_2_U4  ( .A1(
        SubCellInst2_LFInst_11_LFInst_2_n15 ), .A2(SubCellInput[47]), .ZN(
        SubCellInst2_LFInst_11_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst2_LFInst_11_LFInst_2_U3  ( .A(SubCellInput[44]), .B(
        SubCellInput[45]), .ZN(SubCellInst2_LFInst_11_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_1_U12  ( .A1(
        SubCellInst2_LFInst_11_LFInst_1_n18 ), .A2(
        SubCellInst2_LFInst_11_LFInst_1_n17 ), .ZN(MCInst2_MC3_v1_3 [2]) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_1_U11  ( .A1(SubCellInput[45]), .A2(
        SubCellInst2_LFInst_11_LFInst_1_n16 ), .ZN(
        SubCellInst2_LFInst_11_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst2_LFInst_11_LFInst_1_U10  ( .A1(SubCellInput[47]), .A2(
        SubCellInst2_LFInst_11_LFInst_1_n15 ), .ZN(
        SubCellInst2_LFInst_11_LFInst_1_n16 ) );
  AND2_X1 SubCellInst2_LFInst_11_LFInst_1_U9  ( .A1(SubCellInput[44]), .A2(
        SubCellInput[46]), .ZN(SubCellInst2_LFInst_11_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_1_U8  ( .A1(SubCellInput[47]), .A2(
        SubCellInst2_LFInst_11_LFInst_1_n14 ), .ZN(
        SubCellInst2_LFInst_11_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_1_U7  ( .A1(
        SubCellInst2_LFInst_11_LFInst_1_n13 ), .A2(
        SubCellInst2_LFInst_11_LFInst_1_n12 ), .ZN(
        SubCellInst2_LFInst_11_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_1_U6  ( .A1(SubCellInput[44]), .A2(
        SubCellInput[46]), .ZN(SubCellInst2_LFInst_11_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_1_U5  ( .A1(
        SubCellInst2_LFInst_11_LFInst_1_n11 ), .A2(
        SubCellInst2_LFInst_11_LFInst_1_n10 ), .ZN(
        SubCellInst2_LFInst_11_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_1_U4  ( .A1(SubCellInput[44]), .A2(
        SubCellInput[45]), .ZN(SubCellInst2_LFInst_11_LFInst_1_n10 ) );
  INV_X1 SubCellInst2_LFInst_11_LFInst_1_U3  ( .A(SubCellInput[46]), .ZN(
        SubCellInst2_LFInst_11_LFInst_1_n11 ) );
  XNOR2_X1 SubCellInst2_LFInst_11_LFInst_0_U6  ( .A(
        SubCellInst2_LFInst_11_LFInst_0_n6 ), .B(
        SubCellInst2_LFInst_11_LFInst_0_n5 ), .ZN(ShiftRowsOutput2[32]) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_0_U5  ( .A1(SubCellInput[46]), .A2(
        SubCellInst2_LFInst_11_LFInst_0_n4 ), .ZN(
        SubCellInst2_LFInst_11_LFInst_0_n5 ) );
  INV_X1 SubCellInst2_LFInst_11_LFInst_0_U4  ( .A(SubCellInput[45]), .ZN(
        SubCellInst2_LFInst_11_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst2_LFInst_11_LFInst_0_U3  ( .A(SubCellInput[44]), .B(
        SubCellInput[47]), .Z(SubCellInst2_LFInst_11_LFInst_0_n6 ) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_3_U9  ( .A1(
        SubCellInst2_LFInst_12_LFInst_3_n16 ), .A2(
        SubCellInst2_LFInst_12_LFInst_3_n15 ), .ZN(MCInst2_MC3_v0_3 [0]) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_3_U8  ( .A1(SubCellInput[49]), .A2(
        SubCellInst2_LFInst_12_LFInst_3_n14 ), .ZN(
        SubCellInst2_LFInst_12_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst2_LFInst_12_LFInst_3_U7  ( .A(SubCellInput[51]), .B(
        SubCellInput[50]), .Z(SubCellInst2_LFInst_12_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_3_U6  ( .A1(
        SubCellInst2_LFInst_12_LFInst_3_n13 ), .A2(
        SubCellInst2_LFInst_12_LFInst_3_n12 ), .ZN(
        SubCellInst2_LFInst_12_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_3_U5  ( .A1(SubCellInput[48]), .A2(
        SubCellInput[50]), .ZN(SubCellInst2_LFInst_12_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst2_LFInst_12_LFInst_3_U4  ( .A(SubCellInput[48]), .B(
        SubCellInst2_LFInst_12_LFInst_3_n11 ), .ZN(
        SubCellInst2_LFInst_12_LFInst_3_n13 ) );
  OR2_X1 SubCellInst2_LFInst_12_LFInst_3_U3  ( .A1(SubCellInput[51]), .A2(
        SubCellInput[49]), .ZN(SubCellInst2_LFInst_12_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_2_U11  ( .A1(
        SubCellInst2_LFInst_12_LFInst_2_n22 ), .A2(
        SubCellInst2_LFInst_12_LFInst_2_n21 ), .ZN(MCInst2_MC3_v0_3 [3]) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_2_U10  ( .A1(SubCellInput[50]), .A2(
        SubCellInst2_LFInst_12_LFInst_2_n20 ), .ZN(
        SubCellInst2_LFInst_12_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst2_LFInst_12_LFInst_2_U9  ( .A1(SubCellInput[49]), .A2(
        SubCellInst2_LFInst_12_LFInst_2_n19 ), .ZN(
        SubCellInst2_LFInst_12_LFInst_2_n20 ) );
  INV_X1 SubCellInst2_LFInst_12_LFInst_2_U8  ( .A(SubCellInput[51]), .ZN(
        SubCellInst2_LFInst_12_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_2_U7  ( .A1(
        SubCellInst2_LFInst_12_LFInst_2_n18 ), .A2(
        SubCellInst2_LFInst_12_LFInst_2_n17 ), .ZN(
        SubCellInst2_LFInst_12_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst2_LFInst_12_LFInst_2_U6  ( .A(
        SubCellInst2_LFInst_12_LFInst_2_n16 ), .B(SubCellInput[50]), .Z(
        SubCellInst2_LFInst_12_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_2_U5  ( .A1(SubCellInput[48]), .A2(
        SubCellInput[49]), .ZN(SubCellInst2_LFInst_12_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_2_U4  ( .A1(
        SubCellInst2_LFInst_12_LFInst_2_n15 ), .A2(SubCellInput[51]), .ZN(
        SubCellInst2_LFInst_12_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst2_LFInst_12_LFInst_2_U3  ( .A(SubCellInput[48]), .B(
        SubCellInput[49]), .ZN(SubCellInst2_LFInst_12_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_1_U12  ( .A1(
        SubCellInst2_LFInst_12_LFInst_1_n18 ), .A2(
        SubCellInst2_LFInst_12_LFInst_1_n17 ), .ZN(MCInst2_MC3_v0_0 [3]) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_1_U11  ( .A1(SubCellInput[49]), .A2(
        SubCellInst2_LFInst_12_LFInst_1_n16 ), .ZN(
        SubCellInst2_LFInst_12_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst2_LFInst_12_LFInst_1_U10  ( .A1(SubCellInput[51]), .A2(
        SubCellInst2_LFInst_12_LFInst_1_n15 ), .ZN(
        SubCellInst2_LFInst_12_LFInst_1_n16 ) );
  AND2_X1 SubCellInst2_LFInst_12_LFInst_1_U9  ( .A1(SubCellInput[48]), .A2(
        SubCellInput[50]), .ZN(SubCellInst2_LFInst_12_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_1_U8  ( .A1(SubCellInput[51]), .A2(
        SubCellInst2_LFInst_12_LFInst_1_n14 ), .ZN(
        SubCellInst2_LFInst_12_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_1_U7  ( .A1(
        SubCellInst2_LFInst_12_LFInst_1_n13 ), .A2(
        SubCellInst2_LFInst_12_LFInst_1_n12 ), .ZN(
        SubCellInst2_LFInst_12_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_1_U6  ( .A1(SubCellInput[48]), .A2(
        SubCellInput[50]), .ZN(SubCellInst2_LFInst_12_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_1_U5  ( .A1(
        SubCellInst2_LFInst_12_LFInst_1_n11 ), .A2(
        SubCellInst2_LFInst_12_LFInst_1_n10 ), .ZN(
        SubCellInst2_LFInst_12_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_1_U4  ( .A1(SubCellInput[48]), .A2(
        SubCellInput[49]), .ZN(SubCellInst2_LFInst_12_LFInst_1_n10 ) );
  INV_X1 SubCellInst2_LFInst_12_LFInst_1_U3  ( .A(SubCellInput[50]), .ZN(
        SubCellInst2_LFInst_12_LFInst_1_n11 ) );
  XNOR2_X1 SubCellInst2_LFInst_12_LFInst_0_U6  ( .A(
        SubCellInst2_LFInst_12_LFInst_0_n6 ), .B(
        SubCellInst2_LFInst_12_LFInst_0_n5 ), .ZN(ShiftRowsOutput2[48]) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_0_U5  ( .A1(SubCellInput[50]), .A2(
        SubCellInst2_LFInst_12_LFInst_0_n4 ), .ZN(
        SubCellInst2_LFInst_12_LFInst_0_n5 ) );
  INV_X1 SubCellInst2_LFInst_12_LFInst_0_U4  ( .A(SubCellInput[49]), .ZN(
        SubCellInst2_LFInst_12_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst2_LFInst_12_LFInst_0_U3  ( .A(SubCellInput[48]), .B(
        SubCellInput[51]), .Z(SubCellInst2_LFInst_12_LFInst_0_n6 ) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_3_U9  ( .A1(
        SubCellInst2_LFInst_13_LFInst_3_n16 ), .A2(
        SubCellInst2_LFInst_13_LFInst_3_n15 ), .ZN(MCInst2_MC2_v0_3 [0]) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_3_U8  ( .A1(SubCellInput[53]), .A2(
        SubCellInst2_LFInst_13_LFInst_3_n14 ), .ZN(
        SubCellInst2_LFInst_13_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst2_LFInst_13_LFInst_3_U7  ( .A(SubCellInput[55]), .B(
        SubCellInput[54]), .Z(SubCellInst2_LFInst_13_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_3_U6  ( .A1(
        SubCellInst2_LFInst_13_LFInst_3_n13 ), .A2(
        SubCellInst2_LFInst_13_LFInst_3_n12 ), .ZN(
        SubCellInst2_LFInst_13_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_3_U5  ( .A1(SubCellInput[52]), .A2(
        SubCellInput[54]), .ZN(SubCellInst2_LFInst_13_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst2_LFInst_13_LFInst_3_U4  ( .A(SubCellInput[52]), .B(
        SubCellInst2_LFInst_13_LFInst_3_n11 ), .ZN(
        SubCellInst2_LFInst_13_LFInst_3_n13 ) );
  OR2_X1 SubCellInst2_LFInst_13_LFInst_3_U3  ( .A1(SubCellInput[55]), .A2(
        SubCellInput[53]), .ZN(SubCellInst2_LFInst_13_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_2_U11  ( .A1(
        SubCellInst2_LFInst_13_LFInst_2_n22 ), .A2(
        SubCellInst2_LFInst_13_LFInst_2_n21 ), .ZN(MCInst2_MC2_v0_3 [3]) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_2_U10  ( .A1(SubCellInput[54]), .A2(
        SubCellInst2_LFInst_13_LFInst_2_n20 ), .ZN(
        SubCellInst2_LFInst_13_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst2_LFInst_13_LFInst_2_U9  ( .A1(SubCellInput[53]), .A2(
        SubCellInst2_LFInst_13_LFInst_2_n19 ), .ZN(
        SubCellInst2_LFInst_13_LFInst_2_n20 ) );
  INV_X1 SubCellInst2_LFInst_13_LFInst_2_U8  ( .A(SubCellInput[55]), .ZN(
        SubCellInst2_LFInst_13_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_2_U7  ( .A1(
        SubCellInst2_LFInst_13_LFInst_2_n18 ), .A2(
        SubCellInst2_LFInst_13_LFInst_2_n17 ), .ZN(
        SubCellInst2_LFInst_13_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst2_LFInst_13_LFInst_2_U6  ( .A(
        SubCellInst2_LFInst_13_LFInst_2_n16 ), .B(SubCellInput[54]), .Z(
        SubCellInst2_LFInst_13_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_2_U5  ( .A1(SubCellInput[52]), .A2(
        SubCellInput[53]), .ZN(SubCellInst2_LFInst_13_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_2_U4  ( .A1(
        SubCellInst2_LFInst_13_LFInst_2_n15 ), .A2(SubCellInput[55]), .ZN(
        SubCellInst2_LFInst_13_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst2_LFInst_13_LFInst_2_U3  ( .A(SubCellInput[52]), .B(
        SubCellInput[53]), .ZN(SubCellInst2_LFInst_13_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_1_U12  ( .A1(
        SubCellInst2_LFInst_13_LFInst_1_n18 ), .A2(
        SubCellInst2_LFInst_13_LFInst_1_n17 ), .ZN(MCInst2_MC2_v0_0 [3]) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_1_U11  ( .A1(SubCellInput[53]), .A2(
        SubCellInst2_LFInst_13_LFInst_1_n16 ), .ZN(
        SubCellInst2_LFInst_13_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst2_LFInst_13_LFInst_1_U10  ( .A1(SubCellInput[55]), .A2(
        SubCellInst2_LFInst_13_LFInst_1_n15 ), .ZN(
        SubCellInst2_LFInst_13_LFInst_1_n16 ) );
  AND2_X1 SubCellInst2_LFInst_13_LFInst_1_U9  ( .A1(SubCellInput[52]), .A2(
        SubCellInput[54]), .ZN(SubCellInst2_LFInst_13_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_1_U8  ( .A1(SubCellInput[55]), .A2(
        SubCellInst2_LFInst_13_LFInst_1_n14 ), .ZN(
        SubCellInst2_LFInst_13_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_1_U7  ( .A1(
        SubCellInst2_LFInst_13_LFInst_1_n13 ), .A2(
        SubCellInst2_LFInst_13_LFInst_1_n12 ), .ZN(
        SubCellInst2_LFInst_13_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_1_U6  ( .A1(SubCellInput[52]), .A2(
        SubCellInput[54]), .ZN(SubCellInst2_LFInst_13_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_1_U5  ( .A1(
        SubCellInst2_LFInst_13_LFInst_1_n11 ), .A2(
        SubCellInst2_LFInst_13_LFInst_1_n10 ), .ZN(
        SubCellInst2_LFInst_13_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_1_U4  ( .A1(SubCellInput[52]), .A2(
        SubCellInput[53]), .ZN(SubCellInst2_LFInst_13_LFInst_1_n10 ) );
  INV_X1 SubCellInst2_LFInst_13_LFInst_1_U3  ( .A(SubCellInput[54]), .ZN(
        SubCellInst2_LFInst_13_LFInst_1_n11 ) );
  XNOR2_X1 SubCellInst2_LFInst_13_LFInst_0_U6  ( .A(
        SubCellInst2_LFInst_13_LFInst_0_n6 ), .B(
        SubCellInst2_LFInst_13_LFInst_0_n5 ), .ZN(ShiftRowsOutput2[52]) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_0_U5  ( .A1(SubCellInput[54]), .A2(
        SubCellInst2_LFInst_13_LFInst_0_n4 ), .ZN(
        SubCellInst2_LFInst_13_LFInst_0_n5 ) );
  INV_X1 SubCellInst2_LFInst_13_LFInst_0_U4  ( .A(SubCellInput[53]), .ZN(
        SubCellInst2_LFInst_13_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst2_LFInst_13_LFInst_0_U3  ( .A(SubCellInput[52]), .B(
        SubCellInput[55]), .Z(SubCellInst2_LFInst_13_LFInst_0_n6 ) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_3_U9  ( .A1(
        SubCellInst2_LFInst_14_LFInst_3_n16 ), .A2(
        SubCellInst2_LFInst_14_LFInst_3_n15 ), .ZN(MCInst2_MC1_v0_3 [0]) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_3_U8  ( .A1(SubCellInput[57]), .A2(
        SubCellInst2_LFInst_14_LFInst_3_n14 ), .ZN(
        SubCellInst2_LFInst_14_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst2_LFInst_14_LFInst_3_U7  ( .A(SubCellInput[59]), .B(
        SubCellInput[58]), .Z(SubCellInst2_LFInst_14_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_3_U6  ( .A1(
        SubCellInst2_LFInst_14_LFInst_3_n13 ), .A2(
        SubCellInst2_LFInst_14_LFInst_3_n12 ), .ZN(
        SubCellInst2_LFInst_14_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_3_U5  ( .A1(SubCellInput[56]), .A2(
        SubCellInput[58]), .ZN(SubCellInst2_LFInst_14_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst2_LFInst_14_LFInst_3_U4  ( .A(SubCellInput[56]), .B(
        SubCellInst2_LFInst_14_LFInst_3_n11 ), .ZN(
        SubCellInst2_LFInst_14_LFInst_3_n13 ) );
  OR2_X1 SubCellInst2_LFInst_14_LFInst_3_U3  ( .A1(SubCellInput[59]), .A2(
        SubCellInput[57]), .ZN(SubCellInst2_LFInst_14_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_2_U11  ( .A1(
        SubCellInst2_LFInst_14_LFInst_2_n22 ), .A2(
        SubCellInst2_LFInst_14_LFInst_2_n21 ), .ZN(MCInst2_MC1_v0_3 [3]) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_2_U10  ( .A1(SubCellInput[58]), .A2(
        SubCellInst2_LFInst_14_LFInst_2_n20 ), .ZN(
        SubCellInst2_LFInst_14_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst2_LFInst_14_LFInst_2_U9  ( .A1(SubCellInput[57]), .A2(
        SubCellInst2_LFInst_14_LFInst_2_n19 ), .ZN(
        SubCellInst2_LFInst_14_LFInst_2_n20 ) );
  INV_X1 SubCellInst2_LFInst_14_LFInst_2_U8  ( .A(SubCellInput[59]), .ZN(
        SubCellInst2_LFInst_14_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_2_U7  ( .A1(
        SubCellInst2_LFInst_14_LFInst_2_n18 ), .A2(
        SubCellInst2_LFInst_14_LFInst_2_n17 ), .ZN(
        SubCellInst2_LFInst_14_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst2_LFInst_14_LFInst_2_U6  ( .A(
        SubCellInst2_LFInst_14_LFInst_2_n16 ), .B(SubCellInput[58]), .Z(
        SubCellInst2_LFInst_14_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_2_U5  ( .A1(SubCellInput[56]), .A2(
        SubCellInput[57]), .ZN(SubCellInst2_LFInst_14_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_2_U4  ( .A1(
        SubCellInst2_LFInst_14_LFInst_2_n15 ), .A2(SubCellInput[59]), .ZN(
        SubCellInst2_LFInst_14_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst2_LFInst_14_LFInst_2_U3  ( .A(SubCellInput[56]), .B(
        SubCellInput[57]), .ZN(SubCellInst2_LFInst_14_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_1_U12  ( .A1(
        SubCellInst2_LFInst_14_LFInst_1_n18 ), .A2(
        SubCellInst2_LFInst_14_LFInst_1_n17 ), .ZN(MCInst2_MC1_v0_0 [3]) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_1_U11  ( .A1(SubCellInput[57]), .A2(
        SubCellInst2_LFInst_14_LFInst_1_n16 ), .ZN(
        SubCellInst2_LFInst_14_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst2_LFInst_14_LFInst_1_U10  ( .A1(SubCellInput[59]), .A2(
        SubCellInst2_LFInst_14_LFInst_1_n15 ), .ZN(
        SubCellInst2_LFInst_14_LFInst_1_n16 ) );
  AND2_X1 SubCellInst2_LFInst_14_LFInst_1_U9  ( .A1(SubCellInput[56]), .A2(
        SubCellInput[58]), .ZN(SubCellInst2_LFInst_14_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_1_U8  ( .A1(SubCellInput[59]), .A2(
        SubCellInst2_LFInst_14_LFInst_1_n14 ), .ZN(
        SubCellInst2_LFInst_14_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_1_U7  ( .A1(
        SubCellInst2_LFInst_14_LFInst_1_n13 ), .A2(
        SubCellInst2_LFInst_14_LFInst_1_n12 ), .ZN(
        SubCellInst2_LFInst_14_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_1_U6  ( .A1(SubCellInput[56]), .A2(
        SubCellInput[58]), .ZN(SubCellInst2_LFInst_14_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_1_U5  ( .A1(
        SubCellInst2_LFInst_14_LFInst_1_n11 ), .A2(
        SubCellInst2_LFInst_14_LFInst_1_n10 ), .ZN(
        SubCellInst2_LFInst_14_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_1_U4  ( .A1(SubCellInput[56]), .A2(
        SubCellInput[57]), .ZN(SubCellInst2_LFInst_14_LFInst_1_n10 ) );
  INV_X1 SubCellInst2_LFInst_14_LFInst_1_U3  ( .A(SubCellInput[58]), .ZN(
        SubCellInst2_LFInst_14_LFInst_1_n11 ) );
  XNOR2_X1 SubCellInst2_LFInst_14_LFInst_0_U6  ( .A(
        SubCellInst2_LFInst_14_LFInst_0_n6 ), .B(
        SubCellInst2_LFInst_14_LFInst_0_n5 ), .ZN(ShiftRowsOutput2[56]) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_0_U5  ( .A1(SubCellInput[58]), .A2(
        SubCellInst2_LFInst_14_LFInst_0_n4 ), .ZN(
        SubCellInst2_LFInst_14_LFInst_0_n5 ) );
  INV_X1 SubCellInst2_LFInst_14_LFInst_0_U4  ( .A(SubCellInput[57]), .ZN(
        SubCellInst2_LFInst_14_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst2_LFInst_14_LFInst_0_U3  ( .A(SubCellInput[56]), .B(
        SubCellInput[59]), .Z(SubCellInst2_LFInst_14_LFInst_0_n6 ) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_3_U9  ( .A1(
        SubCellInst2_LFInst_15_LFInst_3_n16 ), .A2(
        SubCellInst2_LFInst_15_LFInst_3_n15 ), .ZN(MCInst2_MC0_v0_3 [0]) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_3_U8  ( .A1(SubCellInput[61]), .A2(
        SubCellInst2_LFInst_15_LFInst_3_n14 ), .ZN(
        SubCellInst2_LFInst_15_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst2_LFInst_15_LFInst_3_U7  ( .A(SubCellInput[63]), .B(
        SubCellInput[62]), .Z(SubCellInst2_LFInst_15_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_3_U6  ( .A1(
        SubCellInst2_LFInst_15_LFInst_3_n13 ), .A2(
        SubCellInst2_LFInst_15_LFInst_3_n12 ), .ZN(
        SubCellInst2_LFInst_15_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_3_U5  ( .A1(SubCellInput[60]), .A2(
        SubCellInput[62]), .ZN(SubCellInst2_LFInst_15_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst2_LFInst_15_LFInst_3_U4  ( .A(SubCellInput[60]), .B(
        SubCellInst2_LFInst_15_LFInst_3_n11 ), .ZN(
        SubCellInst2_LFInst_15_LFInst_3_n13 ) );
  OR2_X1 SubCellInst2_LFInst_15_LFInst_3_U3  ( .A1(SubCellInput[63]), .A2(
        SubCellInput[61]), .ZN(SubCellInst2_LFInst_15_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_2_U11  ( .A1(
        SubCellInst2_LFInst_15_LFInst_2_n22 ), .A2(
        SubCellInst2_LFInst_15_LFInst_2_n21 ), .ZN(MCInst2_MC0_v0_3 [3]) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_2_U10  ( .A1(SubCellInput[62]), .A2(
        SubCellInst2_LFInst_15_LFInst_2_n20 ), .ZN(
        SubCellInst2_LFInst_15_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst2_LFInst_15_LFInst_2_U9  ( .A1(SubCellInput[61]), .A2(
        SubCellInst2_LFInst_15_LFInst_2_n19 ), .ZN(
        SubCellInst2_LFInst_15_LFInst_2_n20 ) );
  INV_X1 SubCellInst2_LFInst_15_LFInst_2_U8  ( .A(SubCellInput[63]), .ZN(
        SubCellInst2_LFInst_15_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_2_U7  ( .A1(
        SubCellInst2_LFInst_15_LFInst_2_n18 ), .A2(
        SubCellInst2_LFInst_15_LFInst_2_n17 ), .ZN(
        SubCellInst2_LFInst_15_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst2_LFInst_15_LFInst_2_U6  ( .A(
        SubCellInst2_LFInst_15_LFInst_2_n16 ), .B(SubCellInput[62]), .Z(
        SubCellInst2_LFInst_15_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_2_U5  ( .A1(SubCellInput[60]), .A2(
        SubCellInput[61]), .ZN(SubCellInst2_LFInst_15_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_2_U4  ( .A1(
        SubCellInst2_LFInst_15_LFInst_2_n15 ), .A2(SubCellInput[63]), .ZN(
        SubCellInst2_LFInst_15_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst2_LFInst_15_LFInst_2_U3  ( .A(SubCellInput[60]), .B(
        SubCellInput[61]), .ZN(SubCellInst2_LFInst_15_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_1_U12  ( .A1(
        SubCellInst2_LFInst_15_LFInst_1_n18 ), .A2(
        SubCellInst2_LFInst_15_LFInst_1_n17 ), .ZN(MCInst2_MC0_v0_0 [3]) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_1_U11  ( .A1(SubCellInput[61]), .A2(
        SubCellInst2_LFInst_15_LFInst_1_n16 ), .ZN(
        SubCellInst2_LFInst_15_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst2_LFInst_15_LFInst_1_U10  ( .A1(SubCellInput[63]), .A2(
        SubCellInst2_LFInst_15_LFInst_1_n15 ), .ZN(
        SubCellInst2_LFInst_15_LFInst_1_n16 ) );
  AND2_X1 SubCellInst2_LFInst_15_LFInst_1_U9  ( .A1(SubCellInput[60]), .A2(
        SubCellInput[62]), .ZN(SubCellInst2_LFInst_15_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_1_U8  ( .A1(SubCellInput[63]), .A2(
        SubCellInst2_LFInst_15_LFInst_1_n14 ), .ZN(
        SubCellInst2_LFInst_15_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_1_U7  ( .A1(
        SubCellInst2_LFInst_15_LFInst_1_n13 ), .A2(
        SubCellInst2_LFInst_15_LFInst_1_n12 ), .ZN(
        SubCellInst2_LFInst_15_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_1_U6  ( .A1(SubCellInput[60]), .A2(
        SubCellInput[62]), .ZN(SubCellInst2_LFInst_15_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_1_U5  ( .A1(
        SubCellInst2_LFInst_15_LFInst_1_n11 ), .A2(
        SubCellInst2_LFInst_15_LFInst_1_n10 ), .ZN(
        SubCellInst2_LFInst_15_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_1_U4  ( .A1(SubCellInput[60]), .A2(
        SubCellInput[61]), .ZN(SubCellInst2_LFInst_15_LFInst_1_n10 ) );
  INV_X1 SubCellInst2_LFInst_15_LFInst_1_U3  ( .A(SubCellInput[62]), .ZN(
        SubCellInst2_LFInst_15_LFInst_1_n11 ) );
  XNOR2_X1 SubCellInst2_LFInst_15_LFInst_0_U6  ( .A(
        SubCellInst2_LFInst_15_LFInst_0_n6 ), .B(
        SubCellInst2_LFInst_15_LFInst_0_n5 ), .ZN(ShiftRowsOutput2[60]) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_0_U5  ( .A1(SubCellInput[62]), .A2(
        SubCellInst2_LFInst_15_LFInst_0_n4 ), .ZN(
        SubCellInst2_LFInst_15_LFInst_0_n5 ) );
  INV_X1 SubCellInst2_LFInst_15_LFInst_0_U4  ( .A(SubCellInput[61]), .ZN(
        SubCellInst2_LFInst_15_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst2_LFInst_15_LFInst_0_U3  ( .A(SubCellInput[60]), .B(
        SubCellInput[63]), .Z(SubCellInst2_LFInst_15_LFInst_0_n6 ) );
  XNOR2_X1 MCInst2_MC0_v0_2Inst_0_U4  ( .A(MCInst2_MC0_v0_2Inst_0_n2 ), .B(
        MCInst2_MC0_v0_0 [3]), .ZN(MCInst2_MC0_v0_2 [0]) );
  XNOR2_X1 MCInst2_MC0_v0_2Inst_0_U3  ( .A(MCInst2_MC0_v0_3 [0]), .B(
        ShiftRowsOutput2[60]), .ZN(MCInst2_MC0_v0_2Inst_0_n2 ) );
  XOR2_X1 MCInst2_MC0_v1_1Inst_0_U3  ( .A(MCInst2_MC0_v1_3 [3]), .B(
        MCInst2_MC0_v1_3 [0]), .Z(MCInst2_MC0_v1_1 [0]) );
  XNOR2_X1 MCInst2_MC0_v1_2Inst_0_U4  ( .A(MCInst2_MC0_v1_2Inst_0_n2 ), .B(
        MCInst2_MC0_v1_3 [3]), .ZN(MCInst2_MC0_v1_2 [0]) );
  XNOR2_X1 MCInst2_MC0_v1_2Inst_0_U3  ( .A(MCInst2_MC0_v1_3 [0]), .B(
        MCInst2_MC0_v1_3 [2]), .ZN(MCInst2_MC0_v1_2Inst_0_n2 ) );
  XOR2_X1 MCInst2_MC0_v2_1Inst_0_U3  ( .A(MCInst2_MC0_v2_3 [1]), .B(
        MCInst2_MC0_v2_0 [3]), .Z(MCInst2_MC0_v2_1 [0]) );
  XOR2_X1 MCInst2_MC0_v2_2Inst_0_U3  ( .A(MCInst2_MC0_v2_0 [2]), .B(
        MCInst2_MC0_v2_0 [0]), .Z(MCInst2_MC0_v2_2 [0]) );
  XNOR2_X1 MCInst2_MC0_v2_3Inst_0_U5  ( .A(MCInst2_MC0_v2_3Inst_0_n4 ), .B(
        MCInst2_MC0_v2_3Inst_0_n3 ), .ZN(MCInst2_MC0_v2_3 [0]) );
  XNOR2_X1 MCInst2_MC0_v2_3Inst_0_U4  ( .A(MCInst2_MC0_v2_0 [2]), .B(
        MCInst2_MC0_v2_3 [1]), .ZN(MCInst2_MC0_v2_3Inst_0_n3 ) );
  XOR2_X1 MCInst2_MC0_v2_3Inst_0_U3  ( .A(MCInst2_MC0_v2_0 [3]), .B(
        MCInst2_MC0_v2_0 [0]), .Z(MCInst2_MC0_v2_3Inst_0_n4 ) );
  XOR2_X1 MCInst2_MC0_v3_1Inst_0_U3  ( .A(MCInst2_MC0_v3_0 [3]), .B(
        MCInst2_MC0_v3_2 [2]), .Z(MCInst2_MC0_v3_1 [0]) );
  XOR2_X1 MCInst2_MC0_v3_2Inst_0_U3  ( .A(MCInst2_MC0_v3_2 [3]), .B(
        MCInst2_MC0_v3_0 [2]), .Z(MCInst2_MC0_v3_2 [0]) );
  XNOR2_X1 MCInst2_MC0_v3_3Inst_0_U4  ( .A(MCInst2_MC0_v3_3Inst_0_n2 ), .B(
        MCInst2_MC0_v3_0 [2]), .ZN(MCInst2_MC0_v3_3 [0]) );
  XNOR2_X1 MCInst2_MC0_v3_3Inst_0_U3  ( .A(MCInst2_MC0_v3_2 [2]), .B(
        MCInst2_MC0_v3_2 [3]), .ZN(MCInst2_MC0_v3_3Inst_0_n2 ) );
  XOR2_X1 MCInst2_MC0_v0_0Inst_1_U3  ( .A(MCInst2_MC0_v0_3 [3]), .B(
        MCInst2_MC0_v0_3 [0]), .Z(MCInst2_MC0_v0_0 [1]) );
  XOR2_X1 MCInst2_MC0_v0_1Inst_1_U3  ( .A(MCInst2_MC0_v0_0 [3]), .B(
        MCInst2_MC0_v0_3 [3]), .Z(MCInst2_MC0_v0_1 [1]) );
  XNOR2_X1 MCInst2_MC0_v0_2Inst_1_U4  ( .A(MCInst2_MC0_v0_2Inst_1_n2 ), .B(
        MCInst2_MC0_v0_3 [3]), .ZN(MCInst2_MC0_v0_2 [1]) );
  XNOR2_X1 MCInst2_MC0_v0_2Inst_1_U3  ( .A(MCInst2_MC0_v0_3 [0]), .B(
        ShiftRowsOutput2[60]), .ZN(MCInst2_MC0_v0_2Inst_1_n2 ) );
  XOR2_X1 MCInst2_MC0_v0_3Inst_1_U3  ( .A(ShiftRowsOutput2[60]), .B(
        MCInst2_MC0_v0_3 [0]), .Z(MCInst2_MC0_v0_3 [1]) );
  XOR2_X1 MCInst2_MC0_v1_1Inst_1_U3  ( .A(ShiftRowsOutput2[44]), .B(
        MCInst2_MC0_v1_3 [3]), .Z(MCInst2_MC0_v1_1 [1]) );
  XOR2_X1 MCInst2_MC0_v1_2Inst_1_U3  ( .A(ShiftRowsOutput2[44]), .B(
        MCInst2_MC0_v1_3 [2]), .Z(MCInst2_MC0_v1_2 [1]) );
  XOR2_X1 MCInst2_MC0_v1_3Inst_1_U3  ( .A(ShiftRowsOutput2[44]), .B(
        MCInst2_MC0_v1_3 [0]), .Z(MCInst2_MC0_v1_3 [1]) );
  XOR2_X1 MCInst2_MC0_v2_0Inst_1_U3  ( .A(MCInst2_MC0_v2_3 [1]), .B(
        MCInst2_MC0_v2_0 [0]), .Z(MCInst2_MC0_v2_0 [1]) );
  XNOR2_X1 MCInst2_MC0_v2_1Inst_1_U4  ( .A(MCInst2_MC0_v2_1Inst_1_n2 ), .B(
        MCInst2_MC0_v2_0 [3]), .ZN(MCInst2_MC0_v2_1 [1]) );
  XNOR2_X1 MCInst2_MC0_v2_1Inst_1_U3  ( .A(MCInst2_MC0_v2_0 [0]), .B(
        MCInst2_MC0_v2_0 [2]), .ZN(MCInst2_MC0_v2_1Inst_1_n2 ) );
  XNOR2_X1 MCInst2_MC0_v2_2Inst_1_U5  ( .A(MCInst2_MC0_v2_2Inst_1_n4 ), .B(
        MCInst2_MC0_v2_2Inst_1_n3 ), .ZN(MCInst2_MC0_v2_2 [1]) );
  XNOR2_X1 MCInst2_MC0_v2_2Inst_1_U4  ( .A(MCInst2_MC0_v2_0 [2]), .B(
        MCInst2_MC0_v2_3 [1]), .ZN(MCInst2_MC0_v2_2Inst_1_n3 ) );
  XOR2_X1 MCInst2_MC0_v2_2Inst_1_U3  ( .A(MCInst2_MC0_v2_0 [3]), .B(
        MCInst2_MC0_v2_0 [0]), .Z(MCInst2_MC0_v2_2Inst_1_n4 ) );
  XOR2_X1 MCInst2_MC0_v3_0Inst_1_U3  ( .A(MCInst2_MC0_v3_2 [3]), .B(
        MCInst2_MC0_v3_2 [2]), .Z(MCInst2_MC0_v3_0 [1]) );
  XOR2_X1 MCInst2_MC0_v3_1Inst_1_U3  ( .A(MCInst2_MC0_v3_2 [3]), .B(
        MCInst2_MC0_v3_0 [3]), .Z(MCInst2_MC0_v3_1 [1]) );
  XNOR2_X1 MCInst2_MC0_v3_3Inst_1_U4  ( .A(MCInst2_MC0_v3_3Inst_1_n2 ), .B(
        MCInst2_MC0_v3_0 [3]), .ZN(MCInst2_MC0_v3_3 [1]) );
  XNOR2_X1 MCInst2_MC0_v3_3Inst_1_U3  ( .A(MCInst2_MC0_v3_2 [2]), .B(
        MCInst2_MC0_v3_2 [3]), .ZN(MCInst2_MC0_v3_3Inst_1_n2 ) );
  XOR2_X1 MCInst2_MC0_v0_0Inst_2_U3  ( .A(ShiftRowsOutput2[60]), .B(
        MCInst2_MC0_v0_3 [0]), .Z(MCInst2_MC0_v0_0 [2]) );
  XOR2_X1 MCInst2_MC0_v0_1Inst_2_U3  ( .A(MCInst2_MC0_v0_3 [3]), .B(
        MCInst2_MC0_v0_3 [0]), .Z(MCInst2_MC0_v0_1 [2]) );
  XOR2_X1 MCInst2_MC0_v0_2Inst_2_U3  ( .A(MCInst2_MC0_v0_0 [3]), .B(
        MCInst2_MC0_v0_3 [0]), .Z(MCInst2_MC0_v0_2 [2]) );
  XNOR2_X1 MCInst2_MC0_v1_1Inst_2_U4  ( .A(MCInst2_MC0_v1_1Inst_2_n2 ), .B(
        MCInst2_MC0_v1_3 [2]), .ZN(MCInst2_MC0_v1_1 [2]) );
  XNOR2_X1 MCInst2_MC0_v1_1Inst_2_U3  ( .A(MCInst2_MC0_v1_3 [0]), .B(
        ShiftRowsOutput2[44]), .ZN(MCInst2_MC0_v1_1Inst_2_n2 ) );
  XNOR2_X1 MCInst2_MC0_v1_2Inst_2_U4  ( .A(MCInst2_MC0_v1_2Inst_2_n2 ), .B(
        MCInst2_MC0_v1_3 [2]), .ZN(MCInst2_MC0_v1_2 [2]) );
  XNOR2_X1 MCInst2_MC0_v1_2Inst_2_U3  ( .A(MCInst2_MC0_v1_3 [3]), .B(
        ShiftRowsOutput2[44]), .ZN(MCInst2_MC0_v1_2Inst_2_n2 ) );
  XNOR2_X1 MCInst2_MC0_v2_1Inst_2_U4  ( .A(MCInst2_MC0_v2_1Inst_2_n2 ), .B(
        MCInst2_MC0_v2_0 [3]), .ZN(MCInst2_MC0_v2_1 [2]) );
  XNOR2_X1 MCInst2_MC0_v2_1Inst_2_U3  ( .A(MCInst2_MC0_v2_0 [0]), .B(
        MCInst2_MC0_v2_3 [1]), .ZN(MCInst2_MC0_v2_1Inst_2_n2 ) );
  XNOR2_X1 MCInst2_MC0_v2_2Inst_2_U4  ( .A(MCInst2_MC0_v2_2Inst_2_n2 ), .B(
        MCInst2_MC0_v2_0 [3]), .ZN(MCInst2_MC0_v2_2 [2]) );
  XNOR2_X1 MCInst2_MC0_v2_2Inst_2_U3  ( .A(MCInst2_MC0_v2_0 [0]), .B(
        MCInst2_MC0_v2_0 [2]), .ZN(MCInst2_MC0_v2_2Inst_2_n2 ) );
  XOR2_X1 MCInst2_MC0_v2_3Inst_2_U3  ( .A(MCInst2_MC0_v2_3 [1]), .B(
        MCInst2_MC0_v2_0 [2]), .Z(MCInst2_MC0_v2_3 [2]) );
  XNOR2_X1 MCInst2_MC0_v3_1Inst_2_U4  ( .A(MCInst2_MC0_v3_1Inst_2_n2 ), .B(
        MCInst2_MC0_v3_0 [2]), .ZN(MCInst2_MC0_v3_1 [2]) );
  XNOR2_X1 MCInst2_MC0_v3_1Inst_2_U3  ( .A(MCInst2_MC0_v3_2 [2]), .B(
        MCInst2_MC0_v3_2 [3]), .ZN(MCInst2_MC0_v3_1Inst_2_n2 ) );
  XOR2_X1 MCInst2_MC0_v3_3Inst_2_U3  ( .A(MCInst2_MC0_v3_0 [2]), .B(
        MCInst2_MC0_v3_2 [2]), .Z(MCInst2_MC0_v3_3 [2]) );
  XOR2_X1 MCInst2_MC0_v0_1Inst_3_U3  ( .A(ShiftRowsOutput2[60]), .B(
        MCInst2_MC0_v0_3 [0]), .Z(MCInst2_MC0_v0_1 [3]) );
  XOR2_X1 MCInst2_MC0_v0_2Inst_3_U3  ( .A(ShiftRowsOutput2[60]), .B(
        MCInst2_MC0_v0_3 [3]), .Z(MCInst2_MC0_v0_2 [3]) );
  XOR2_X1 MCInst2_MC0_v1_1Inst_3_U3  ( .A(MCInst2_MC0_v1_3 [2]), .B(
        MCInst2_MC0_v1_3 [3]), .Z(MCInst2_MC0_v1_1 [3]) );
  XNOR2_X1 MCInst2_MC0_v1_2Inst_3_U5  ( .A(MCInst2_MC0_v1_2Inst_3_n4 ), .B(
        MCInst2_MC0_v1_2Inst_3_n3 ), .ZN(MCInst2_MC0_v1_2 [3]) );
  XNOR2_X1 MCInst2_MC0_v1_2Inst_3_U4  ( .A(MCInst2_MC0_v1_3 [2]), .B(
        ShiftRowsOutput2[44]), .ZN(MCInst2_MC0_v1_2Inst_3_n3 ) );
  XOR2_X1 MCInst2_MC0_v1_2Inst_3_U3  ( .A(MCInst2_MC0_v1_3 [3]), .B(
        MCInst2_MC0_v1_3 [0]), .Z(MCInst2_MC0_v1_2Inst_3_n4 ) );
  XOR2_X1 MCInst2_MC0_v2_1Inst_3_U3  ( .A(MCInst2_MC0_v2_0 [2]), .B(
        MCInst2_MC0_v2_0 [0]), .Z(MCInst2_MC0_v2_1 [3]) );
  XNOR2_X1 MCInst2_MC0_v2_2Inst_3_U4  ( .A(MCInst2_MC0_v2_2Inst_3_n2 ), .B(
        MCInst2_MC0_v2_0 [3]), .ZN(MCInst2_MC0_v2_2 [3]) );
  XNOR2_X1 MCInst2_MC0_v2_2Inst_3_U3  ( .A(MCInst2_MC0_v2_0 [0]), .B(
        MCInst2_MC0_v2_3 [1]), .ZN(MCInst2_MC0_v2_2Inst_3_n2 ) );
  XNOR2_X1 MCInst2_MC0_v2_3Inst_3_U4  ( .A(MCInst2_MC0_v2_3Inst_3_n2 ), .B(
        MCInst2_MC0_v2_0 [2]), .ZN(MCInst2_MC0_v2_3 [3]) );
  XNOR2_X1 MCInst2_MC0_v2_3Inst_3_U3  ( .A(MCInst2_MC0_v2_0 [3]), .B(
        MCInst2_MC0_v2_3 [1]), .ZN(MCInst2_MC0_v2_3Inst_3_n2 ) );
  XOR2_X1 MCInst2_MC0_v3_1Inst_3_U3  ( .A(MCInst2_MC0_v3_0 [2]), .B(
        MCInst2_MC0_v3_0 [3]), .Z(MCInst2_MC0_v3_1 [3]) );
  XOR2_X1 MCInst2_MC0_v3_3Inst_3_U3  ( .A(MCInst2_MC0_v3_2 [3]), .B(
        MCInst2_MC0_v3_0 [3]), .Z(MCInst2_MC0_v3_3 [3]) );
  XNOR2_X1 MCInst2_MC0_r0Inst_XORInst_0_0_U3  ( .A(
        MCInst2_MC0_r0Inst_XORInst_0_0_n5 ), .B(
        MCInst2_MC0_r0Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[60]) );
  XNOR2_X1 MCInst2_MC0_r0Inst_XORInst_0_0_U2  ( .A(MCInst2_MC0_v3_2 [2]), 
        .B(MCInst2_MC0_v2_0 [0]), .ZN(MCInst2_MC0_r0Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst2_MC0_r0Inst_XORInst_0_0_U1  ( .A(MCInst2_MC0_v0_3 [3]), .B(
        ShiftRowsOutput2[44]), .Z(MCInst2_MC0_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst2_MC0_r0Inst_XORInst_0_1_U3  ( .A(
        MCInst2_MC0_r0Inst_XORInst_0_1_n5 ), .B(
        MCInst2_MC0_r0Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[61]) );
  XNOR2_X1 MCInst2_MC0_r0Inst_XORInst_0_1_U2  ( .A(MCInst2_MC0_v3_0 [1]), 
        .B(MCInst2_MC0_v2_0 [1]), .ZN(MCInst2_MC0_r0Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst2_MC0_r0Inst_XORInst_0_1_U1  ( .A(MCInst2_MC0_v0_0 [1]), .B(
        MCInst2_MC0_v1_3 [2]), .Z(MCInst2_MC0_r0Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst2_MC0_r0Inst_XORInst_0_2_U3  ( .A(
        MCInst2_MC0_r0Inst_XORInst_0_2_n5 ), .B(
        MCInst2_MC0_r0Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[62]) );
  XNOR2_X1 MCInst2_MC0_r0Inst_XORInst_0_2_U2  ( .A(MCInst2_MC0_v3_0 [2]), 
        .B(MCInst2_MC0_v2_0 [2]), .ZN(MCInst2_MC0_r0Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst2_MC0_r0Inst_XORInst_0_2_U1  ( .A(MCInst2_MC0_v0_0 [2]), .B(
        MCInst2_MC0_v1_3 [3]), .Z(MCInst2_MC0_r0Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst2_MC0_r0Inst_XORInst_0_3_U3  ( .A(
        MCInst2_MC0_r0Inst_XORInst_0_3_n5 ), .B(
        MCInst2_MC0_r0Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[63]) );
  XNOR2_X1 MCInst2_MC0_r0Inst_XORInst_0_3_U2  ( .A(MCInst2_MC0_v3_0 [3]), 
        .B(MCInst2_MC0_v2_0 [3]), .ZN(MCInst2_MC0_r0Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst2_MC0_r0Inst_XORInst_0_3_U1  ( .A(MCInst2_MC0_v0_0 [3]), .B(
        MCInst2_MC0_v1_3 [0]), .Z(MCInst2_MC0_r0Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst2_MC0_r1Inst_XORInst_0_0_U3  ( .A(
        MCInst2_MC0_r1Inst_XORInst_0_0_n5 ), .B(
        MCInst2_MC0_r1Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[44]) );
  XNOR2_X1 MCInst2_MC0_r1Inst_XORInst_0_0_U2  ( .A(MCInst2_MC0_v3_1 [0]), 
        .B(MCInst2_MC0_v2_1 [0]), .ZN(MCInst2_MC0_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst2_MC0_r1Inst_XORInst_0_0_U1  ( .A(MCInst2_MC0_v0_0 [3]), .B(
        MCInst2_MC0_v1_1 [0]), .Z(MCInst2_MC0_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst2_MC0_r1Inst_XORInst_0_1_U3  ( .A(
        MCInst2_MC0_r1Inst_XORInst_0_1_n5 ), .B(
        MCInst2_MC0_r1Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[45]) );
  XNOR2_X1 MCInst2_MC0_r1Inst_XORInst_0_1_U2  ( .A(MCInst2_MC0_v3_1 [1]), 
        .B(MCInst2_MC0_v2_1 [1]), .ZN(MCInst2_MC0_r1Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst2_MC0_r1Inst_XORInst_0_1_U1  ( .A(MCInst2_MC0_v0_1 [1]), .B(
        MCInst2_MC0_v1_1 [1]), .Z(MCInst2_MC0_r1Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst2_MC0_r1Inst_XORInst_0_2_U3  ( .A(
        MCInst2_MC0_r1Inst_XORInst_0_2_n5 ), .B(
        MCInst2_MC0_r1Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[46]) );
  XNOR2_X1 MCInst2_MC0_r1Inst_XORInst_0_2_U2  ( .A(MCInst2_MC0_v3_1 [2]), 
        .B(MCInst2_MC0_v2_1 [2]), .ZN(MCInst2_MC0_r1Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst2_MC0_r1Inst_XORInst_0_2_U1  ( .A(MCInst2_MC0_v0_1 [2]), .B(
        MCInst2_MC0_v1_1 [2]), .Z(MCInst2_MC0_r1Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst2_MC0_r1Inst_XORInst_0_3_U3  ( .A(
        MCInst2_MC0_r1Inst_XORInst_0_3_n5 ), .B(
        MCInst2_MC0_r1Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[47]) );
  XNOR2_X1 MCInst2_MC0_r1Inst_XORInst_0_3_U2  ( .A(MCInst2_MC0_v3_1 [3]), 
        .B(MCInst2_MC0_v2_1 [3]), .ZN(MCInst2_MC0_r1Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst2_MC0_r1Inst_XORInst_0_3_U1  ( .A(MCInst2_MC0_v0_1 [3]), .B(
        MCInst2_MC0_v1_1 [3]), .Z(MCInst2_MC0_r1Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst2_MC0_r2Inst_XORInst_0_0_U3  ( .A(
        MCInst2_MC0_r2Inst_XORInst_0_0_n5 ), .B(
        MCInst2_MC0_r2Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[28]) );
  XNOR2_X1 MCInst2_MC0_r2Inst_XORInst_0_0_U2  ( .A(MCInst2_MC0_v3_2 [0]), 
        .B(MCInst2_MC0_v2_2 [0]), .ZN(MCInst2_MC0_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst2_MC0_r2Inst_XORInst_0_0_U1  ( .A(MCInst2_MC0_v0_2 [0]), .B(
        MCInst2_MC0_v1_2 [0]), .Z(MCInst2_MC0_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst2_MC0_r2Inst_XORInst_0_1_U3  ( .A(
        MCInst2_MC0_r2Inst_XORInst_0_1_n5 ), .B(
        MCInst2_MC0_r2Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[29]) );
  XNOR2_X1 MCInst2_MC0_r2Inst_XORInst_0_1_U2  ( .A(MCInst2_MC0_v3_0 [3]), 
        .B(MCInst2_MC0_v2_2 [1]), .ZN(MCInst2_MC0_r2Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst2_MC0_r2Inst_XORInst_0_1_U1  ( .A(MCInst2_MC0_v0_2 [1]), .B(
        MCInst2_MC0_v1_2 [1]), .Z(MCInst2_MC0_r2Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst2_MC0_r2Inst_XORInst_0_2_U3  ( .A(
        MCInst2_MC0_r2Inst_XORInst_0_2_n5 ), .B(
        MCInst2_MC0_r2Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[30]) );
  XNOR2_X1 MCInst2_MC0_r2Inst_XORInst_0_2_U2  ( .A(MCInst2_MC0_v3_2 [2]), 
        .B(MCInst2_MC0_v2_2 [2]), .ZN(MCInst2_MC0_r2Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst2_MC0_r2Inst_XORInst_0_2_U1  ( .A(MCInst2_MC0_v0_2 [2]), .B(
        MCInst2_MC0_v1_2 [2]), .Z(MCInst2_MC0_r2Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst2_MC0_r2Inst_XORInst_0_3_U3  ( .A(
        MCInst2_MC0_r2Inst_XORInst_0_3_n5 ), .B(
        MCInst2_MC0_r2Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[31]) );
  XNOR2_X1 MCInst2_MC0_r2Inst_XORInst_0_3_U2  ( .A(MCInst2_MC0_v3_2 [3]), 
        .B(MCInst2_MC0_v2_2 [3]), .ZN(MCInst2_MC0_r2Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst2_MC0_r2Inst_XORInst_0_3_U1  ( .A(MCInst2_MC0_v0_2 [3]), .B(
        MCInst2_MC0_v1_2 [3]), .Z(MCInst2_MC0_r2Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst2_MC0_r3Inst_XORInst_0_0_U3  ( .A(
        MCInst2_MC0_r3Inst_XORInst_0_0_n5 ), .B(
        MCInst2_MC0_r3Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[12]) );
  XNOR2_X1 MCInst2_MC0_r3Inst_XORInst_0_0_U2  ( .A(MCInst2_MC0_v3_3 [0]), 
        .B(MCInst2_MC0_v2_3 [0]), .ZN(MCInst2_MC0_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst2_MC0_r3Inst_XORInst_0_0_U1  ( .A(MCInst2_MC0_v0_3 [0]), .B(
        MCInst2_MC0_v1_3 [0]), .Z(MCInst2_MC0_r3Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst2_MC0_r3Inst_XORInst_0_1_U3  ( .A(
        MCInst2_MC0_r3Inst_XORInst_0_1_n5 ), .B(
        MCInst2_MC0_r3Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[13]) );
  XNOR2_X1 MCInst2_MC0_r3Inst_XORInst_0_1_U2  ( .A(MCInst2_MC0_v3_3 [1]), 
        .B(MCInst2_MC0_v2_3 [1]), .ZN(MCInst2_MC0_r3Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst2_MC0_r3Inst_XORInst_0_1_U1  ( .A(MCInst2_MC0_v0_3 [1]), .B(
        MCInst2_MC0_v1_3 [1]), .Z(MCInst2_MC0_r3Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst2_MC0_r3Inst_XORInst_0_2_U3  ( .A(
        MCInst2_MC0_r3Inst_XORInst_0_2_n5 ), .B(
        MCInst2_MC0_r3Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[14]) );
  XNOR2_X1 MCInst2_MC0_r3Inst_XORInst_0_2_U2  ( .A(MCInst2_MC0_v3_3 [2]), 
        .B(MCInst2_MC0_v2_3 [2]), .ZN(MCInst2_MC0_r3Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst2_MC0_r3Inst_XORInst_0_2_U1  ( .A(MCInst2_MC0_v0_0 [3]), .B(
        MCInst2_MC0_v1_3 [2]), .Z(MCInst2_MC0_r3Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst2_MC0_r3Inst_XORInst_0_3_U3  ( .A(
        MCInst2_MC0_r3Inst_XORInst_0_3_n5 ), .B(
        MCInst2_MC0_r3Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[15]) );
  XNOR2_X1 MCInst2_MC0_r3Inst_XORInst_0_3_U2  ( .A(MCInst2_MC0_v3_3 [3]), 
        .B(MCInst2_MC0_v2_3 [3]), .ZN(MCInst2_MC0_r3Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst2_MC0_r3Inst_XORInst_0_3_U1  ( .A(MCInst2_MC0_v0_3 [3]), .B(
        MCInst2_MC0_v1_3 [3]), .Z(MCInst2_MC0_r3Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst2_MC1_v0_2Inst_0_U4  ( .A(MCInst2_MC1_v0_2Inst_0_n2 ), .B(
        MCInst2_MC1_v0_0 [3]), .ZN(MCInst2_MC1_v0_2 [0]) );
  XNOR2_X1 MCInst2_MC1_v0_2Inst_0_U3  ( .A(MCInst2_MC1_v0_3 [0]), .B(
        ShiftRowsOutput2[56]), .ZN(MCInst2_MC1_v0_2Inst_0_n2 ) );
  XOR2_X1 MCInst2_MC1_v1_1Inst_0_U3  ( .A(MCInst2_MC1_v1_3 [3]), .B(
        MCInst2_MC1_v1_3 [0]), .Z(MCInst2_MC1_v1_1 [0]) );
  XNOR2_X1 MCInst2_MC1_v1_2Inst_0_U4  ( .A(MCInst2_MC1_v1_2Inst_0_n2 ), .B(
        MCInst2_MC1_v1_3 [3]), .ZN(MCInst2_MC1_v1_2 [0]) );
  XNOR2_X1 MCInst2_MC1_v1_2Inst_0_U3  ( .A(MCInst2_MC1_v1_3 [0]), .B(
        MCInst2_MC1_v1_3 [2]), .ZN(MCInst2_MC1_v1_2Inst_0_n2 ) );
  XOR2_X1 MCInst2_MC1_v2_1Inst_0_U3  ( .A(MCInst2_MC1_v2_3 [1]), .B(
        MCInst2_MC1_v2_0 [3]), .Z(MCInst2_MC1_v2_1 [0]) );
  XOR2_X1 MCInst2_MC1_v2_2Inst_0_U3  ( .A(MCInst2_MC1_v2_0 [2]), .B(
        MCInst2_MC1_v2_0 [0]), .Z(MCInst2_MC1_v2_2 [0]) );
  XNOR2_X1 MCInst2_MC1_v2_3Inst_0_U5  ( .A(MCInst2_MC1_v2_3Inst_0_n4 ), .B(
        MCInst2_MC1_v2_3Inst_0_n3 ), .ZN(MCInst2_MC1_v2_3 [0]) );
  XNOR2_X1 MCInst2_MC1_v2_3Inst_0_U4  ( .A(MCInst2_MC1_v2_0 [2]), .B(
        MCInst2_MC1_v2_3 [1]), .ZN(MCInst2_MC1_v2_3Inst_0_n3 ) );
  XOR2_X1 MCInst2_MC1_v2_3Inst_0_U3  ( .A(MCInst2_MC1_v2_0 [3]), .B(
        MCInst2_MC1_v2_0 [0]), .Z(MCInst2_MC1_v2_3Inst_0_n4 ) );
  XOR2_X1 MCInst2_MC1_v3_1Inst_0_U3  ( .A(MCInst2_MC1_v3_0 [3]), .B(
        MCInst2_MC1_v3_2 [2]), .Z(MCInst2_MC1_v3_1 [0]) );
  XOR2_X1 MCInst2_MC1_v3_2Inst_0_U3  ( .A(MCInst2_MC1_v3_2 [3]), .B(
        MCInst2_MC1_v3_0 [2]), .Z(MCInst2_MC1_v3_2 [0]) );
  XNOR2_X1 MCInst2_MC1_v3_3Inst_0_U4  ( .A(MCInst2_MC1_v3_3Inst_0_n2 ), .B(
        MCInst2_MC1_v3_0 [2]), .ZN(MCInst2_MC1_v3_3 [0]) );
  XNOR2_X1 MCInst2_MC1_v3_3Inst_0_U3  ( .A(MCInst2_MC1_v3_2 [2]), .B(
        MCInst2_MC1_v3_2 [3]), .ZN(MCInst2_MC1_v3_3Inst_0_n2 ) );
  XOR2_X1 MCInst2_MC1_v0_0Inst_1_U3  ( .A(MCInst2_MC1_v0_3 [3]), .B(
        MCInst2_MC1_v0_3 [0]), .Z(MCInst2_MC1_v0_0 [1]) );
  XOR2_X1 MCInst2_MC1_v0_1Inst_1_U3  ( .A(MCInst2_MC1_v0_0 [3]), .B(
        MCInst2_MC1_v0_3 [3]), .Z(MCInst2_MC1_v0_1 [1]) );
  XNOR2_X1 MCInst2_MC1_v0_2Inst_1_U4  ( .A(MCInst2_MC1_v0_2Inst_1_n2 ), .B(
        MCInst2_MC1_v0_3 [3]), .ZN(MCInst2_MC1_v0_2 [1]) );
  XNOR2_X1 MCInst2_MC1_v0_2Inst_1_U3  ( .A(MCInst2_MC1_v0_3 [0]), .B(
        ShiftRowsOutput2[56]), .ZN(MCInst2_MC1_v0_2Inst_1_n2 ) );
  XOR2_X1 MCInst2_MC1_v0_3Inst_1_U3  ( .A(ShiftRowsOutput2[56]), .B(
        MCInst2_MC1_v0_3 [0]), .Z(MCInst2_MC1_v0_3 [1]) );
  XOR2_X1 MCInst2_MC1_v1_1Inst_1_U3  ( .A(ShiftRowsOutput2[40]), .B(
        MCInst2_MC1_v1_3 [3]), .Z(MCInst2_MC1_v1_1 [1]) );
  XOR2_X1 MCInst2_MC1_v1_2Inst_1_U3  ( .A(ShiftRowsOutput2[40]), .B(
        MCInst2_MC1_v1_3 [2]), .Z(MCInst2_MC1_v1_2 [1]) );
  XOR2_X1 MCInst2_MC1_v1_3Inst_1_U3  ( .A(ShiftRowsOutput2[40]), .B(
        MCInst2_MC1_v1_3 [0]), .Z(MCInst2_MC1_v1_3 [1]) );
  XOR2_X1 MCInst2_MC1_v2_0Inst_1_U3  ( .A(MCInst2_MC1_v2_3 [1]), .B(
        MCInst2_MC1_v2_0 [0]), .Z(MCInst2_MC1_v2_0 [1]) );
  XNOR2_X1 MCInst2_MC1_v2_1Inst_1_U4  ( .A(MCInst2_MC1_v2_1Inst_1_n2 ), .B(
        MCInst2_MC1_v2_0 [3]), .ZN(MCInst2_MC1_v2_1 [1]) );
  XNOR2_X1 MCInst2_MC1_v2_1Inst_1_U3  ( .A(MCInst2_MC1_v2_0 [0]), .B(
        MCInst2_MC1_v2_0 [2]), .ZN(MCInst2_MC1_v2_1Inst_1_n2 ) );
  XNOR2_X1 MCInst2_MC1_v2_2Inst_1_U5  ( .A(MCInst2_MC1_v2_2Inst_1_n4 ), .B(
        MCInst2_MC1_v2_2Inst_1_n3 ), .ZN(MCInst2_MC1_v2_2 [1]) );
  XNOR2_X1 MCInst2_MC1_v2_2Inst_1_U4  ( .A(MCInst2_MC1_v2_0 [2]), .B(
        MCInst2_MC1_v2_3 [1]), .ZN(MCInst2_MC1_v2_2Inst_1_n3 ) );
  XOR2_X1 MCInst2_MC1_v2_2Inst_1_U3  ( .A(MCInst2_MC1_v2_0 [3]), .B(
        MCInst2_MC1_v2_0 [0]), .Z(MCInst2_MC1_v2_2Inst_1_n4 ) );
  XOR2_X1 MCInst2_MC1_v3_0Inst_1_U3  ( .A(MCInst2_MC1_v3_2 [3]), .B(
        MCInst2_MC1_v3_2 [2]), .Z(MCInst2_MC1_v3_0 [1]) );
  XOR2_X1 MCInst2_MC1_v3_1Inst_1_U3  ( .A(MCInst2_MC1_v3_2 [3]), .B(
        MCInst2_MC1_v3_0 [3]), .Z(MCInst2_MC1_v3_1 [1]) );
  XNOR2_X1 MCInst2_MC1_v3_3Inst_1_U4  ( .A(MCInst2_MC1_v3_3Inst_1_n2 ), .B(
        MCInst2_MC1_v3_0 [3]), .ZN(MCInst2_MC1_v3_3 [1]) );
  XNOR2_X1 MCInst2_MC1_v3_3Inst_1_U3  ( .A(MCInst2_MC1_v3_2 [2]), .B(
        MCInst2_MC1_v3_2 [3]), .ZN(MCInst2_MC1_v3_3Inst_1_n2 ) );
  XOR2_X1 MCInst2_MC1_v0_0Inst_2_U3  ( .A(ShiftRowsOutput2[56]), .B(
        MCInst2_MC1_v0_3 [0]), .Z(MCInst2_MC1_v0_0 [2]) );
  XOR2_X1 MCInst2_MC1_v0_1Inst_2_U3  ( .A(MCInst2_MC1_v0_3 [3]), .B(
        MCInst2_MC1_v0_3 [0]), .Z(MCInst2_MC1_v0_1 [2]) );
  XOR2_X1 MCInst2_MC1_v0_2Inst_2_U3  ( .A(MCInst2_MC1_v0_0 [3]), .B(
        MCInst2_MC1_v0_3 [0]), .Z(MCInst2_MC1_v0_2 [2]) );
  XNOR2_X1 MCInst2_MC1_v1_1Inst_2_U4  ( .A(MCInst2_MC1_v1_1Inst_2_n2 ), .B(
        MCInst2_MC1_v1_3 [2]), .ZN(MCInst2_MC1_v1_1 [2]) );
  XNOR2_X1 MCInst2_MC1_v1_1Inst_2_U3  ( .A(MCInst2_MC1_v1_3 [0]), .B(
        ShiftRowsOutput2[40]), .ZN(MCInst2_MC1_v1_1Inst_2_n2 ) );
  XNOR2_X1 MCInst2_MC1_v1_2Inst_2_U4  ( .A(MCInst2_MC1_v1_2Inst_2_n2 ), .B(
        MCInst2_MC1_v1_3 [2]), .ZN(MCInst2_MC1_v1_2 [2]) );
  XNOR2_X1 MCInst2_MC1_v1_2Inst_2_U3  ( .A(MCInst2_MC1_v1_3 [3]), .B(
        ShiftRowsOutput2[40]), .ZN(MCInst2_MC1_v1_2Inst_2_n2 ) );
  XNOR2_X1 MCInst2_MC1_v2_1Inst_2_U4  ( .A(MCInst2_MC1_v2_1Inst_2_n2 ), .B(
        MCInst2_MC1_v2_0 [3]), .ZN(MCInst2_MC1_v2_1 [2]) );
  XNOR2_X1 MCInst2_MC1_v2_1Inst_2_U3  ( .A(MCInst2_MC1_v2_0 [0]), .B(
        MCInst2_MC1_v2_3 [1]), .ZN(MCInst2_MC1_v2_1Inst_2_n2 ) );
  XNOR2_X1 MCInst2_MC1_v2_2Inst_2_U4  ( .A(MCInst2_MC1_v2_2Inst_2_n2 ), .B(
        MCInst2_MC1_v2_0 [3]), .ZN(MCInst2_MC1_v2_2 [2]) );
  XNOR2_X1 MCInst2_MC1_v2_2Inst_2_U3  ( .A(MCInst2_MC1_v2_0 [0]), .B(
        MCInst2_MC1_v2_0 [2]), .ZN(MCInst2_MC1_v2_2Inst_2_n2 ) );
  XOR2_X1 MCInst2_MC1_v2_3Inst_2_U3  ( .A(MCInst2_MC1_v2_3 [1]), .B(
        MCInst2_MC1_v2_0 [2]), .Z(MCInst2_MC1_v2_3 [2]) );
  XNOR2_X1 MCInst2_MC1_v3_1Inst_2_U4  ( .A(MCInst2_MC1_v3_1Inst_2_n2 ), .B(
        MCInst2_MC1_v3_0 [2]), .ZN(MCInst2_MC1_v3_1 [2]) );
  XNOR2_X1 MCInst2_MC1_v3_1Inst_2_U3  ( .A(MCInst2_MC1_v3_2 [2]), .B(
        MCInst2_MC1_v3_2 [3]), .ZN(MCInst2_MC1_v3_1Inst_2_n2 ) );
  XOR2_X1 MCInst2_MC1_v3_3Inst_2_U3  ( .A(MCInst2_MC1_v3_0 [2]), .B(
        MCInst2_MC1_v3_2 [2]), .Z(MCInst2_MC1_v3_3 [2]) );
  XOR2_X1 MCInst2_MC1_v0_1Inst_3_U3  ( .A(ShiftRowsOutput2[56]), .B(
        MCInst2_MC1_v0_3 [0]), .Z(MCInst2_MC1_v0_1 [3]) );
  XOR2_X1 MCInst2_MC1_v0_2Inst_3_U3  ( .A(ShiftRowsOutput2[56]), .B(
        MCInst2_MC1_v0_3 [3]), .Z(MCInst2_MC1_v0_2 [3]) );
  XOR2_X1 MCInst2_MC1_v1_1Inst_3_U3  ( .A(MCInst2_MC1_v1_3 [2]), .B(
        MCInst2_MC1_v1_3 [3]), .Z(MCInst2_MC1_v1_1 [3]) );
  XNOR2_X1 MCInst2_MC1_v1_2Inst_3_U5  ( .A(MCInst2_MC1_v1_2Inst_3_n4 ), .B(
        MCInst2_MC1_v1_2Inst_3_n3 ), .ZN(MCInst2_MC1_v1_2 [3]) );
  XNOR2_X1 MCInst2_MC1_v1_2Inst_3_U4  ( .A(MCInst2_MC1_v1_3 [2]), .B(
        ShiftRowsOutput2[40]), .ZN(MCInst2_MC1_v1_2Inst_3_n3 ) );
  XOR2_X1 MCInst2_MC1_v1_2Inst_3_U3  ( .A(MCInst2_MC1_v1_3 [3]), .B(
        MCInst2_MC1_v1_3 [0]), .Z(MCInst2_MC1_v1_2Inst_3_n4 ) );
  XOR2_X1 MCInst2_MC1_v2_1Inst_3_U3  ( .A(MCInst2_MC1_v2_0 [2]), .B(
        MCInst2_MC1_v2_0 [0]), .Z(MCInst2_MC1_v2_1 [3]) );
  XNOR2_X1 MCInst2_MC1_v2_2Inst_3_U4  ( .A(MCInst2_MC1_v2_2Inst_3_n2 ), .B(
        MCInst2_MC1_v2_0 [3]), .ZN(MCInst2_MC1_v2_2 [3]) );
  XNOR2_X1 MCInst2_MC1_v2_2Inst_3_U3  ( .A(MCInst2_MC1_v2_0 [0]), .B(
        MCInst2_MC1_v2_3 [1]), .ZN(MCInst2_MC1_v2_2Inst_3_n2 ) );
  XNOR2_X1 MCInst2_MC1_v2_3Inst_3_U4  ( .A(MCInst2_MC1_v2_3Inst_3_n2 ), .B(
        MCInst2_MC1_v2_0 [2]), .ZN(MCInst2_MC1_v2_3 [3]) );
  XNOR2_X1 MCInst2_MC1_v2_3Inst_3_U3  ( .A(MCInst2_MC1_v2_0 [3]), .B(
        MCInst2_MC1_v2_3 [1]), .ZN(MCInst2_MC1_v2_3Inst_3_n2 ) );
  XOR2_X1 MCInst2_MC1_v3_1Inst_3_U3  ( .A(MCInst2_MC1_v3_0 [2]), .B(
        MCInst2_MC1_v3_0 [3]), .Z(MCInst2_MC1_v3_1 [3]) );
  XOR2_X1 MCInst2_MC1_v3_3Inst_3_U3  ( .A(MCInst2_MC1_v3_2 [3]), .B(
        MCInst2_MC1_v3_0 [3]), .Z(MCInst2_MC1_v3_3 [3]) );
  XNOR2_X1 MCInst2_MC1_r0Inst_XORInst_0_0_U3  ( .A(
        MCInst2_MC1_r0Inst_XORInst_0_0_n5 ), .B(
        MCInst2_MC1_r0Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[56]) );
  XNOR2_X1 MCInst2_MC1_r0Inst_XORInst_0_0_U2  ( .A(MCInst2_MC1_v3_2 [2]), 
        .B(MCInst2_MC1_v2_0 [0]), .ZN(MCInst2_MC1_r0Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst2_MC1_r0Inst_XORInst_0_0_U1  ( .A(MCInst2_MC1_v0_3 [3]), .B(
        ShiftRowsOutput2[40]), .Z(MCInst2_MC1_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst2_MC1_r0Inst_XORInst_0_1_U3  ( .A(
        MCInst2_MC1_r0Inst_XORInst_0_1_n5 ), .B(
        MCInst2_MC1_r0Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[57]) );
  XNOR2_X1 MCInst2_MC1_r0Inst_XORInst_0_1_U2  ( .A(MCInst2_MC1_v3_0 [1]), 
        .B(MCInst2_MC1_v2_0 [1]), .ZN(MCInst2_MC1_r0Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst2_MC1_r0Inst_XORInst_0_1_U1  ( .A(MCInst2_MC1_v0_0 [1]), .B(
        MCInst2_MC1_v1_3 [2]), .Z(MCInst2_MC1_r0Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst2_MC1_r0Inst_XORInst_0_2_U3  ( .A(
        MCInst2_MC1_r0Inst_XORInst_0_2_n5 ), .B(
        MCInst2_MC1_r0Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[58]) );
  XNOR2_X1 MCInst2_MC1_r0Inst_XORInst_0_2_U2  ( .A(MCInst2_MC1_v3_0 [2]), 
        .B(MCInst2_MC1_v2_0 [2]), .ZN(MCInst2_MC1_r0Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst2_MC1_r0Inst_XORInst_0_2_U1  ( .A(MCInst2_MC1_v0_0 [2]), .B(
        MCInst2_MC1_v1_3 [3]), .Z(MCInst2_MC1_r0Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst2_MC1_r0Inst_XORInst_0_3_U3  ( .A(
        MCInst2_MC1_r0Inst_XORInst_0_3_n5 ), .B(
        MCInst2_MC1_r0Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[59]) );
  XNOR2_X1 MCInst2_MC1_r0Inst_XORInst_0_3_U2  ( .A(MCInst2_MC1_v3_0 [3]), 
        .B(MCInst2_MC1_v2_0 [3]), .ZN(MCInst2_MC1_r0Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst2_MC1_r0Inst_XORInst_0_3_U1  ( .A(MCInst2_MC1_v0_0 [3]), .B(
        MCInst2_MC1_v1_3 [0]), .Z(MCInst2_MC1_r0Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst2_MC1_r1Inst_XORInst_0_0_U3  ( .A(
        MCInst2_MC1_r1Inst_XORInst_0_0_n5 ), .B(
        MCInst2_MC1_r1Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[40]) );
  XNOR2_X1 MCInst2_MC1_r1Inst_XORInst_0_0_U2  ( .A(MCInst2_MC1_v3_1 [0]), 
        .B(MCInst2_MC1_v2_1 [0]), .ZN(MCInst2_MC1_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst2_MC1_r1Inst_XORInst_0_0_U1  ( .A(MCInst2_MC1_v0_0 [3]), .B(
        MCInst2_MC1_v1_1 [0]), .Z(MCInst2_MC1_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst2_MC1_r1Inst_XORInst_0_1_U3  ( .A(
        MCInst2_MC1_r1Inst_XORInst_0_1_n5 ), .B(
        MCInst2_MC1_r1Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[41]) );
  XNOR2_X1 MCInst2_MC1_r1Inst_XORInst_0_1_U2  ( .A(MCInst2_MC1_v3_1 [1]), 
        .B(MCInst2_MC1_v2_1 [1]), .ZN(MCInst2_MC1_r1Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst2_MC1_r1Inst_XORInst_0_1_U1  ( .A(MCInst2_MC1_v0_1 [1]), .B(
        MCInst2_MC1_v1_1 [1]), .Z(MCInst2_MC1_r1Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst2_MC1_r1Inst_XORInst_0_2_U3  ( .A(
        MCInst2_MC1_r1Inst_XORInst_0_2_n5 ), .B(
        MCInst2_MC1_r1Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[42]) );
  XNOR2_X1 MCInst2_MC1_r1Inst_XORInst_0_2_U2  ( .A(MCInst2_MC1_v3_1 [2]), 
        .B(MCInst2_MC1_v2_1 [2]), .ZN(MCInst2_MC1_r1Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst2_MC1_r1Inst_XORInst_0_2_U1  ( .A(MCInst2_MC1_v0_1 [2]), .B(
        MCInst2_MC1_v1_1 [2]), .Z(MCInst2_MC1_r1Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst2_MC1_r1Inst_XORInst_0_3_U3  ( .A(
        MCInst2_MC1_r1Inst_XORInst_0_3_n5 ), .B(
        MCInst2_MC1_r1Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[43]) );
  XNOR2_X1 MCInst2_MC1_r1Inst_XORInst_0_3_U2  ( .A(MCInst2_MC1_v3_1 [3]), 
        .B(MCInst2_MC1_v2_1 [3]), .ZN(MCInst2_MC1_r1Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst2_MC1_r1Inst_XORInst_0_3_U1  ( .A(MCInst2_MC1_v0_1 [3]), .B(
        MCInst2_MC1_v1_1 [3]), .Z(MCInst2_MC1_r1Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst2_MC1_r2Inst_XORInst_0_0_U3  ( .A(
        MCInst2_MC1_r2Inst_XORInst_0_0_n5 ), .B(
        MCInst2_MC1_r2Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[24]) );
  XNOR2_X1 MCInst2_MC1_r2Inst_XORInst_0_0_U2  ( .A(MCInst2_MC1_v3_2 [0]), 
        .B(MCInst2_MC1_v2_2 [0]), .ZN(MCInst2_MC1_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst2_MC1_r2Inst_XORInst_0_0_U1  ( .A(MCInst2_MC1_v0_2 [0]), .B(
        MCInst2_MC1_v1_2 [0]), .Z(MCInst2_MC1_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst2_MC1_r2Inst_XORInst_0_1_U3  ( .A(
        MCInst2_MC1_r2Inst_XORInst_0_1_n5 ), .B(
        MCInst2_MC1_r2Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[25]) );
  XNOR2_X1 MCInst2_MC1_r2Inst_XORInst_0_1_U2  ( .A(MCInst2_MC1_v3_0 [3]), 
        .B(MCInst2_MC1_v2_2 [1]), .ZN(MCInst2_MC1_r2Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst2_MC1_r2Inst_XORInst_0_1_U1  ( .A(MCInst2_MC1_v0_2 [1]), .B(
        MCInst2_MC1_v1_2 [1]), .Z(MCInst2_MC1_r2Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst2_MC1_r2Inst_XORInst_0_2_U3  ( .A(
        MCInst2_MC1_r2Inst_XORInst_0_2_n5 ), .B(
        MCInst2_MC1_r2Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[26]) );
  XNOR2_X1 MCInst2_MC1_r2Inst_XORInst_0_2_U2  ( .A(MCInst2_MC1_v3_2 [2]), 
        .B(MCInst2_MC1_v2_2 [2]), .ZN(MCInst2_MC1_r2Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst2_MC1_r2Inst_XORInst_0_2_U1  ( .A(MCInst2_MC1_v0_2 [2]), .B(
        MCInst2_MC1_v1_2 [2]), .Z(MCInst2_MC1_r2Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst2_MC1_r2Inst_XORInst_0_3_U3  ( .A(
        MCInst2_MC1_r2Inst_XORInst_0_3_n5 ), .B(
        MCInst2_MC1_r2Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[27]) );
  XNOR2_X1 MCInst2_MC1_r2Inst_XORInst_0_3_U2  ( .A(MCInst2_MC1_v3_2 [3]), 
        .B(MCInst2_MC1_v2_2 [3]), .ZN(MCInst2_MC1_r2Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst2_MC1_r2Inst_XORInst_0_3_U1  ( .A(MCInst2_MC1_v0_2 [3]), .B(
        MCInst2_MC1_v1_2 [3]), .Z(MCInst2_MC1_r2Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst2_MC1_r3Inst_XORInst_0_0_U3  ( .A(
        MCInst2_MC1_r3Inst_XORInst_0_0_n5 ), .B(
        MCInst2_MC1_r3Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[8]) );
  XNOR2_X1 MCInst2_MC1_r3Inst_XORInst_0_0_U2  ( .A(MCInst2_MC1_v3_3 [0]), 
        .B(MCInst2_MC1_v2_3 [0]), .ZN(MCInst2_MC1_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst2_MC1_r3Inst_XORInst_0_0_U1  ( .A(MCInst2_MC1_v0_3 [0]), .B(
        MCInst2_MC1_v1_3 [0]), .Z(MCInst2_MC1_r3Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst2_MC1_r3Inst_XORInst_0_1_U3  ( .A(
        MCInst2_MC1_r3Inst_XORInst_0_1_n5 ), .B(
        MCInst2_MC1_r3Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[9]) );
  XNOR2_X1 MCInst2_MC1_r3Inst_XORInst_0_1_U2  ( .A(MCInst2_MC1_v3_3 [1]), 
        .B(MCInst2_MC1_v2_3 [1]), .ZN(MCInst2_MC1_r3Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst2_MC1_r3Inst_XORInst_0_1_U1  ( .A(MCInst2_MC1_v0_3 [1]), .B(
        MCInst2_MC1_v1_3 [1]), .Z(MCInst2_MC1_r3Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst2_MC1_r3Inst_XORInst_0_2_U3  ( .A(
        MCInst2_MC1_r3Inst_XORInst_0_2_n5 ), .B(
        MCInst2_MC1_r3Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[10]) );
  XNOR2_X1 MCInst2_MC1_r3Inst_XORInst_0_2_U2  ( .A(MCInst2_MC1_v3_3 [2]), 
        .B(MCInst2_MC1_v2_3 [2]), .ZN(MCInst2_MC1_r3Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst2_MC1_r3Inst_XORInst_0_2_U1  ( .A(MCInst2_MC1_v0_0 [3]), .B(
        MCInst2_MC1_v1_3 [2]), .Z(MCInst2_MC1_r3Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst2_MC1_r3Inst_XORInst_0_3_U3  ( .A(
        MCInst2_MC1_r3Inst_XORInst_0_3_n5 ), .B(
        MCInst2_MC1_r3Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[11]) );
  XNOR2_X1 MCInst2_MC1_r3Inst_XORInst_0_3_U2  ( .A(MCInst2_MC1_v3_3 [3]), 
        .B(MCInst2_MC1_v2_3 [3]), .ZN(MCInst2_MC1_r3Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst2_MC1_r3Inst_XORInst_0_3_U1  ( .A(MCInst2_MC1_v0_3 [3]), .B(
        MCInst2_MC1_v1_3 [3]), .Z(MCInst2_MC1_r3Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst2_MC2_v0_2Inst_0_U4  ( .A(MCInst2_MC2_v0_2Inst_0_n2 ), .B(
        MCInst2_MC2_v0_0 [3]), .ZN(MCInst2_MC2_v0_2 [0]) );
  XNOR2_X1 MCInst2_MC2_v0_2Inst_0_U3  ( .A(MCInst2_MC2_v0_3 [0]), .B(
        ShiftRowsOutput2[52]), .ZN(MCInst2_MC2_v0_2Inst_0_n2 ) );
  XOR2_X1 MCInst2_MC2_v1_1Inst_0_U3  ( .A(MCInst2_MC2_v1_3 [3]), .B(
        MCInst2_MC2_v1_3 [0]), .Z(MCInst2_MC2_v1_1 [0]) );
  XNOR2_X1 MCInst2_MC2_v1_2Inst_0_U4  ( .A(MCInst2_MC2_v1_2Inst_0_n2 ), .B(
        MCInst2_MC2_v1_3 [3]), .ZN(MCInst2_MC2_v1_2 [0]) );
  XNOR2_X1 MCInst2_MC2_v1_2Inst_0_U3  ( .A(MCInst2_MC2_v1_3 [0]), .B(
        MCInst2_MC2_v1_3 [2]), .ZN(MCInst2_MC2_v1_2Inst_0_n2 ) );
  XOR2_X1 MCInst2_MC2_v2_1Inst_0_U3  ( .A(MCInst2_MC2_v2_3 [1]), .B(
        MCInst2_MC2_v2_0 [3]), .Z(MCInst2_MC2_v2_1 [0]) );
  XOR2_X1 MCInst2_MC2_v2_2Inst_0_U3  ( .A(MCInst2_MC2_v2_0 [2]), .B(
        MCInst2_MC2_v2_0 [0]), .Z(MCInst2_MC2_v2_2 [0]) );
  XNOR2_X1 MCInst2_MC2_v2_3Inst_0_U5  ( .A(MCInst2_MC2_v2_3Inst_0_n4 ), .B(
        MCInst2_MC2_v2_3Inst_0_n3 ), .ZN(MCInst2_MC2_v2_3 [0]) );
  XNOR2_X1 MCInst2_MC2_v2_3Inst_0_U4  ( .A(MCInst2_MC2_v2_0 [2]), .B(
        MCInst2_MC2_v2_3 [1]), .ZN(MCInst2_MC2_v2_3Inst_0_n3 ) );
  XOR2_X1 MCInst2_MC2_v2_3Inst_0_U3  ( .A(MCInst2_MC2_v2_0 [3]), .B(
        MCInst2_MC2_v2_0 [0]), .Z(MCInst2_MC2_v2_3Inst_0_n4 ) );
  XOR2_X1 MCInst2_MC2_v3_1Inst_0_U3  ( .A(MCInst2_MC2_v3_0 [3]), .B(
        MCInst2_MC2_v3_2 [2]), .Z(MCInst2_MC2_v3_1 [0]) );
  XOR2_X1 MCInst2_MC2_v3_2Inst_0_U3  ( .A(MCInst2_MC2_v3_2 [3]), .B(
        MCInst2_MC2_v3_0 [2]), .Z(MCInst2_MC2_v3_2 [0]) );
  XNOR2_X1 MCInst2_MC2_v3_3Inst_0_U4  ( .A(MCInst2_MC2_v3_3Inst_0_n2 ), .B(
        MCInst2_MC2_v3_0 [2]), .ZN(MCInst2_MC2_v3_3 [0]) );
  XNOR2_X1 MCInst2_MC2_v3_3Inst_0_U3  ( .A(MCInst2_MC2_v3_2 [2]), .B(
        MCInst2_MC2_v3_2 [3]), .ZN(MCInst2_MC2_v3_3Inst_0_n2 ) );
  XOR2_X1 MCInst2_MC2_v0_0Inst_1_U3  ( .A(MCInst2_MC2_v0_3 [3]), .B(
        MCInst2_MC2_v0_3 [0]), .Z(MCInst2_MC2_v0_0 [1]) );
  XOR2_X1 MCInst2_MC2_v0_1Inst_1_U3  ( .A(MCInst2_MC2_v0_0 [3]), .B(
        MCInst2_MC2_v0_3 [3]), .Z(MCInst2_MC2_v0_1 [1]) );
  XNOR2_X1 MCInst2_MC2_v0_2Inst_1_U4  ( .A(MCInst2_MC2_v0_2Inst_1_n2 ), .B(
        MCInst2_MC2_v0_3 [3]), .ZN(MCInst2_MC2_v0_2 [1]) );
  XNOR2_X1 MCInst2_MC2_v0_2Inst_1_U3  ( .A(MCInst2_MC2_v0_3 [0]), .B(
        ShiftRowsOutput2[52]), .ZN(MCInst2_MC2_v0_2Inst_1_n2 ) );
  XOR2_X1 MCInst2_MC2_v0_3Inst_1_U3  ( .A(ShiftRowsOutput2[52]), .B(
        MCInst2_MC2_v0_3 [0]), .Z(MCInst2_MC2_v0_3 [1]) );
  XOR2_X1 MCInst2_MC2_v1_1Inst_1_U3  ( .A(ShiftRowsOutput2[36]), .B(
        MCInst2_MC2_v1_3 [3]), .Z(MCInst2_MC2_v1_1 [1]) );
  XOR2_X1 MCInst2_MC2_v1_2Inst_1_U3  ( .A(ShiftRowsOutput2[36]), .B(
        MCInst2_MC2_v1_3 [2]), .Z(MCInst2_MC2_v1_2 [1]) );
  XOR2_X1 MCInst2_MC2_v1_3Inst_1_U3  ( .A(ShiftRowsOutput2[36]), .B(
        MCInst2_MC2_v1_3 [0]), .Z(MCInst2_MC2_v1_3 [1]) );
  XOR2_X1 MCInst2_MC2_v2_0Inst_1_U3  ( .A(MCInst2_MC2_v2_3 [1]), .B(
        MCInst2_MC2_v2_0 [0]), .Z(MCInst2_MC2_v2_0 [1]) );
  XNOR2_X1 MCInst2_MC2_v2_1Inst_1_U4  ( .A(MCInst2_MC2_v2_1Inst_1_n2 ), .B(
        MCInst2_MC2_v2_0 [3]), .ZN(MCInst2_MC2_v2_1 [1]) );
  XNOR2_X1 MCInst2_MC2_v2_1Inst_1_U3  ( .A(MCInst2_MC2_v2_0 [0]), .B(
        MCInst2_MC2_v2_0 [2]), .ZN(MCInst2_MC2_v2_1Inst_1_n2 ) );
  XNOR2_X1 MCInst2_MC2_v2_2Inst_1_U5  ( .A(MCInst2_MC2_v2_2Inst_1_n4 ), .B(
        MCInst2_MC2_v2_2Inst_1_n3 ), .ZN(MCInst2_MC2_v2_2 [1]) );
  XNOR2_X1 MCInst2_MC2_v2_2Inst_1_U4  ( .A(MCInst2_MC2_v2_0 [2]), .B(
        MCInst2_MC2_v2_3 [1]), .ZN(MCInst2_MC2_v2_2Inst_1_n3 ) );
  XOR2_X1 MCInst2_MC2_v2_2Inst_1_U3  ( .A(MCInst2_MC2_v2_0 [3]), .B(
        MCInst2_MC2_v2_0 [0]), .Z(MCInst2_MC2_v2_2Inst_1_n4 ) );
  XOR2_X1 MCInst2_MC2_v3_0Inst_1_U3  ( .A(MCInst2_MC2_v3_2 [3]), .B(
        MCInst2_MC2_v3_2 [2]), .Z(MCInst2_MC2_v3_0 [1]) );
  XOR2_X1 MCInst2_MC2_v3_1Inst_1_U3  ( .A(MCInst2_MC2_v3_2 [3]), .B(
        MCInst2_MC2_v3_0 [3]), .Z(MCInst2_MC2_v3_1 [1]) );
  XNOR2_X1 MCInst2_MC2_v3_3Inst_1_U4  ( .A(MCInst2_MC2_v3_3Inst_1_n2 ), .B(
        MCInst2_MC2_v3_0 [3]), .ZN(MCInst2_MC2_v3_3 [1]) );
  XNOR2_X1 MCInst2_MC2_v3_3Inst_1_U3  ( .A(MCInst2_MC2_v3_2 [2]), .B(
        MCInst2_MC2_v3_2 [3]), .ZN(MCInst2_MC2_v3_3Inst_1_n2 ) );
  XOR2_X1 MCInst2_MC2_v0_0Inst_2_U3  ( .A(ShiftRowsOutput2[52]), .B(
        MCInst2_MC2_v0_3 [0]), .Z(MCInst2_MC2_v0_0 [2]) );
  XOR2_X1 MCInst2_MC2_v0_1Inst_2_U3  ( .A(MCInst2_MC2_v0_3 [3]), .B(
        MCInst2_MC2_v0_3 [0]), .Z(MCInst2_MC2_v0_1 [2]) );
  XOR2_X1 MCInst2_MC2_v0_2Inst_2_U3  ( .A(MCInst2_MC2_v0_0 [3]), .B(
        MCInst2_MC2_v0_3 [0]), .Z(MCInst2_MC2_v0_2 [2]) );
  XNOR2_X1 MCInst2_MC2_v1_1Inst_2_U4  ( .A(MCInst2_MC2_v1_1Inst_2_n2 ), .B(
        MCInst2_MC2_v1_3 [2]), .ZN(MCInst2_MC2_v1_1 [2]) );
  XNOR2_X1 MCInst2_MC2_v1_1Inst_2_U3  ( .A(MCInst2_MC2_v1_3 [0]), .B(
        ShiftRowsOutput2[36]), .ZN(MCInst2_MC2_v1_1Inst_2_n2 ) );
  XNOR2_X1 MCInst2_MC2_v1_2Inst_2_U4  ( .A(MCInst2_MC2_v1_2Inst_2_n2 ), .B(
        MCInst2_MC2_v1_3 [2]), .ZN(MCInst2_MC2_v1_2 [2]) );
  XNOR2_X1 MCInst2_MC2_v1_2Inst_2_U3  ( .A(MCInst2_MC2_v1_3 [3]), .B(
        ShiftRowsOutput2[36]), .ZN(MCInst2_MC2_v1_2Inst_2_n2 ) );
  XNOR2_X1 MCInst2_MC2_v2_1Inst_2_U4  ( .A(MCInst2_MC2_v2_1Inst_2_n2 ), .B(
        MCInst2_MC2_v2_0 [3]), .ZN(MCInst2_MC2_v2_1 [2]) );
  XNOR2_X1 MCInst2_MC2_v2_1Inst_2_U3  ( .A(MCInst2_MC2_v2_0 [0]), .B(
        MCInst2_MC2_v2_3 [1]), .ZN(MCInst2_MC2_v2_1Inst_2_n2 ) );
  XNOR2_X1 MCInst2_MC2_v2_2Inst_2_U4  ( .A(MCInst2_MC2_v2_2Inst_2_n2 ), .B(
        MCInst2_MC2_v2_0 [3]), .ZN(MCInst2_MC2_v2_2 [2]) );
  XNOR2_X1 MCInst2_MC2_v2_2Inst_2_U3  ( .A(MCInst2_MC2_v2_0 [0]), .B(
        MCInst2_MC2_v2_0 [2]), .ZN(MCInst2_MC2_v2_2Inst_2_n2 ) );
  XOR2_X1 MCInst2_MC2_v2_3Inst_2_U3  ( .A(MCInst2_MC2_v2_3 [1]), .B(
        MCInst2_MC2_v2_0 [2]), .Z(MCInst2_MC2_v2_3 [2]) );
  XNOR2_X1 MCInst2_MC2_v3_1Inst_2_U4  ( .A(MCInst2_MC2_v3_1Inst_2_n2 ), .B(
        MCInst2_MC2_v3_0 [2]), .ZN(MCInst2_MC2_v3_1 [2]) );
  XNOR2_X1 MCInst2_MC2_v3_1Inst_2_U3  ( .A(MCInst2_MC2_v3_2 [2]), .B(
        MCInst2_MC2_v3_2 [3]), .ZN(MCInst2_MC2_v3_1Inst_2_n2 ) );
  XOR2_X1 MCInst2_MC2_v3_3Inst_2_U3  ( .A(MCInst2_MC2_v3_0 [2]), .B(
        MCInst2_MC2_v3_2 [2]), .Z(MCInst2_MC2_v3_3 [2]) );
  XOR2_X1 MCInst2_MC2_v0_1Inst_3_U3  ( .A(ShiftRowsOutput2[52]), .B(
        MCInst2_MC2_v0_3 [0]), .Z(MCInst2_MC2_v0_1 [3]) );
  XOR2_X1 MCInst2_MC2_v0_2Inst_3_U3  ( .A(ShiftRowsOutput2[52]), .B(
        MCInst2_MC2_v0_3 [3]), .Z(MCInst2_MC2_v0_2 [3]) );
  XOR2_X1 MCInst2_MC2_v1_1Inst_3_U3  ( .A(MCInst2_MC2_v1_3 [2]), .B(
        MCInst2_MC2_v1_3 [3]), .Z(MCInst2_MC2_v1_1 [3]) );
  XNOR2_X1 MCInst2_MC2_v1_2Inst_3_U5  ( .A(MCInst2_MC2_v1_2Inst_3_n4 ), .B(
        MCInst2_MC2_v1_2Inst_3_n3 ), .ZN(MCInst2_MC2_v1_2 [3]) );
  XNOR2_X1 MCInst2_MC2_v1_2Inst_3_U4  ( .A(MCInst2_MC2_v1_3 [2]), .B(
        ShiftRowsOutput2[36]), .ZN(MCInst2_MC2_v1_2Inst_3_n3 ) );
  XOR2_X1 MCInst2_MC2_v1_2Inst_3_U3  ( .A(MCInst2_MC2_v1_3 [3]), .B(
        MCInst2_MC2_v1_3 [0]), .Z(MCInst2_MC2_v1_2Inst_3_n4 ) );
  XOR2_X1 MCInst2_MC2_v2_1Inst_3_U3  ( .A(MCInst2_MC2_v2_0 [2]), .B(
        MCInst2_MC2_v2_0 [0]), .Z(MCInst2_MC2_v2_1 [3]) );
  XNOR2_X1 MCInst2_MC2_v2_2Inst_3_U4  ( .A(MCInst2_MC2_v2_2Inst_3_n2 ), .B(
        MCInst2_MC2_v2_0 [3]), .ZN(MCInst2_MC2_v2_2 [3]) );
  XNOR2_X1 MCInst2_MC2_v2_2Inst_3_U3  ( .A(MCInst2_MC2_v2_0 [0]), .B(
        MCInst2_MC2_v2_3 [1]), .ZN(MCInst2_MC2_v2_2Inst_3_n2 ) );
  XNOR2_X1 MCInst2_MC2_v2_3Inst_3_U4  ( .A(MCInst2_MC2_v2_3Inst_3_n2 ), .B(
        MCInst2_MC2_v2_0 [2]), .ZN(MCInst2_MC2_v2_3 [3]) );
  XNOR2_X1 MCInst2_MC2_v2_3Inst_3_U3  ( .A(MCInst2_MC2_v2_0 [3]), .B(
        MCInst2_MC2_v2_3 [1]), .ZN(MCInst2_MC2_v2_3Inst_3_n2 ) );
  XOR2_X1 MCInst2_MC2_v3_1Inst_3_U3  ( .A(MCInst2_MC2_v3_0 [2]), .B(
        MCInst2_MC2_v3_0 [3]), .Z(MCInst2_MC2_v3_1 [3]) );
  XOR2_X1 MCInst2_MC2_v3_3Inst_3_U3  ( .A(MCInst2_MC2_v3_2 [3]), .B(
        MCInst2_MC2_v3_0 [3]), .Z(MCInst2_MC2_v3_3 [3]) );
  XNOR2_X1 MCInst2_MC2_r0Inst_XORInst_0_0_U3  ( .A(
        MCInst2_MC2_r0Inst_XORInst_0_0_n5 ), .B(
        MCInst2_MC2_r0Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[52]) );
  XNOR2_X1 MCInst2_MC2_r0Inst_XORInst_0_0_U2  ( .A(MCInst2_MC2_v3_2 [2]), 
        .B(MCInst2_MC2_v2_0 [0]), .ZN(MCInst2_MC2_r0Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst2_MC2_r0Inst_XORInst_0_0_U1  ( .A(MCInst2_MC2_v0_3 [3]), .B(
        ShiftRowsOutput2[36]), .Z(MCInst2_MC2_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst2_MC2_r0Inst_XORInst_0_1_U3  ( .A(
        MCInst2_MC2_r0Inst_XORInst_0_1_n5 ), .B(
        MCInst2_MC2_r0Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[53]) );
  XNOR2_X1 MCInst2_MC2_r0Inst_XORInst_0_1_U2  ( .A(MCInst2_MC2_v3_0 [1]), 
        .B(MCInst2_MC2_v2_0 [1]), .ZN(MCInst2_MC2_r0Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst2_MC2_r0Inst_XORInst_0_1_U1  ( .A(MCInst2_MC2_v0_0 [1]), .B(
        MCInst2_MC2_v1_3 [2]), .Z(MCInst2_MC2_r0Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst2_MC2_r0Inst_XORInst_0_2_U3  ( .A(
        MCInst2_MC2_r0Inst_XORInst_0_2_n5 ), .B(
        MCInst2_MC2_r0Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[54]) );
  XNOR2_X1 MCInst2_MC2_r0Inst_XORInst_0_2_U2  ( .A(MCInst2_MC2_v3_0 [2]), 
        .B(MCInst2_MC2_v2_0 [2]), .ZN(MCInst2_MC2_r0Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst2_MC2_r0Inst_XORInst_0_2_U1  ( .A(MCInst2_MC2_v0_0 [2]), .B(
        MCInst2_MC2_v1_3 [3]), .Z(MCInst2_MC2_r0Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst2_MC2_r0Inst_XORInst_0_3_U3  ( .A(
        MCInst2_MC2_r0Inst_XORInst_0_3_n5 ), .B(
        MCInst2_MC2_r0Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[55]) );
  XNOR2_X1 MCInst2_MC2_r0Inst_XORInst_0_3_U2  ( .A(MCInst2_MC2_v3_0 [3]), 
        .B(MCInst2_MC2_v2_0 [3]), .ZN(MCInst2_MC2_r0Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst2_MC2_r0Inst_XORInst_0_3_U1  ( .A(MCInst2_MC2_v0_0 [3]), .B(
        MCInst2_MC2_v1_3 [0]), .Z(MCInst2_MC2_r0Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst2_MC2_r1Inst_XORInst_0_0_U3  ( .A(
        MCInst2_MC2_r1Inst_XORInst_0_0_n5 ), .B(
        MCInst2_MC2_r1Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[36]) );
  XNOR2_X1 MCInst2_MC2_r1Inst_XORInst_0_0_U2  ( .A(MCInst2_MC2_v3_1 [0]), 
        .B(MCInst2_MC2_v2_1 [0]), .ZN(MCInst2_MC2_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst2_MC2_r1Inst_XORInst_0_0_U1  ( .A(MCInst2_MC2_v0_0 [3]), .B(
        MCInst2_MC2_v1_1 [0]), .Z(MCInst2_MC2_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst2_MC2_r1Inst_XORInst_0_1_U3  ( .A(
        MCInst2_MC2_r1Inst_XORInst_0_1_n5 ), .B(
        MCInst2_MC2_r1Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[37]) );
  XNOR2_X1 MCInst2_MC2_r1Inst_XORInst_0_1_U2  ( .A(MCInst2_MC2_v3_1 [1]), 
        .B(MCInst2_MC2_v2_1 [1]), .ZN(MCInst2_MC2_r1Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst2_MC2_r1Inst_XORInst_0_1_U1  ( .A(MCInst2_MC2_v0_1 [1]), .B(
        MCInst2_MC2_v1_1 [1]), .Z(MCInst2_MC2_r1Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst2_MC2_r1Inst_XORInst_0_2_U3  ( .A(
        MCInst2_MC2_r1Inst_XORInst_0_2_n5 ), .B(
        MCInst2_MC2_r1Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[38]) );
  XNOR2_X1 MCInst2_MC2_r1Inst_XORInst_0_2_U2  ( .A(MCInst2_MC2_v3_1 [2]), 
        .B(MCInst2_MC2_v2_1 [2]), .ZN(MCInst2_MC2_r1Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst2_MC2_r1Inst_XORInst_0_2_U1  ( .A(MCInst2_MC2_v0_1 [2]), .B(
        MCInst2_MC2_v1_1 [2]), .Z(MCInst2_MC2_r1Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst2_MC2_r1Inst_XORInst_0_3_U3  ( .A(
        MCInst2_MC2_r1Inst_XORInst_0_3_n5 ), .B(
        MCInst2_MC2_r1Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[39]) );
  XNOR2_X1 MCInst2_MC2_r1Inst_XORInst_0_3_U2  ( .A(MCInst2_MC2_v3_1 [3]), 
        .B(MCInst2_MC2_v2_1 [3]), .ZN(MCInst2_MC2_r1Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst2_MC2_r1Inst_XORInst_0_3_U1  ( .A(MCInst2_MC2_v0_1 [3]), .B(
        MCInst2_MC2_v1_1 [3]), .Z(MCInst2_MC2_r1Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst2_MC2_r2Inst_XORInst_0_0_U3  ( .A(
        MCInst2_MC2_r2Inst_XORInst_0_0_n5 ), .B(
        MCInst2_MC2_r2Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[20]) );
  XNOR2_X1 MCInst2_MC2_r2Inst_XORInst_0_0_U2  ( .A(MCInst2_MC2_v3_2 [0]), 
        .B(MCInst2_MC2_v2_2 [0]), .ZN(MCInst2_MC2_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst2_MC2_r2Inst_XORInst_0_0_U1  ( .A(MCInst2_MC2_v0_2 [0]), .B(
        MCInst2_MC2_v1_2 [0]), .Z(MCInst2_MC2_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst2_MC2_r2Inst_XORInst_0_1_U3  ( .A(
        MCInst2_MC2_r2Inst_XORInst_0_1_n5 ), .B(
        MCInst2_MC2_r2Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[21]) );
  XNOR2_X1 MCInst2_MC2_r2Inst_XORInst_0_1_U2  ( .A(MCInst2_MC2_v3_0 [3]), 
        .B(MCInst2_MC2_v2_2 [1]), .ZN(MCInst2_MC2_r2Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst2_MC2_r2Inst_XORInst_0_1_U1  ( .A(MCInst2_MC2_v0_2 [1]), .B(
        MCInst2_MC2_v1_2 [1]), .Z(MCInst2_MC2_r2Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst2_MC2_r2Inst_XORInst_0_2_U3  ( .A(
        MCInst2_MC2_r2Inst_XORInst_0_2_n5 ), .B(
        MCInst2_MC2_r2Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[22]) );
  XNOR2_X1 MCInst2_MC2_r2Inst_XORInst_0_2_U2  ( .A(MCInst2_MC2_v3_2 [2]), 
        .B(MCInst2_MC2_v2_2 [2]), .ZN(MCInst2_MC2_r2Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst2_MC2_r2Inst_XORInst_0_2_U1  ( .A(MCInst2_MC2_v0_2 [2]), .B(
        MCInst2_MC2_v1_2 [2]), .Z(MCInst2_MC2_r2Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst2_MC2_r2Inst_XORInst_0_3_U3  ( .A(
        MCInst2_MC2_r2Inst_XORInst_0_3_n5 ), .B(
        MCInst2_MC2_r2Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[23]) );
  XNOR2_X1 MCInst2_MC2_r2Inst_XORInst_0_3_U2  ( .A(MCInst2_MC2_v3_2 [3]), 
        .B(MCInst2_MC2_v2_2 [3]), .ZN(MCInst2_MC2_r2Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst2_MC2_r2Inst_XORInst_0_3_U1  ( .A(MCInst2_MC2_v0_2 [3]), .B(
        MCInst2_MC2_v1_2 [3]), .Z(MCInst2_MC2_r2Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst2_MC2_r3Inst_XORInst_0_0_U3  ( .A(
        MCInst2_MC2_r3Inst_XORInst_0_0_n5 ), .B(
        MCInst2_MC2_r3Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[4]) );
  XNOR2_X1 MCInst2_MC2_r3Inst_XORInst_0_0_U2  ( .A(MCInst2_MC2_v3_3 [0]), 
        .B(MCInst2_MC2_v2_3 [0]), .ZN(MCInst2_MC2_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst2_MC2_r3Inst_XORInst_0_0_U1  ( .A(MCInst2_MC2_v0_3 [0]), .B(
        MCInst2_MC2_v1_3 [0]), .Z(MCInst2_MC2_r3Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst2_MC2_r3Inst_XORInst_0_1_U3  ( .A(
        MCInst2_MC2_r3Inst_XORInst_0_1_n5 ), .B(
        MCInst2_MC2_r3Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[5]) );
  XNOR2_X1 MCInst2_MC2_r3Inst_XORInst_0_1_U2  ( .A(MCInst2_MC2_v3_3 [1]), 
        .B(MCInst2_MC2_v2_3 [1]), .ZN(MCInst2_MC2_r3Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst2_MC2_r3Inst_XORInst_0_1_U1  ( .A(MCInst2_MC2_v0_3 [1]), .B(
        MCInst2_MC2_v1_3 [1]), .Z(MCInst2_MC2_r3Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst2_MC2_r3Inst_XORInst_0_2_U3  ( .A(
        MCInst2_MC2_r3Inst_XORInst_0_2_n5 ), .B(
        MCInst2_MC2_r3Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[6]) );
  XNOR2_X1 MCInst2_MC2_r3Inst_XORInst_0_2_U2  ( .A(MCInst2_MC2_v3_3 [2]), 
        .B(MCInst2_MC2_v2_3 [2]), .ZN(MCInst2_MC2_r3Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst2_MC2_r3Inst_XORInst_0_2_U1  ( .A(MCInst2_MC2_v0_0 [3]), .B(
        MCInst2_MC2_v1_3 [2]), .Z(MCInst2_MC2_r3Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst2_MC2_r3Inst_XORInst_0_3_U3  ( .A(
        MCInst2_MC2_r3Inst_XORInst_0_3_n5 ), .B(
        MCInst2_MC2_r3Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[7]) );
  XNOR2_X1 MCInst2_MC2_r3Inst_XORInst_0_3_U2  ( .A(MCInst2_MC2_v3_3 [3]), 
        .B(MCInst2_MC2_v2_3 [3]), .ZN(MCInst2_MC2_r3Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst2_MC2_r3Inst_XORInst_0_3_U1  ( .A(MCInst2_MC2_v0_3 [3]), .B(
        MCInst2_MC2_v1_3 [3]), .Z(MCInst2_MC2_r3Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst2_MC3_v0_2Inst_0_U4  ( .A(MCInst2_MC3_v0_2Inst_0_n2 ), .B(
        MCInst2_MC3_v0_0 [3]), .ZN(MCInst2_MC3_v0_2 [0]) );
  XNOR2_X1 MCInst2_MC3_v0_2Inst_0_U3  ( .A(MCInst2_MC3_v0_3 [0]), .B(
        ShiftRowsOutput2[48]), .ZN(MCInst2_MC3_v0_2Inst_0_n2 ) );
  XOR2_X1 MCInst2_MC3_v1_1Inst_0_U3  ( .A(MCInst2_MC3_v1_3 [3]), .B(
        MCInst2_MC3_v1_3 [0]), .Z(MCInst2_MC3_v1_1 [0]) );
  XNOR2_X1 MCInst2_MC3_v1_2Inst_0_U4  ( .A(MCInst2_MC3_v1_2Inst_0_n2 ), .B(
        MCInst2_MC3_v1_3 [3]), .ZN(MCInst2_MC3_v1_2 [0]) );
  XNOR2_X1 MCInst2_MC3_v1_2Inst_0_U3  ( .A(MCInst2_MC3_v1_3 [0]), .B(
        MCInst2_MC3_v1_3 [2]), .ZN(MCInst2_MC3_v1_2Inst_0_n2 ) );
  XOR2_X1 MCInst2_MC3_v2_1Inst_0_U3  ( .A(MCInst2_MC3_v2_3 [1]), .B(
        MCInst2_MC3_v2_0 [3]), .Z(MCInst2_MC3_v2_1 [0]) );
  XOR2_X1 MCInst2_MC3_v2_2Inst_0_U3  ( .A(MCInst2_MC3_v2_0 [2]), .B(
        MCInst2_MC3_v2_0 [0]), .Z(MCInst2_MC3_v2_2 [0]) );
  XNOR2_X1 MCInst2_MC3_v2_3Inst_0_U5  ( .A(MCInst2_MC3_v2_3Inst_0_n4 ), .B(
        MCInst2_MC3_v2_3Inst_0_n3 ), .ZN(MCInst2_MC3_v2_3 [0]) );
  XNOR2_X1 MCInst2_MC3_v2_3Inst_0_U4  ( .A(MCInst2_MC3_v2_0 [2]), .B(
        MCInst2_MC3_v2_3 [1]), .ZN(MCInst2_MC3_v2_3Inst_0_n3 ) );
  XOR2_X1 MCInst2_MC3_v2_3Inst_0_U3  ( .A(MCInst2_MC3_v2_0 [3]), .B(
        MCInst2_MC3_v2_0 [0]), .Z(MCInst2_MC3_v2_3Inst_0_n4 ) );
  XOR2_X1 MCInst2_MC3_v3_1Inst_0_U3  ( .A(MCInst2_MC3_v3_0 [3]), .B(
        MCInst2_MC3_v3_2 [2]), .Z(MCInst2_MC3_v3_1 [0]) );
  XOR2_X1 MCInst2_MC3_v3_2Inst_0_U3  ( .A(MCInst2_MC3_v3_2 [3]), .B(
        MCInst2_MC3_v3_0 [2]), .Z(MCInst2_MC3_v3_2 [0]) );
  XNOR2_X1 MCInst2_MC3_v3_3Inst_0_U4  ( .A(MCInst2_MC3_v3_3Inst_0_n2 ), .B(
        MCInst2_MC3_v3_0 [2]), .ZN(MCInst2_MC3_v3_3 [0]) );
  XNOR2_X1 MCInst2_MC3_v3_3Inst_0_U3  ( .A(MCInst2_MC3_v3_2 [2]), .B(
        MCInst2_MC3_v3_2 [3]), .ZN(MCInst2_MC3_v3_3Inst_0_n2 ) );
  XOR2_X1 MCInst2_MC3_v0_0Inst_1_U3  ( .A(MCInst2_MC3_v0_3 [3]), .B(
        MCInst2_MC3_v0_3 [0]), .Z(MCInst2_MC3_v0_0 [1]) );
  XOR2_X1 MCInst2_MC3_v0_1Inst_1_U3  ( .A(MCInst2_MC3_v0_0 [3]), .B(
        MCInst2_MC3_v0_3 [3]), .Z(MCInst2_MC3_v0_1 [1]) );
  XNOR2_X1 MCInst2_MC3_v0_2Inst_1_U4  ( .A(MCInst2_MC3_v0_2Inst_1_n2 ), .B(
        MCInst2_MC3_v0_3 [3]), .ZN(MCInst2_MC3_v0_2 [1]) );
  XNOR2_X1 MCInst2_MC3_v0_2Inst_1_U3  ( .A(MCInst2_MC3_v0_3 [0]), .B(
        ShiftRowsOutput2[48]), .ZN(MCInst2_MC3_v0_2Inst_1_n2 ) );
  XOR2_X1 MCInst2_MC3_v0_3Inst_1_U3  ( .A(ShiftRowsOutput2[48]), .B(
        MCInst2_MC3_v0_3 [0]), .Z(MCInst2_MC3_v0_3 [1]) );
  XOR2_X1 MCInst2_MC3_v1_1Inst_1_U3  ( .A(ShiftRowsOutput2[32]), .B(
        MCInst2_MC3_v1_3 [3]), .Z(MCInst2_MC3_v1_1 [1]) );
  XOR2_X1 MCInst2_MC3_v1_2Inst_1_U3  ( .A(ShiftRowsOutput2[32]), .B(
        MCInst2_MC3_v1_3 [2]), .Z(MCInst2_MC3_v1_2 [1]) );
  XOR2_X1 MCInst2_MC3_v1_3Inst_1_U3  ( .A(ShiftRowsOutput2[32]), .B(
        MCInst2_MC3_v1_3 [0]), .Z(MCInst2_MC3_v1_3 [1]) );
  XOR2_X1 MCInst2_MC3_v2_0Inst_1_U3  ( .A(MCInst2_MC3_v2_3 [1]), .B(
        MCInst2_MC3_v2_0 [0]), .Z(MCInst2_MC3_v2_0 [1]) );
  XNOR2_X1 MCInst2_MC3_v2_1Inst_1_U4  ( .A(MCInst2_MC3_v2_1Inst_1_n2 ), .B(
        MCInst2_MC3_v2_0 [3]), .ZN(MCInst2_MC3_v2_1 [1]) );
  XNOR2_X1 MCInst2_MC3_v2_1Inst_1_U3  ( .A(MCInst2_MC3_v2_0 [0]), .B(
        MCInst2_MC3_v2_0 [2]), .ZN(MCInst2_MC3_v2_1Inst_1_n2 ) );
  XNOR2_X1 MCInst2_MC3_v2_2Inst_1_U5  ( .A(MCInst2_MC3_v2_2Inst_1_n4 ), .B(
        MCInst2_MC3_v2_2Inst_1_n3 ), .ZN(MCInst2_MC3_v2_2 [1]) );
  XNOR2_X1 MCInst2_MC3_v2_2Inst_1_U4  ( .A(MCInst2_MC3_v2_0 [2]), .B(
        MCInst2_MC3_v2_3 [1]), .ZN(MCInst2_MC3_v2_2Inst_1_n3 ) );
  XOR2_X1 MCInst2_MC3_v2_2Inst_1_U3  ( .A(MCInst2_MC3_v2_0 [3]), .B(
        MCInst2_MC3_v2_0 [0]), .Z(MCInst2_MC3_v2_2Inst_1_n4 ) );
  XOR2_X1 MCInst2_MC3_v3_0Inst_1_U3  ( .A(MCInst2_MC3_v3_2 [3]), .B(
        MCInst2_MC3_v3_2 [2]), .Z(MCInst2_MC3_v3_0 [1]) );
  XOR2_X1 MCInst2_MC3_v3_1Inst_1_U3  ( .A(MCInst2_MC3_v3_2 [3]), .B(
        MCInst2_MC3_v3_0 [3]), .Z(MCInst2_MC3_v3_1 [1]) );
  XNOR2_X1 MCInst2_MC3_v3_3Inst_1_U4  ( .A(MCInst2_MC3_v3_3Inst_1_n2 ), .B(
        MCInst2_MC3_v3_0 [3]), .ZN(MCInst2_MC3_v3_3 [1]) );
  XNOR2_X1 MCInst2_MC3_v3_3Inst_1_U3  ( .A(MCInst2_MC3_v3_2 [2]), .B(
        MCInst2_MC3_v3_2 [3]), .ZN(MCInst2_MC3_v3_3Inst_1_n2 ) );
  XOR2_X1 MCInst2_MC3_v0_0Inst_2_U3  ( .A(ShiftRowsOutput2[48]), .B(
        MCInst2_MC3_v0_3 [0]), .Z(MCInst2_MC3_v0_0 [2]) );
  XOR2_X1 MCInst2_MC3_v0_1Inst_2_U3  ( .A(MCInst2_MC3_v0_3 [3]), .B(
        MCInst2_MC3_v0_3 [0]), .Z(MCInst2_MC3_v0_1 [2]) );
  XOR2_X1 MCInst2_MC3_v0_2Inst_2_U3  ( .A(MCInst2_MC3_v0_0 [3]), .B(
        MCInst2_MC3_v0_3 [0]), .Z(MCInst2_MC3_v0_2 [2]) );
  XNOR2_X1 MCInst2_MC3_v1_1Inst_2_U4  ( .A(MCInst2_MC3_v1_1Inst_2_n2 ), .B(
        MCInst2_MC3_v1_3 [2]), .ZN(MCInst2_MC3_v1_1 [2]) );
  XNOR2_X1 MCInst2_MC3_v1_1Inst_2_U3  ( .A(MCInst2_MC3_v1_3 [0]), .B(
        ShiftRowsOutput2[32]), .ZN(MCInst2_MC3_v1_1Inst_2_n2 ) );
  XNOR2_X1 MCInst2_MC3_v1_2Inst_2_U4  ( .A(MCInst2_MC3_v1_2Inst_2_n2 ), .B(
        MCInst2_MC3_v1_3 [2]), .ZN(MCInst2_MC3_v1_2 [2]) );
  XNOR2_X1 MCInst2_MC3_v1_2Inst_2_U3  ( .A(MCInst2_MC3_v1_3 [3]), .B(
        ShiftRowsOutput2[32]), .ZN(MCInst2_MC3_v1_2Inst_2_n2 ) );
  XNOR2_X1 MCInst2_MC3_v2_1Inst_2_U4  ( .A(MCInst2_MC3_v2_1Inst_2_n2 ), .B(
        MCInst2_MC3_v2_0 [3]), .ZN(MCInst2_MC3_v2_1 [2]) );
  XNOR2_X1 MCInst2_MC3_v2_1Inst_2_U3  ( .A(MCInst2_MC3_v2_0 [0]), .B(
        MCInst2_MC3_v2_3 [1]), .ZN(MCInst2_MC3_v2_1Inst_2_n2 ) );
  XNOR2_X1 MCInst2_MC3_v2_2Inst_2_U4  ( .A(MCInst2_MC3_v2_2Inst_2_n2 ), .B(
        MCInst2_MC3_v2_0 [3]), .ZN(MCInst2_MC3_v2_2 [2]) );
  XNOR2_X1 MCInst2_MC3_v2_2Inst_2_U3  ( .A(MCInst2_MC3_v2_0 [0]), .B(
        MCInst2_MC3_v2_0 [2]), .ZN(MCInst2_MC3_v2_2Inst_2_n2 ) );
  XOR2_X1 MCInst2_MC3_v2_3Inst_2_U3  ( .A(MCInst2_MC3_v2_3 [1]), .B(
        MCInst2_MC3_v2_0 [2]), .Z(MCInst2_MC3_v2_3 [2]) );
  XNOR2_X1 MCInst2_MC3_v3_1Inst_2_U4  ( .A(MCInst2_MC3_v3_1Inst_2_n2 ), .B(
        MCInst2_MC3_v3_0 [2]), .ZN(MCInst2_MC3_v3_1 [2]) );
  XNOR2_X1 MCInst2_MC3_v3_1Inst_2_U3  ( .A(MCInst2_MC3_v3_2 [2]), .B(
        MCInst2_MC3_v3_2 [3]), .ZN(MCInst2_MC3_v3_1Inst_2_n2 ) );
  XOR2_X1 MCInst2_MC3_v3_3Inst_2_U3  ( .A(MCInst2_MC3_v3_0 [2]), .B(
        MCInst2_MC3_v3_2 [2]), .Z(MCInst2_MC3_v3_3 [2]) );
  XOR2_X1 MCInst2_MC3_v0_1Inst_3_U3  ( .A(ShiftRowsOutput2[48]), .B(
        MCInst2_MC3_v0_3 [0]), .Z(MCInst2_MC3_v0_1 [3]) );
  XOR2_X1 MCInst2_MC3_v0_2Inst_3_U3  ( .A(ShiftRowsOutput2[48]), .B(
        MCInst2_MC3_v0_3 [3]), .Z(MCInst2_MC3_v0_2 [3]) );
  XOR2_X1 MCInst2_MC3_v1_1Inst_3_U3  ( .A(MCInst2_MC3_v1_3 [2]), .B(
        MCInst2_MC3_v1_3 [3]), .Z(MCInst2_MC3_v1_1 [3]) );
  XNOR2_X1 MCInst2_MC3_v1_2Inst_3_U5  ( .A(MCInst2_MC3_v1_2Inst_3_n4 ), .B(
        MCInst2_MC3_v1_2Inst_3_n3 ), .ZN(MCInst2_MC3_v1_2 [3]) );
  XNOR2_X1 MCInst2_MC3_v1_2Inst_3_U4  ( .A(MCInst2_MC3_v1_3 [2]), .B(
        ShiftRowsOutput2[32]), .ZN(MCInst2_MC3_v1_2Inst_3_n3 ) );
  XOR2_X1 MCInst2_MC3_v1_2Inst_3_U3  ( .A(MCInst2_MC3_v1_3 [3]), .B(
        MCInst2_MC3_v1_3 [0]), .Z(MCInst2_MC3_v1_2Inst_3_n4 ) );
  XOR2_X1 MCInst2_MC3_v2_1Inst_3_U3  ( .A(MCInst2_MC3_v2_0 [2]), .B(
        MCInst2_MC3_v2_0 [0]), .Z(MCInst2_MC3_v2_1 [3]) );
  XNOR2_X1 MCInst2_MC3_v2_2Inst_3_U4  ( .A(MCInst2_MC3_v2_2Inst_3_n2 ), .B(
        MCInst2_MC3_v2_0 [3]), .ZN(MCInst2_MC3_v2_2 [3]) );
  XNOR2_X1 MCInst2_MC3_v2_2Inst_3_U3  ( .A(MCInst2_MC3_v2_0 [0]), .B(
        MCInst2_MC3_v2_3 [1]), .ZN(MCInst2_MC3_v2_2Inst_3_n2 ) );
  XNOR2_X1 MCInst2_MC3_v2_3Inst_3_U4  ( .A(MCInst2_MC3_v2_3Inst_3_n2 ), .B(
        MCInst2_MC3_v2_0 [2]), .ZN(MCInst2_MC3_v2_3 [3]) );
  XNOR2_X1 MCInst2_MC3_v2_3Inst_3_U3  ( .A(MCInst2_MC3_v2_0 [3]), .B(
        MCInst2_MC3_v2_3 [1]), .ZN(MCInst2_MC3_v2_3Inst_3_n2 ) );
  XOR2_X1 MCInst2_MC3_v3_1Inst_3_U3  ( .A(MCInst2_MC3_v3_0 [2]), .B(
        MCInst2_MC3_v3_0 [3]), .Z(MCInst2_MC3_v3_1 [3]) );
  XOR2_X1 MCInst2_MC3_v3_3Inst_3_U3  ( .A(MCInst2_MC3_v3_2 [3]), .B(
        MCInst2_MC3_v3_0 [3]), .Z(MCInst2_MC3_v3_3 [3]) );
  XNOR2_X1 MCInst2_MC3_r0Inst_XORInst_0_0_U3  ( .A(
        MCInst2_MC3_r0Inst_XORInst_0_0_n5 ), .B(
        MCInst2_MC3_r0Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[48]) );
  XNOR2_X1 MCInst2_MC3_r0Inst_XORInst_0_0_U2  ( .A(MCInst2_MC3_v3_2 [2]), 
        .B(MCInst2_MC3_v2_0 [0]), .ZN(MCInst2_MC3_r0Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst2_MC3_r0Inst_XORInst_0_0_U1  ( .A(MCInst2_MC3_v0_3 [3]), .B(
        ShiftRowsOutput2[32]), .Z(MCInst2_MC3_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst2_MC3_r0Inst_XORInst_0_1_U3  ( .A(
        MCInst2_MC3_r0Inst_XORInst_0_1_n5 ), .B(
        MCInst2_MC3_r0Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[49]) );
  XNOR2_X1 MCInst2_MC3_r0Inst_XORInst_0_1_U2  ( .A(MCInst2_MC3_v3_0 [1]), 
        .B(MCInst2_MC3_v2_0 [1]), .ZN(MCInst2_MC3_r0Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst2_MC3_r0Inst_XORInst_0_1_U1  ( .A(MCInst2_MC3_v0_0 [1]), .B(
        MCInst2_MC3_v1_3 [2]), .Z(MCInst2_MC3_r0Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst2_MC3_r0Inst_XORInst_0_2_U3  ( .A(
        MCInst2_MC3_r0Inst_XORInst_0_2_n5 ), .B(
        MCInst2_MC3_r0Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[50]) );
  XNOR2_X1 MCInst2_MC3_r0Inst_XORInst_0_2_U2  ( .A(MCInst2_MC3_v3_0 [2]), 
        .B(MCInst2_MC3_v2_0 [2]), .ZN(MCInst2_MC3_r0Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst2_MC3_r0Inst_XORInst_0_2_U1  ( .A(MCInst2_MC3_v0_0 [2]), .B(
        MCInst2_MC3_v1_3 [3]), .Z(MCInst2_MC3_r0Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst2_MC3_r0Inst_XORInst_0_3_U3  ( .A(
        MCInst2_MC3_r0Inst_XORInst_0_3_n5 ), .B(
        MCInst2_MC3_r0Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[51]) );
  XNOR2_X1 MCInst2_MC3_r0Inst_XORInst_0_3_U2  ( .A(MCInst2_MC3_v3_0 [3]), 
        .B(MCInst2_MC3_v2_0 [3]), .ZN(MCInst2_MC3_r0Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst2_MC3_r0Inst_XORInst_0_3_U1  ( .A(MCInst2_MC3_v0_0 [3]), .B(
        MCInst2_MC3_v1_3 [0]), .Z(MCInst2_MC3_r0Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst2_MC3_r1Inst_XORInst_0_0_U3  ( .A(
        MCInst2_MC3_r1Inst_XORInst_0_0_n5 ), .B(
        MCInst2_MC3_r1Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[32]) );
  XNOR2_X1 MCInst2_MC3_r1Inst_XORInst_0_0_U2  ( .A(MCInst2_MC3_v3_1 [0]), 
        .B(MCInst2_MC3_v2_1 [0]), .ZN(MCInst2_MC3_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst2_MC3_r1Inst_XORInst_0_0_U1  ( .A(MCInst2_MC3_v0_0 [3]), .B(
        MCInst2_MC3_v1_1 [0]), .Z(MCInst2_MC3_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst2_MC3_r1Inst_XORInst_0_1_U3  ( .A(
        MCInst2_MC3_r1Inst_XORInst_0_1_n5 ), .B(
        MCInst2_MC3_r1Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[33]) );
  XNOR2_X1 MCInst2_MC3_r1Inst_XORInst_0_1_U2  ( .A(MCInst2_MC3_v3_1 [1]), 
        .B(MCInst2_MC3_v2_1 [1]), .ZN(MCInst2_MC3_r1Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst2_MC3_r1Inst_XORInst_0_1_U1  ( .A(MCInst2_MC3_v0_1 [1]), .B(
        MCInst2_MC3_v1_1 [1]), .Z(MCInst2_MC3_r1Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst2_MC3_r1Inst_XORInst_0_2_U3  ( .A(
        MCInst2_MC3_r1Inst_XORInst_0_2_n5 ), .B(
        MCInst2_MC3_r1Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[34]) );
  XNOR2_X1 MCInst2_MC3_r1Inst_XORInst_0_2_U2  ( .A(MCInst2_MC3_v3_1 [2]), 
        .B(MCInst2_MC3_v2_1 [2]), .ZN(MCInst2_MC3_r1Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst2_MC3_r1Inst_XORInst_0_2_U1  ( .A(MCInst2_MC3_v0_1 [2]), .B(
        MCInst2_MC3_v1_1 [2]), .Z(MCInst2_MC3_r1Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst2_MC3_r1Inst_XORInst_0_3_U3  ( .A(
        MCInst2_MC3_r1Inst_XORInst_0_3_n5 ), .B(
        MCInst2_MC3_r1Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[35]) );
  XNOR2_X1 MCInst2_MC3_r1Inst_XORInst_0_3_U2  ( .A(MCInst2_MC3_v3_1 [3]), 
        .B(MCInst2_MC3_v2_1 [3]), .ZN(MCInst2_MC3_r1Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst2_MC3_r1Inst_XORInst_0_3_U1  ( .A(MCInst2_MC3_v0_1 [3]), .B(
        MCInst2_MC3_v1_1 [3]), .Z(MCInst2_MC3_r1Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst2_MC3_r2Inst_XORInst_0_0_U3  ( .A(
        MCInst2_MC3_r2Inst_XORInst_0_0_n5 ), .B(
        MCInst2_MC3_r2Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[16]) );
  XNOR2_X1 MCInst2_MC3_r2Inst_XORInst_0_0_U2  ( .A(MCInst2_MC3_v3_2 [0]), 
        .B(MCInst2_MC3_v2_2 [0]), .ZN(MCInst2_MC3_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst2_MC3_r2Inst_XORInst_0_0_U1  ( .A(MCInst2_MC3_v0_2 [0]), .B(
        MCInst2_MC3_v1_2 [0]), .Z(MCInst2_MC3_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst2_MC3_r2Inst_XORInst_0_1_U3  ( .A(
        MCInst2_MC3_r2Inst_XORInst_0_1_n5 ), .B(
        MCInst2_MC3_r2Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[17]) );
  XNOR2_X1 MCInst2_MC3_r2Inst_XORInst_0_1_U2  ( .A(MCInst2_MC3_v3_0 [3]), 
        .B(MCInst2_MC3_v2_2 [1]), .ZN(MCInst2_MC3_r2Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst2_MC3_r2Inst_XORInst_0_1_U1  ( .A(MCInst2_MC3_v0_2 [1]), .B(
        MCInst2_MC3_v1_2 [1]), .Z(MCInst2_MC3_r2Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst2_MC3_r2Inst_XORInst_0_2_U3  ( .A(
        MCInst2_MC3_r2Inst_XORInst_0_2_n5 ), .B(
        MCInst2_MC3_r2Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[18]) );
  XNOR2_X1 MCInst2_MC3_r2Inst_XORInst_0_2_U2  ( .A(MCInst2_MC3_v3_2 [2]), 
        .B(MCInst2_MC3_v2_2 [2]), .ZN(MCInst2_MC3_r2Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst2_MC3_r2Inst_XORInst_0_2_U1  ( .A(MCInst2_MC3_v0_2 [2]), .B(
        MCInst2_MC3_v1_2 [2]), .Z(MCInst2_MC3_r2Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst2_MC3_r2Inst_XORInst_0_3_U3  ( .A(
        MCInst2_MC3_r2Inst_XORInst_0_3_n5 ), .B(
        MCInst2_MC3_r2Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[19]) );
  XNOR2_X1 MCInst2_MC3_r2Inst_XORInst_0_3_U2  ( .A(MCInst2_MC3_v3_2 [3]), 
        .B(MCInst2_MC3_v2_2 [3]), .ZN(MCInst2_MC3_r2Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst2_MC3_r2Inst_XORInst_0_3_U1  ( .A(MCInst2_MC3_v0_2 [3]), .B(
        MCInst2_MC3_v1_2 [3]), .Z(MCInst2_MC3_r2Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst2_MC3_r3Inst_XORInst_0_0_U3  ( .A(
        MCInst2_MC3_r3Inst_XORInst_0_0_n5 ), .B(
        MCInst2_MC3_r3Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[0]) );
  XNOR2_X1 MCInst2_MC3_r3Inst_XORInst_0_0_U2  ( .A(MCInst2_MC3_v3_3 [0]), 
        .B(MCInst2_MC3_v2_3 [0]), .ZN(MCInst2_MC3_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst2_MC3_r3Inst_XORInst_0_0_U1  ( .A(MCInst2_MC3_v0_3 [0]), .B(
        MCInst2_MC3_v1_3 [0]), .Z(MCInst2_MC3_r3Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst2_MC3_r3Inst_XORInst_0_1_U3  ( .A(
        MCInst2_MC3_r3Inst_XORInst_0_1_n5 ), .B(
        MCInst2_MC3_r3Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[1]) );
  XNOR2_X1 MCInst2_MC3_r3Inst_XORInst_0_1_U2  ( .A(MCInst2_MC3_v3_3 [1]), 
        .B(MCInst2_MC3_v2_3 [1]), .ZN(MCInst2_MC3_r3Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst2_MC3_r3Inst_XORInst_0_1_U1  ( .A(MCInst2_MC3_v0_3 [1]), .B(
        MCInst2_MC3_v1_3 [1]), .Z(MCInst2_MC3_r3Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst2_MC3_r3Inst_XORInst_0_2_U3  ( .A(
        MCInst2_MC3_r3Inst_XORInst_0_2_n5 ), .B(
        MCInst2_MC3_r3Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[2]) );
  XNOR2_X1 MCInst2_MC3_r3Inst_XORInst_0_2_U2  ( .A(MCInst2_MC3_v3_3 [2]), 
        .B(MCInst2_MC3_v2_3 [2]), .ZN(MCInst2_MC3_r3Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst2_MC3_r3Inst_XORInst_0_2_U1  ( .A(MCInst2_MC3_v0_0 [3]), .B(
        MCInst2_MC3_v1_3 [2]), .Z(MCInst2_MC3_r3Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst2_MC3_r3Inst_XORInst_0_3_U3  ( .A(
        MCInst2_MC3_r3Inst_XORInst_0_3_n5 ), .B(
        MCInst2_MC3_r3Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[3]) );
  XNOR2_X1 MCInst2_MC3_r3Inst_XORInst_0_3_U2  ( .A(MCInst2_MC3_v3_3 [3]), 
        .B(MCInst2_MC3_v2_3 [3]), .ZN(MCInst2_MC3_r3Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst2_MC3_r3Inst_XORInst_0_3_U1  ( .A(MCInst2_MC3_v0_3 [3]), .B(
        MCInst2_MC3_v1_3 [3]), .Z(MCInst2_MC3_r3Inst_XORInst_0_3_n5 ) );
endmodule

