module Cipher ( clk, rst, EncDec, Input, Key, Tweak, Output, ErrorFlag );
  input [63:0] Input;
  input [191:0] Key;
  output [63:0] Output;
  (* FIRMER="clock" *)input clk;
  (* FIRMER="control" *)input rst;
  output ErrorFlag;
  wire   n8, n9, \MCInst_XOR_r0_Inst_0_n3 , \MCInst_XOR_r0_Inst_1_n3 ,
         \MCInst_XOR_r0_Inst_2_n3 , \MCInst_XOR_r0_Inst_3_n3 ,
         \MCInst_XOR_r0_Inst_4_n3 , \MCInst_XOR_r0_Inst_5_n3 ,
         \MCInst_XOR_r0_Inst_6_n3 , \MCInst_XOR_r0_Inst_7_n3 ,
         \MCInst_XOR_r0_Inst_8_n3 , \MCInst_XOR_r0_Inst_9_n3 ,
         \MCInst_XOR_r0_Inst_10_n3 , \MCInst_XOR_r0_Inst_11_n3 ,
         \MCInst_XOR_r0_Inst_12_n3 , \MCInst_XOR_r0_Inst_13_n3 ,
         \MCInst_XOR_r0_Inst_14_n3 , \MCInst_XOR_r0_Inst_15_n3 ,
         \SubCellInst_LFInst_0_LFInst_0_n11 ,
         \SubCellInst_LFInst_0_LFInst_0_n10 ,
         \SubCellInst_LFInst_0_LFInst_0_n9 ,
         \SubCellInst_LFInst_0_LFInst_0_n8 ,
         \SubCellInst_LFInst_0_LFInst_0_n7 ,
         \SubCellInst_LFInst_0_LFInst_1_n6 ,
         \SubCellInst_LFInst_0_LFInst_1_n5 ,
         \SubCellInst_LFInst_0_LFInst_1_n4 ,
         \SubCellInst_LFInst_0_LFInst_2_n11 ,
         \SubCellInst_LFInst_0_LFInst_2_n10 ,
         \SubCellInst_LFInst_0_LFInst_2_n9 ,
         \SubCellInst_LFInst_0_LFInst_2_n8 ,
         \SubCellInst_LFInst_0_LFInst_2_n7 ,
         \SubCellInst_LFInst_0_LFInst_3_n6 ,
         \SubCellInst_LFInst_0_LFInst_3_n5 ,
         \SubCellInst_LFInst_0_LFInst_3_n4 ,
         \SubCellInst_LFInst_1_LFInst_0_n11 ,
         \SubCellInst_LFInst_1_LFInst_0_n10 ,
         \SubCellInst_LFInst_1_LFInst_0_n9 ,
         \SubCellInst_LFInst_1_LFInst_0_n8 ,
         \SubCellInst_LFInst_1_LFInst_0_n7 ,
         \SubCellInst_LFInst_1_LFInst_1_n6 ,
         \SubCellInst_LFInst_1_LFInst_1_n5 ,
         \SubCellInst_LFInst_1_LFInst_1_n4 ,
         \SubCellInst_LFInst_1_LFInst_2_n11 ,
         \SubCellInst_LFInst_1_LFInst_2_n10 ,
         \SubCellInst_LFInst_1_LFInst_2_n9 ,
         \SubCellInst_LFInst_1_LFInst_2_n8 ,
         \SubCellInst_LFInst_1_LFInst_2_n7 ,
         \SubCellInst_LFInst_1_LFInst_3_n6 ,
         \SubCellInst_LFInst_1_LFInst_3_n5 ,
         \SubCellInst_LFInst_1_LFInst_3_n4 ,
         \SubCellInst_LFInst_2_LFInst_0_n11 ,
         \SubCellInst_LFInst_2_LFInst_0_n10 ,
         \SubCellInst_LFInst_2_LFInst_0_n9 ,
         \SubCellInst_LFInst_2_LFInst_0_n8 ,
         \SubCellInst_LFInst_2_LFInst_0_n7 ,
         \SubCellInst_LFInst_2_LFInst_1_n6 ,
         \SubCellInst_LFInst_2_LFInst_1_n5 ,
         \SubCellInst_LFInst_2_LFInst_1_n4 ,
         \SubCellInst_LFInst_2_LFInst_2_n11 ,
         \SubCellInst_LFInst_2_LFInst_2_n10 ,
         \SubCellInst_LFInst_2_LFInst_2_n9 ,
         \SubCellInst_LFInst_2_LFInst_2_n8 ,
         \SubCellInst_LFInst_2_LFInst_2_n7 ,
         \SubCellInst_LFInst_2_LFInst_3_n6 ,
         \SubCellInst_LFInst_2_LFInst_3_n5 ,
         \SubCellInst_LFInst_2_LFInst_3_n4 ,
         \SubCellInst_LFInst_3_LFInst_0_n11 ,
         \SubCellInst_LFInst_3_LFInst_0_n10 ,
         \SubCellInst_LFInst_3_LFInst_0_n9 ,
         \SubCellInst_LFInst_3_LFInst_0_n8 ,
         \SubCellInst_LFInst_3_LFInst_0_n7 ,
         \SubCellInst_LFInst_3_LFInst_1_n6 ,
         \SubCellInst_LFInst_3_LFInst_1_n5 ,
         \SubCellInst_LFInst_3_LFInst_1_n4 ,
         \SubCellInst_LFInst_3_LFInst_2_n11 ,
         \SubCellInst_LFInst_3_LFInst_2_n10 ,
         \SubCellInst_LFInst_3_LFInst_2_n9 ,
         \SubCellInst_LFInst_3_LFInst_2_n8 ,
         \SubCellInst_LFInst_3_LFInst_2_n7 ,
         \SubCellInst_LFInst_3_LFInst_3_n6 ,
         \SubCellInst_LFInst_3_LFInst_3_n5 ,
         \SubCellInst_LFInst_3_LFInst_3_n4 ,
         \SubCellInst_LFInst_4_LFInst_0_n11 ,
         \SubCellInst_LFInst_4_LFInst_0_n10 ,
         \SubCellInst_LFInst_4_LFInst_0_n9 ,
         \SubCellInst_LFInst_4_LFInst_0_n8 ,
         \SubCellInst_LFInst_4_LFInst_0_n7 ,
         \SubCellInst_LFInst_4_LFInst_1_n6 ,
         \SubCellInst_LFInst_4_LFInst_1_n5 ,
         \SubCellInst_LFInst_4_LFInst_1_n4 ,
         \SubCellInst_LFInst_4_LFInst_2_n11 ,
         \SubCellInst_LFInst_4_LFInst_2_n10 ,
         \SubCellInst_LFInst_4_LFInst_2_n9 ,
         \SubCellInst_LFInst_4_LFInst_2_n8 ,
         \SubCellInst_LFInst_4_LFInst_2_n7 ,
         \SubCellInst_LFInst_4_LFInst_3_n6 ,
         \SubCellInst_LFInst_4_LFInst_3_n5 ,
         \SubCellInst_LFInst_4_LFInst_3_n4 ,
         \SubCellInst_LFInst_5_LFInst_0_n11 ,
         \SubCellInst_LFInst_5_LFInst_0_n10 ,
         \SubCellInst_LFInst_5_LFInst_0_n9 ,
         \SubCellInst_LFInst_5_LFInst_0_n8 ,
         \SubCellInst_LFInst_5_LFInst_0_n7 ,
         \SubCellInst_LFInst_5_LFInst_1_n6 ,
         \SubCellInst_LFInst_5_LFInst_1_n5 ,
         \SubCellInst_LFInst_5_LFInst_1_n4 ,
         \SubCellInst_LFInst_5_LFInst_2_n11 ,
         \SubCellInst_LFInst_5_LFInst_2_n10 ,
         \SubCellInst_LFInst_5_LFInst_2_n9 ,
         \SubCellInst_LFInst_5_LFInst_2_n8 ,
         \SubCellInst_LFInst_5_LFInst_2_n7 ,
         \SubCellInst_LFInst_5_LFInst_3_n6 ,
         \SubCellInst_LFInst_5_LFInst_3_n5 ,
         \SubCellInst_LFInst_5_LFInst_3_n4 ,
         \SubCellInst_LFInst_6_LFInst_0_n11 ,
         \SubCellInst_LFInst_6_LFInst_0_n10 ,
         \SubCellInst_LFInst_6_LFInst_0_n9 ,
         \SubCellInst_LFInst_6_LFInst_0_n8 ,
         \SubCellInst_LFInst_6_LFInst_0_n7 ,
         \SubCellInst_LFInst_6_LFInst_1_n6 ,
         \SubCellInst_LFInst_6_LFInst_1_n5 ,
         \SubCellInst_LFInst_6_LFInst_1_n4 ,
         \SubCellInst_LFInst_6_LFInst_2_n11 ,
         \SubCellInst_LFInst_6_LFInst_2_n10 ,
         \SubCellInst_LFInst_6_LFInst_2_n9 ,
         \SubCellInst_LFInst_6_LFInst_2_n8 ,
         \SubCellInst_LFInst_6_LFInst_2_n7 ,
         \SubCellInst_LFInst_6_LFInst_3_n6 ,
         \SubCellInst_LFInst_6_LFInst_3_n5 ,
         \SubCellInst_LFInst_6_LFInst_3_n4 ,
         \SubCellInst_LFInst_7_LFInst_0_n11 ,
         \SubCellInst_LFInst_7_LFInst_0_n10 ,
         \SubCellInst_LFInst_7_LFInst_0_n9 ,
         \SubCellInst_LFInst_7_LFInst_0_n8 ,
         \SubCellInst_LFInst_7_LFInst_0_n7 ,
         \SubCellInst_LFInst_7_LFInst_1_n6 ,
         \SubCellInst_LFInst_7_LFInst_1_n5 ,
         \SubCellInst_LFInst_7_LFInst_1_n4 ,
         \SubCellInst_LFInst_7_LFInst_2_n11 ,
         \SubCellInst_LFInst_7_LFInst_2_n10 ,
         \SubCellInst_LFInst_7_LFInst_2_n9 ,
         \SubCellInst_LFInst_7_LFInst_2_n8 ,
         \SubCellInst_LFInst_7_LFInst_2_n7 ,
         \SubCellInst_LFInst_7_LFInst_3_n6 ,
         \SubCellInst_LFInst_7_LFInst_3_n5 ,
         \SubCellInst_LFInst_7_LFInst_3_n4 ,
         \SubCellInst_LFInst_8_LFInst_0_n11 ,
         \SubCellInst_LFInst_8_LFInst_0_n10 ,
         \SubCellInst_LFInst_8_LFInst_0_n9 ,
         \SubCellInst_LFInst_8_LFInst_0_n8 ,
         \SubCellInst_LFInst_8_LFInst_0_n7 ,
         \SubCellInst_LFInst_8_LFInst_1_n6 ,
         \SubCellInst_LFInst_8_LFInst_1_n5 ,
         \SubCellInst_LFInst_8_LFInst_1_n4 ,
         \SubCellInst_LFInst_8_LFInst_2_n11 ,
         \SubCellInst_LFInst_8_LFInst_2_n10 ,
         \SubCellInst_LFInst_8_LFInst_2_n9 ,
         \SubCellInst_LFInst_8_LFInst_2_n8 ,
         \SubCellInst_LFInst_8_LFInst_2_n7 ,
         \SubCellInst_LFInst_8_LFInst_3_n6 ,
         \SubCellInst_LFInst_8_LFInst_3_n5 ,
         \SubCellInst_LFInst_8_LFInst_3_n4 ,
         \SubCellInst_LFInst_9_LFInst_0_n11 ,
         \SubCellInst_LFInst_9_LFInst_0_n10 ,
         \SubCellInst_LFInst_9_LFInst_0_n9 ,
         \SubCellInst_LFInst_9_LFInst_0_n8 ,
         \SubCellInst_LFInst_9_LFInst_0_n7 ,
         \SubCellInst_LFInst_9_LFInst_1_n6 ,
         \SubCellInst_LFInst_9_LFInst_1_n5 ,
         \SubCellInst_LFInst_9_LFInst_1_n4 ,
         \SubCellInst_LFInst_9_LFInst_2_n11 ,
         \SubCellInst_LFInst_9_LFInst_2_n10 ,
         \SubCellInst_LFInst_9_LFInst_2_n9 ,
         \SubCellInst_LFInst_9_LFInst_2_n8 ,
         \SubCellInst_LFInst_9_LFInst_2_n7 ,
         \SubCellInst_LFInst_9_LFInst_3_n6 ,
         \SubCellInst_LFInst_9_LFInst_3_n5 ,
         \SubCellInst_LFInst_9_LFInst_3_n4 ,
         \SubCellInst_LFInst_10_LFInst_0_n11 ,
         \SubCellInst_LFInst_10_LFInst_0_n10 ,
         \SubCellInst_LFInst_10_LFInst_0_n9 ,
         \SubCellInst_LFInst_10_LFInst_0_n8 ,
         \SubCellInst_LFInst_10_LFInst_0_n7 ,
         \SubCellInst_LFInst_10_LFInst_1_n6 ,
         \SubCellInst_LFInst_10_LFInst_1_n5 ,
         \SubCellInst_LFInst_10_LFInst_1_n4 ,
         \SubCellInst_LFInst_10_LFInst_2_n11 ,
         \SubCellInst_LFInst_10_LFInst_2_n10 ,
         \SubCellInst_LFInst_10_LFInst_2_n9 ,
         \SubCellInst_LFInst_10_LFInst_2_n8 ,
         \SubCellInst_LFInst_10_LFInst_2_n7 ,
         \SubCellInst_LFInst_10_LFInst_3_n6 ,
         \SubCellInst_LFInst_10_LFInst_3_n5 ,
         \SubCellInst_LFInst_10_LFInst_3_n4 ,
         \SubCellInst_LFInst_11_LFInst_0_n11 ,
         \SubCellInst_LFInst_11_LFInst_0_n10 ,
         \SubCellInst_LFInst_11_LFInst_0_n9 ,
         \SubCellInst_LFInst_11_LFInst_0_n8 ,
         \SubCellInst_LFInst_11_LFInst_0_n7 ,
         \SubCellInst_LFInst_11_LFInst_1_n6 ,
         \SubCellInst_LFInst_11_LFInst_1_n5 ,
         \SubCellInst_LFInst_11_LFInst_1_n4 ,
         \SubCellInst_LFInst_11_LFInst_2_n11 ,
         \SubCellInst_LFInst_11_LFInst_2_n10 ,
         \SubCellInst_LFInst_11_LFInst_2_n9 ,
         \SubCellInst_LFInst_11_LFInst_2_n8 ,
         \SubCellInst_LFInst_11_LFInst_2_n7 ,
         \SubCellInst_LFInst_11_LFInst_3_n6 ,
         \SubCellInst_LFInst_11_LFInst_3_n5 ,
         \SubCellInst_LFInst_11_LFInst_3_n4 ,
         \SubCellInst_LFInst_12_LFInst_0_n11 ,
         \SubCellInst_LFInst_12_LFInst_0_n10 ,
         \SubCellInst_LFInst_12_LFInst_0_n9 ,
         \SubCellInst_LFInst_12_LFInst_0_n8 ,
         \SubCellInst_LFInst_12_LFInst_0_n7 ,
         \SubCellInst_LFInst_12_LFInst_1_n6 ,
         \SubCellInst_LFInst_12_LFInst_1_n5 ,
         \SubCellInst_LFInst_12_LFInst_1_n4 ,
         \SubCellInst_LFInst_12_LFInst_2_n11 ,
         \SubCellInst_LFInst_12_LFInst_2_n10 ,
         \SubCellInst_LFInst_12_LFInst_2_n9 ,
         \SubCellInst_LFInst_12_LFInst_2_n8 ,
         \SubCellInst_LFInst_12_LFInst_2_n7 ,
         \SubCellInst_LFInst_12_LFInst_3_n6 ,
         \SubCellInst_LFInst_12_LFInst_3_n5 ,
         \SubCellInst_LFInst_12_LFInst_3_n4 ,
         \SubCellInst_LFInst_13_LFInst_0_n11 ,
         \SubCellInst_LFInst_13_LFInst_0_n10 ,
         \SubCellInst_LFInst_13_LFInst_0_n9 ,
         \SubCellInst_LFInst_13_LFInst_0_n8 ,
         \SubCellInst_LFInst_13_LFInst_0_n7 ,
         \SubCellInst_LFInst_13_LFInst_1_n6 ,
         \SubCellInst_LFInst_13_LFInst_1_n5 ,
         \SubCellInst_LFInst_13_LFInst_1_n4 ,
         \SubCellInst_LFInst_13_LFInst_2_n11 ,
         \SubCellInst_LFInst_13_LFInst_2_n10 ,
         \SubCellInst_LFInst_13_LFInst_2_n9 ,
         \SubCellInst_LFInst_13_LFInst_2_n8 ,
         \SubCellInst_LFInst_13_LFInst_2_n7 ,
         \SubCellInst_LFInst_13_LFInst_3_n6 ,
         \SubCellInst_LFInst_13_LFInst_3_n5 ,
         \SubCellInst_LFInst_13_LFInst_3_n4 ,
         \SubCellInst_LFInst_14_LFInst_0_n11 ,
         \SubCellInst_LFInst_14_LFInst_0_n10 ,
         \SubCellInst_LFInst_14_LFInst_0_n9 ,
         \SubCellInst_LFInst_14_LFInst_0_n8 ,
         \SubCellInst_LFInst_14_LFInst_0_n7 ,
         \SubCellInst_LFInst_14_LFInst_1_n6 ,
         \SubCellInst_LFInst_14_LFInst_1_n5 ,
         \SubCellInst_LFInst_14_LFInst_1_n4 ,
         \SubCellInst_LFInst_14_LFInst_2_n11 ,
         \SubCellInst_LFInst_14_LFInst_2_n10 ,
         \SubCellInst_LFInst_14_LFInst_2_n9 ,
         \SubCellInst_LFInst_14_LFInst_2_n8 ,
         \SubCellInst_LFInst_14_LFInst_2_n7 ,
         \SubCellInst_LFInst_14_LFInst_3_n6 ,
         \SubCellInst_LFInst_14_LFInst_3_n5 ,
         \SubCellInst_LFInst_14_LFInst_3_n4 ,
         \SubCellInst_LFInst_15_LFInst_0_n11 ,
         \SubCellInst_LFInst_15_LFInst_0_n10 ,
         \SubCellInst_LFInst_15_LFInst_0_n9 ,
         \SubCellInst_LFInst_15_LFInst_0_n8 ,
         \SubCellInst_LFInst_15_LFInst_0_n7 ,
         \SubCellInst_LFInst_15_LFInst_1_n6 ,
         \SubCellInst_LFInst_15_LFInst_1_n5 ,
         \SubCellInst_LFInst_15_LFInst_1_n4 ,
         \SubCellInst_LFInst_15_LFInst_2_n11 ,
         \SubCellInst_LFInst_15_LFInst_2_n10 ,
         \SubCellInst_LFInst_15_LFInst_2_n9 ,
         \SubCellInst_LFInst_15_LFInst_2_n8 ,
         \SubCellInst_LFInst_15_LFInst_2_n7 ,
         \SubCellInst_LFInst_15_LFInst_3_n6 ,
         \SubCellInst_LFInst_15_LFInst_3_n5 ,
         \SubCellInst_LFInst_15_LFInst_3_n4 , \MCInst2_XOR_r0_Inst_0_n3 ,
         \MCInst2_XOR_r0_Inst_1_n3 , \MCInst2_XOR_r0_Inst_2_n3 ,
         \MCInst2_XOR_r0_Inst_3_n3 , \MCInst2_XOR_r0_Inst_4_n3 ,
         \MCInst2_XOR_r0_Inst_5_n3 , \MCInst2_XOR_r0_Inst_6_n3 ,
         \MCInst2_XOR_r0_Inst_7_n3 , \MCInst2_XOR_r0_Inst_8_n3 ,
         \MCInst2_XOR_r0_Inst_9_n3 , \MCInst2_XOR_r0_Inst_10_n3 ,
         \MCInst2_XOR_r0_Inst_11_n3 , \MCInst2_XOR_r0_Inst_12_n3 ,
         \MCInst2_XOR_r0_Inst_13_n3 , \MCInst2_XOR_r0_Inst_14_n3 ,
         \MCInst2_XOR_r0_Inst_15_n3 , \SubCellInst2_LFInst_0_LFInst_0_n11 ,
         \SubCellInst2_LFInst_0_LFInst_0_n10 ,
         \SubCellInst2_LFInst_0_LFInst_0_n9 ,
         \SubCellInst2_LFInst_0_LFInst_0_n8 ,
         \SubCellInst2_LFInst_0_LFInst_0_n7 ,
         \SubCellInst2_LFInst_0_LFInst_1_n6 ,
         \SubCellInst2_LFInst_0_LFInst_1_n5 ,
         \SubCellInst2_LFInst_0_LFInst_1_n4 ,
         \SubCellInst2_LFInst_0_LFInst_2_n11 ,
         \SubCellInst2_LFInst_0_LFInst_2_n10 ,
         \SubCellInst2_LFInst_0_LFInst_2_n9 ,
         \SubCellInst2_LFInst_0_LFInst_2_n8 ,
         \SubCellInst2_LFInst_0_LFInst_2_n7 ,
         \SubCellInst2_LFInst_0_LFInst_3_n6 ,
         \SubCellInst2_LFInst_0_LFInst_3_n5 ,
         \SubCellInst2_LFInst_0_LFInst_3_n4 ,
         \SubCellInst2_LFInst_1_LFInst_0_n11 ,
         \SubCellInst2_LFInst_1_LFInst_0_n10 ,
         \SubCellInst2_LFInst_1_LFInst_0_n9 ,
         \SubCellInst2_LFInst_1_LFInst_0_n8 ,
         \SubCellInst2_LFInst_1_LFInst_0_n7 ,
         \SubCellInst2_LFInst_1_LFInst_1_n6 ,
         \SubCellInst2_LFInst_1_LFInst_1_n5 ,
         \SubCellInst2_LFInst_1_LFInst_1_n4 ,
         \SubCellInst2_LFInst_1_LFInst_2_n11 ,
         \SubCellInst2_LFInst_1_LFInst_2_n10 ,
         \SubCellInst2_LFInst_1_LFInst_2_n9 ,
         \SubCellInst2_LFInst_1_LFInst_2_n8 ,
         \SubCellInst2_LFInst_1_LFInst_2_n7 ,
         \SubCellInst2_LFInst_1_LFInst_3_n6 ,
         \SubCellInst2_LFInst_1_LFInst_3_n5 ,
         \SubCellInst2_LFInst_1_LFInst_3_n4 ,
         \SubCellInst2_LFInst_2_LFInst_0_n11 ,
         \SubCellInst2_LFInst_2_LFInst_0_n10 ,
         \SubCellInst2_LFInst_2_LFInst_0_n9 ,
         \SubCellInst2_LFInst_2_LFInst_0_n8 ,
         \SubCellInst2_LFInst_2_LFInst_0_n7 ,
         \SubCellInst2_LFInst_2_LFInst_1_n6 ,
         \SubCellInst2_LFInst_2_LFInst_1_n5 ,
         \SubCellInst2_LFInst_2_LFInst_1_n4 ,
         \SubCellInst2_LFInst_2_LFInst_2_n11 ,
         \SubCellInst2_LFInst_2_LFInst_2_n10 ,
         \SubCellInst2_LFInst_2_LFInst_2_n9 ,
         \SubCellInst2_LFInst_2_LFInst_2_n8 ,
         \SubCellInst2_LFInst_2_LFInst_2_n7 ,
         \SubCellInst2_LFInst_2_LFInst_3_n6 ,
         \SubCellInst2_LFInst_2_LFInst_3_n5 ,
         \SubCellInst2_LFInst_2_LFInst_3_n4 ,
         \SubCellInst2_LFInst_3_LFInst_0_n11 ,
         \SubCellInst2_LFInst_3_LFInst_0_n10 ,
         \SubCellInst2_LFInst_3_LFInst_0_n9 ,
         \SubCellInst2_LFInst_3_LFInst_0_n8 ,
         \SubCellInst2_LFInst_3_LFInst_0_n7 ,
         \SubCellInst2_LFInst_3_LFInst_1_n6 ,
         \SubCellInst2_LFInst_3_LFInst_1_n5 ,
         \SubCellInst2_LFInst_3_LFInst_1_n4 ,
         \SubCellInst2_LFInst_3_LFInst_2_n11 ,
         \SubCellInst2_LFInst_3_LFInst_2_n10 ,
         \SubCellInst2_LFInst_3_LFInst_2_n9 ,
         \SubCellInst2_LFInst_3_LFInst_2_n8 ,
         \SubCellInst2_LFInst_3_LFInst_2_n7 ,
         \SubCellInst2_LFInst_3_LFInst_3_n6 ,
         \SubCellInst2_LFInst_3_LFInst_3_n5 ,
         \SubCellInst2_LFInst_3_LFInst_3_n4 ,
         \SubCellInst2_LFInst_4_LFInst_0_n11 ,
         \SubCellInst2_LFInst_4_LFInst_0_n10 ,
         \SubCellInst2_LFInst_4_LFInst_0_n9 ,
         \SubCellInst2_LFInst_4_LFInst_0_n8 ,
         \SubCellInst2_LFInst_4_LFInst_0_n7 ,
         \SubCellInst2_LFInst_4_LFInst_1_n6 ,
         \SubCellInst2_LFInst_4_LFInst_1_n5 ,
         \SubCellInst2_LFInst_4_LFInst_1_n4 ,
         \SubCellInst2_LFInst_4_LFInst_2_n11 ,
         \SubCellInst2_LFInst_4_LFInst_2_n10 ,
         \SubCellInst2_LFInst_4_LFInst_2_n9 ,
         \SubCellInst2_LFInst_4_LFInst_2_n8 ,
         \SubCellInst2_LFInst_4_LFInst_2_n7 ,
         \SubCellInst2_LFInst_4_LFInst_3_n6 ,
         \SubCellInst2_LFInst_4_LFInst_3_n5 ,
         \SubCellInst2_LFInst_4_LFInst_3_n4 ,
         \SubCellInst2_LFInst_5_LFInst_0_n11 ,
         \SubCellInst2_LFInst_5_LFInst_0_n10 ,
         \SubCellInst2_LFInst_5_LFInst_0_n9 ,
         \SubCellInst2_LFInst_5_LFInst_0_n8 ,
         \SubCellInst2_LFInst_5_LFInst_0_n7 ,
         \SubCellInst2_LFInst_5_LFInst_1_n6 ,
         \SubCellInst2_LFInst_5_LFInst_1_n5 ,
         \SubCellInst2_LFInst_5_LFInst_1_n4 ,
         \SubCellInst2_LFInst_5_LFInst_2_n11 ,
         \SubCellInst2_LFInst_5_LFInst_2_n10 ,
         \SubCellInst2_LFInst_5_LFInst_2_n9 ,
         \SubCellInst2_LFInst_5_LFInst_2_n8 ,
         \SubCellInst2_LFInst_5_LFInst_2_n7 ,
         \SubCellInst2_LFInst_5_LFInst_3_n6 ,
         \SubCellInst2_LFInst_5_LFInst_3_n5 ,
         \SubCellInst2_LFInst_5_LFInst_3_n4 ,
         \SubCellInst2_LFInst_6_LFInst_0_n11 ,
         \SubCellInst2_LFInst_6_LFInst_0_n10 ,
         \SubCellInst2_LFInst_6_LFInst_0_n9 ,
         \SubCellInst2_LFInst_6_LFInst_0_n8 ,
         \SubCellInst2_LFInst_6_LFInst_0_n7 ,
         \SubCellInst2_LFInst_6_LFInst_1_n6 ,
         \SubCellInst2_LFInst_6_LFInst_1_n5 ,
         \SubCellInst2_LFInst_6_LFInst_1_n4 ,
         \SubCellInst2_LFInst_6_LFInst_2_n11 ,
         \SubCellInst2_LFInst_6_LFInst_2_n10 ,
         \SubCellInst2_LFInst_6_LFInst_2_n9 ,
         \SubCellInst2_LFInst_6_LFInst_2_n8 ,
         \SubCellInst2_LFInst_6_LFInst_2_n7 ,
         \SubCellInst2_LFInst_6_LFInst_3_n6 ,
         \SubCellInst2_LFInst_6_LFInst_3_n5 ,
         \SubCellInst2_LFInst_6_LFInst_3_n4 ,
         \SubCellInst2_LFInst_7_LFInst_0_n11 ,
         \SubCellInst2_LFInst_7_LFInst_0_n10 ,
         \SubCellInst2_LFInst_7_LFInst_0_n9 ,
         \SubCellInst2_LFInst_7_LFInst_0_n8 ,
         \SubCellInst2_LFInst_7_LFInst_0_n7 ,
         \SubCellInst2_LFInst_7_LFInst_1_n6 ,
         \SubCellInst2_LFInst_7_LFInst_1_n5 ,
         \SubCellInst2_LFInst_7_LFInst_1_n4 ,
         \SubCellInst2_LFInst_7_LFInst_2_n11 ,
         \SubCellInst2_LFInst_7_LFInst_2_n10 ,
         \SubCellInst2_LFInst_7_LFInst_2_n9 ,
         \SubCellInst2_LFInst_7_LFInst_2_n8 ,
         \SubCellInst2_LFInst_7_LFInst_2_n7 ,
         \SubCellInst2_LFInst_7_LFInst_3_n6 ,
         \SubCellInst2_LFInst_7_LFInst_3_n5 ,
         \SubCellInst2_LFInst_7_LFInst_3_n4 ,
         \SubCellInst2_LFInst_8_LFInst_0_n11 ,
         \SubCellInst2_LFInst_8_LFInst_0_n10 ,
         \SubCellInst2_LFInst_8_LFInst_0_n9 ,
         \SubCellInst2_LFInst_8_LFInst_0_n8 ,
         \SubCellInst2_LFInst_8_LFInst_0_n7 ,
         \SubCellInst2_LFInst_8_LFInst_1_n6 ,
         \SubCellInst2_LFInst_8_LFInst_1_n5 ,
         \SubCellInst2_LFInst_8_LFInst_1_n4 ,
         \SubCellInst2_LFInst_8_LFInst_2_n11 ,
         \SubCellInst2_LFInst_8_LFInst_2_n10 ,
         \SubCellInst2_LFInst_8_LFInst_2_n9 ,
         \SubCellInst2_LFInst_8_LFInst_2_n8 ,
         \SubCellInst2_LFInst_8_LFInst_2_n7 ,
         \SubCellInst2_LFInst_8_LFInst_3_n6 ,
         \SubCellInst2_LFInst_8_LFInst_3_n5 ,
         \SubCellInst2_LFInst_8_LFInst_3_n4 ,
         \SubCellInst2_LFInst_9_LFInst_0_n11 ,
         \SubCellInst2_LFInst_9_LFInst_0_n10 ,
         \SubCellInst2_LFInst_9_LFInst_0_n9 ,
         \SubCellInst2_LFInst_9_LFInst_0_n8 ,
         \SubCellInst2_LFInst_9_LFInst_0_n7 ,
         \SubCellInst2_LFInst_9_LFInst_1_n6 ,
         \SubCellInst2_LFInst_9_LFInst_1_n5 ,
         \SubCellInst2_LFInst_9_LFInst_1_n4 ,
         \SubCellInst2_LFInst_9_LFInst_2_n11 ,
         \SubCellInst2_LFInst_9_LFInst_2_n10 ,
         \SubCellInst2_LFInst_9_LFInst_2_n9 ,
         \SubCellInst2_LFInst_9_LFInst_2_n8 ,
         \SubCellInst2_LFInst_9_LFInst_2_n7 ,
         \SubCellInst2_LFInst_9_LFInst_3_n6 ,
         \SubCellInst2_LFInst_9_LFInst_3_n5 ,
         \SubCellInst2_LFInst_9_LFInst_3_n4 ,
         \SubCellInst2_LFInst_10_LFInst_0_n11 ,
         \SubCellInst2_LFInst_10_LFInst_0_n10 ,
         \SubCellInst2_LFInst_10_LFInst_0_n9 ,
         \SubCellInst2_LFInst_10_LFInst_0_n8 ,
         \SubCellInst2_LFInst_10_LFInst_0_n7 ,
         \SubCellInst2_LFInst_10_LFInst_1_n6 ,
         \SubCellInst2_LFInst_10_LFInst_1_n5 ,
         \SubCellInst2_LFInst_10_LFInst_1_n4 ,
         \SubCellInst2_LFInst_10_LFInst_2_n11 ,
         \SubCellInst2_LFInst_10_LFInst_2_n10 ,
         \SubCellInst2_LFInst_10_LFInst_2_n9 ,
         \SubCellInst2_LFInst_10_LFInst_2_n8 ,
         \SubCellInst2_LFInst_10_LFInst_2_n7 ,
         \SubCellInst2_LFInst_10_LFInst_3_n6 ,
         \SubCellInst2_LFInst_10_LFInst_3_n5 ,
         \SubCellInst2_LFInst_10_LFInst_3_n4 ,
         \SubCellInst2_LFInst_11_LFInst_0_n11 ,
         \SubCellInst2_LFInst_11_LFInst_0_n10 ,
         \SubCellInst2_LFInst_11_LFInst_0_n9 ,
         \SubCellInst2_LFInst_11_LFInst_0_n8 ,
         \SubCellInst2_LFInst_11_LFInst_0_n7 ,
         \SubCellInst2_LFInst_11_LFInst_1_n6 ,
         \SubCellInst2_LFInst_11_LFInst_1_n5 ,
         \SubCellInst2_LFInst_11_LFInst_1_n4 ,
         \SubCellInst2_LFInst_11_LFInst_2_n11 ,
         \SubCellInst2_LFInst_11_LFInst_2_n10 ,
         \SubCellInst2_LFInst_11_LFInst_2_n9 ,
         \SubCellInst2_LFInst_11_LFInst_2_n8 ,
         \SubCellInst2_LFInst_11_LFInst_2_n7 ,
         \SubCellInst2_LFInst_11_LFInst_3_n6 ,
         \SubCellInst2_LFInst_11_LFInst_3_n5 ,
         \SubCellInst2_LFInst_11_LFInst_3_n4 ,
         \SubCellInst2_LFInst_12_LFInst_0_n11 ,
         \SubCellInst2_LFInst_12_LFInst_0_n10 ,
         \SubCellInst2_LFInst_12_LFInst_0_n9 ,
         \SubCellInst2_LFInst_12_LFInst_0_n8 ,
         \SubCellInst2_LFInst_12_LFInst_0_n7 ,
         \SubCellInst2_LFInst_12_LFInst_1_n6 ,
         \SubCellInst2_LFInst_12_LFInst_1_n5 ,
         \SubCellInst2_LFInst_12_LFInst_1_n4 ,
         \SubCellInst2_LFInst_12_LFInst_2_n11 ,
         \SubCellInst2_LFInst_12_LFInst_2_n10 ,
         \SubCellInst2_LFInst_12_LFInst_2_n9 ,
         \SubCellInst2_LFInst_12_LFInst_2_n8 ,
         \SubCellInst2_LFInst_12_LFInst_2_n7 ,
         \SubCellInst2_LFInst_12_LFInst_3_n6 ,
         \SubCellInst2_LFInst_12_LFInst_3_n5 ,
         \SubCellInst2_LFInst_12_LFInst_3_n4 ,
         \SubCellInst2_LFInst_13_LFInst_0_n11 ,
         \SubCellInst2_LFInst_13_LFInst_0_n10 ,
         \SubCellInst2_LFInst_13_LFInst_0_n9 ,
         \SubCellInst2_LFInst_13_LFInst_0_n8 ,
         \SubCellInst2_LFInst_13_LFInst_0_n7 ,
         \SubCellInst2_LFInst_13_LFInst_1_n6 ,
         \SubCellInst2_LFInst_13_LFInst_1_n5 ,
         \SubCellInst2_LFInst_13_LFInst_1_n4 ,
         \SubCellInst2_LFInst_13_LFInst_2_n11 ,
         \SubCellInst2_LFInst_13_LFInst_2_n10 ,
         \SubCellInst2_LFInst_13_LFInst_2_n9 ,
         \SubCellInst2_LFInst_13_LFInst_2_n8 ,
         \SubCellInst2_LFInst_13_LFInst_2_n7 ,
         \SubCellInst2_LFInst_13_LFInst_3_n6 ,
         \SubCellInst2_LFInst_13_LFInst_3_n5 ,
         \SubCellInst2_LFInst_13_LFInst_3_n4 ,
         \SubCellInst2_LFInst_14_LFInst_0_n11 ,
         \SubCellInst2_LFInst_14_LFInst_0_n10 ,
         \SubCellInst2_LFInst_14_LFInst_0_n9 ,
         \SubCellInst2_LFInst_14_LFInst_0_n8 ,
         \SubCellInst2_LFInst_14_LFInst_0_n7 ,
         \SubCellInst2_LFInst_14_LFInst_1_n6 ,
         \SubCellInst2_LFInst_14_LFInst_1_n5 ,
         \SubCellInst2_LFInst_14_LFInst_1_n4 ,
         \SubCellInst2_LFInst_14_LFInst_2_n11 ,
         \SubCellInst2_LFInst_14_LFInst_2_n10 ,
         \SubCellInst2_LFInst_14_LFInst_2_n9 ,
         \SubCellInst2_LFInst_14_LFInst_2_n8 ,
         \SubCellInst2_LFInst_14_LFInst_2_n7 ,
         \SubCellInst2_LFInst_14_LFInst_3_n6 ,
         \SubCellInst2_LFInst_14_LFInst_3_n5 ,
         \SubCellInst2_LFInst_14_LFInst_3_n4 ,
         \SubCellInst2_LFInst_15_LFInst_0_n11 ,
         \SubCellInst2_LFInst_15_LFInst_0_n10 ,
         \SubCellInst2_LFInst_15_LFInst_0_n9 ,
         \SubCellInst2_LFInst_15_LFInst_0_n8 ,
         \SubCellInst2_LFInst_15_LFInst_0_n7 ,
         \SubCellInst2_LFInst_15_LFInst_1_n6 ,
         \SubCellInst2_LFInst_15_LFInst_1_n5 ,
         \SubCellInst2_LFInst_15_LFInst_1_n4 ,
         \SubCellInst2_LFInst_15_LFInst_2_n11 ,
         \SubCellInst2_LFInst_15_LFInst_2_n10 ,
         \SubCellInst2_LFInst_15_LFInst_2_n9 ,
         \SubCellInst2_LFInst_15_LFInst_2_n8 ,
         \SubCellInst2_LFInst_15_LFInst_2_n7 ,
         \SubCellInst2_LFInst_15_LFInst_3_n6 ,
         \SubCellInst2_LFInst_15_LFInst_3_n5 ,
         \SubCellInst2_LFInst_15_LFInst_3_n4 , \MCInst3_XOR_r0_Inst_0_n3 ,
         \MCInst3_XOR_r0_Inst_1_n3 , \MCInst3_XOR_r0_Inst_2_n3 ,
         \MCInst3_XOR_r0_Inst_3_n3 , \MCInst3_XOR_r0_Inst_4_n3 ,
         \MCInst3_XOR_r0_Inst_5_n3 , \MCInst3_XOR_r0_Inst_6_n3 ,
         \MCInst3_XOR_r0_Inst_7_n3 , \MCInst3_XOR_r0_Inst_8_n3 ,
         \MCInst3_XOR_r0_Inst_9_n3 , \MCInst3_XOR_r0_Inst_10_n3 ,
         \MCInst3_XOR_r0_Inst_11_n3 , \MCInst3_XOR_r0_Inst_12_n3 ,
         \MCInst3_XOR_r0_Inst_13_n3 , \MCInst3_XOR_r0_Inst_14_n3 ,
         \MCInst3_XOR_r0_Inst_15_n3 , \SubCellInst3_LFInst_0_LFInst_0_n11 ,
         \SubCellInst3_LFInst_0_LFInst_0_n10 ,
         \SubCellInst3_LFInst_0_LFInst_0_n9 ,
         \SubCellInst3_LFInst_0_LFInst_0_n8 ,
         \SubCellInst3_LFInst_0_LFInst_0_n7 ,
         \SubCellInst3_LFInst_0_LFInst_1_n6 ,
         \SubCellInst3_LFInst_0_LFInst_1_n5 ,
         \SubCellInst3_LFInst_0_LFInst_1_n4 ,
         \SubCellInst3_LFInst_0_LFInst_2_n11 ,
         \SubCellInst3_LFInst_0_LFInst_2_n10 ,
         \SubCellInst3_LFInst_0_LFInst_2_n9 ,
         \SubCellInst3_LFInst_0_LFInst_2_n8 ,
         \SubCellInst3_LFInst_0_LFInst_2_n7 ,
         \SubCellInst3_LFInst_0_LFInst_3_n6 ,
         \SubCellInst3_LFInst_0_LFInst_3_n5 ,
         \SubCellInst3_LFInst_0_LFInst_3_n4 ,
         \SubCellInst3_LFInst_1_LFInst_0_n11 ,
         \SubCellInst3_LFInst_1_LFInst_0_n10 ,
         \SubCellInst3_LFInst_1_LFInst_0_n9 ,
         \SubCellInst3_LFInst_1_LFInst_0_n8 ,
         \SubCellInst3_LFInst_1_LFInst_0_n7 ,
         \SubCellInst3_LFInst_1_LFInst_1_n6 ,
         \SubCellInst3_LFInst_1_LFInst_1_n5 ,
         \SubCellInst3_LFInst_1_LFInst_1_n4 ,
         \SubCellInst3_LFInst_1_LFInst_2_n11 ,
         \SubCellInst3_LFInst_1_LFInst_2_n10 ,
         \SubCellInst3_LFInst_1_LFInst_2_n9 ,
         \SubCellInst3_LFInst_1_LFInst_2_n8 ,
         \SubCellInst3_LFInst_1_LFInst_2_n7 ,
         \SubCellInst3_LFInst_1_LFInst_3_n6 ,
         \SubCellInst3_LFInst_1_LFInst_3_n5 ,
         \SubCellInst3_LFInst_1_LFInst_3_n4 ,
         \SubCellInst3_LFInst_2_LFInst_0_n11 ,
         \SubCellInst3_LFInst_2_LFInst_0_n10 ,
         \SubCellInst3_LFInst_2_LFInst_0_n9 ,
         \SubCellInst3_LFInst_2_LFInst_0_n8 ,
         \SubCellInst3_LFInst_2_LFInst_0_n7 ,
         \SubCellInst3_LFInst_2_LFInst_1_n6 ,
         \SubCellInst3_LFInst_2_LFInst_1_n5 ,
         \SubCellInst3_LFInst_2_LFInst_1_n4 ,
         \SubCellInst3_LFInst_2_LFInst_2_n11 ,
         \SubCellInst3_LFInst_2_LFInst_2_n10 ,
         \SubCellInst3_LFInst_2_LFInst_2_n9 ,
         \SubCellInst3_LFInst_2_LFInst_2_n8 ,
         \SubCellInst3_LFInst_2_LFInst_2_n7 ,
         \SubCellInst3_LFInst_2_LFInst_3_n6 ,
         \SubCellInst3_LFInst_2_LFInst_3_n5 ,
         \SubCellInst3_LFInst_2_LFInst_3_n4 ,
         \SubCellInst3_LFInst_3_LFInst_0_n11 ,
         \SubCellInst3_LFInst_3_LFInst_0_n10 ,
         \SubCellInst3_LFInst_3_LFInst_0_n9 ,
         \SubCellInst3_LFInst_3_LFInst_0_n8 ,
         \SubCellInst3_LFInst_3_LFInst_0_n7 ,
         \SubCellInst3_LFInst_3_LFInst_1_n6 ,
         \SubCellInst3_LFInst_3_LFInst_1_n5 ,
         \SubCellInst3_LFInst_3_LFInst_1_n4 ,
         \SubCellInst3_LFInst_3_LFInst_2_n11 ,
         \SubCellInst3_LFInst_3_LFInst_2_n10 ,
         \SubCellInst3_LFInst_3_LFInst_2_n9 ,
         \SubCellInst3_LFInst_3_LFInst_2_n8 ,
         \SubCellInst3_LFInst_3_LFInst_2_n7 ,
         \SubCellInst3_LFInst_3_LFInst_3_n6 ,
         \SubCellInst3_LFInst_3_LFInst_3_n5 ,
         \SubCellInst3_LFInst_3_LFInst_3_n4 ,
         \SubCellInst3_LFInst_4_LFInst_0_n11 ,
         \SubCellInst3_LFInst_4_LFInst_0_n10 ,
         \SubCellInst3_LFInst_4_LFInst_0_n9 ,
         \SubCellInst3_LFInst_4_LFInst_0_n8 ,
         \SubCellInst3_LFInst_4_LFInst_0_n7 ,
         \SubCellInst3_LFInst_4_LFInst_1_n6 ,
         \SubCellInst3_LFInst_4_LFInst_1_n5 ,
         \SubCellInst3_LFInst_4_LFInst_1_n4 ,
         \SubCellInst3_LFInst_4_LFInst_2_n11 ,
         \SubCellInst3_LFInst_4_LFInst_2_n10 ,
         \SubCellInst3_LFInst_4_LFInst_2_n9 ,
         \SubCellInst3_LFInst_4_LFInst_2_n8 ,
         \SubCellInst3_LFInst_4_LFInst_2_n7 ,
         \SubCellInst3_LFInst_4_LFInst_3_n6 ,
         \SubCellInst3_LFInst_4_LFInst_3_n5 ,
         \SubCellInst3_LFInst_4_LFInst_3_n4 ,
         \SubCellInst3_LFInst_5_LFInst_0_n11 ,
         \SubCellInst3_LFInst_5_LFInst_0_n10 ,
         \SubCellInst3_LFInst_5_LFInst_0_n9 ,
         \SubCellInst3_LFInst_5_LFInst_0_n8 ,
         \SubCellInst3_LFInst_5_LFInst_0_n7 ,
         \SubCellInst3_LFInst_5_LFInst_1_n6 ,
         \SubCellInst3_LFInst_5_LFInst_1_n5 ,
         \SubCellInst3_LFInst_5_LFInst_1_n4 ,
         \SubCellInst3_LFInst_5_LFInst_2_n11 ,
         \SubCellInst3_LFInst_5_LFInst_2_n10 ,
         \SubCellInst3_LFInst_5_LFInst_2_n9 ,
         \SubCellInst3_LFInst_5_LFInst_2_n8 ,
         \SubCellInst3_LFInst_5_LFInst_2_n7 ,
         \SubCellInst3_LFInst_5_LFInst_3_n6 ,
         \SubCellInst3_LFInst_5_LFInst_3_n5 ,
         \SubCellInst3_LFInst_5_LFInst_3_n4 ,
         \SubCellInst3_LFInst_6_LFInst_0_n11 ,
         \SubCellInst3_LFInst_6_LFInst_0_n10 ,
         \SubCellInst3_LFInst_6_LFInst_0_n9 ,
         \SubCellInst3_LFInst_6_LFInst_0_n8 ,
         \SubCellInst3_LFInst_6_LFInst_0_n7 ,
         \SubCellInst3_LFInst_6_LFInst_1_n6 ,
         \SubCellInst3_LFInst_6_LFInst_1_n5 ,
         \SubCellInst3_LFInst_6_LFInst_1_n4 ,
         \SubCellInst3_LFInst_6_LFInst_2_n11 ,
         \SubCellInst3_LFInst_6_LFInst_2_n10 ,
         \SubCellInst3_LFInst_6_LFInst_2_n9 ,
         \SubCellInst3_LFInst_6_LFInst_2_n8 ,
         \SubCellInst3_LFInst_6_LFInst_2_n7 ,
         \SubCellInst3_LFInst_6_LFInst_3_n6 ,
         \SubCellInst3_LFInst_6_LFInst_3_n5 ,
         \SubCellInst3_LFInst_6_LFInst_3_n4 ,
         \SubCellInst3_LFInst_7_LFInst_0_n11 ,
         \SubCellInst3_LFInst_7_LFInst_0_n10 ,
         \SubCellInst3_LFInst_7_LFInst_0_n9 ,
         \SubCellInst3_LFInst_7_LFInst_0_n8 ,
         \SubCellInst3_LFInst_7_LFInst_0_n7 ,
         \SubCellInst3_LFInst_7_LFInst_1_n6 ,
         \SubCellInst3_LFInst_7_LFInst_1_n5 ,
         \SubCellInst3_LFInst_7_LFInst_1_n4 ,
         \SubCellInst3_LFInst_7_LFInst_2_n11 ,
         \SubCellInst3_LFInst_7_LFInst_2_n10 ,
         \SubCellInst3_LFInst_7_LFInst_2_n9 ,
         \SubCellInst3_LFInst_7_LFInst_2_n8 ,
         \SubCellInst3_LFInst_7_LFInst_2_n7 ,
         \SubCellInst3_LFInst_7_LFInst_3_n6 ,
         \SubCellInst3_LFInst_7_LFInst_3_n5 ,
         \SubCellInst3_LFInst_7_LFInst_3_n4 ,
         \SubCellInst3_LFInst_8_LFInst_0_n11 ,
         \SubCellInst3_LFInst_8_LFInst_0_n10 ,
         \SubCellInst3_LFInst_8_LFInst_0_n9 ,
         \SubCellInst3_LFInst_8_LFInst_0_n8 ,
         \SubCellInst3_LFInst_8_LFInst_0_n7 ,
         \SubCellInst3_LFInst_8_LFInst_1_n6 ,
         \SubCellInst3_LFInst_8_LFInst_1_n5 ,
         \SubCellInst3_LFInst_8_LFInst_1_n4 ,
         \SubCellInst3_LFInst_8_LFInst_2_n11 ,
         \SubCellInst3_LFInst_8_LFInst_2_n10 ,
         \SubCellInst3_LFInst_8_LFInst_2_n9 ,
         \SubCellInst3_LFInst_8_LFInst_2_n8 ,
         \SubCellInst3_LFInst_8_LFInst_2_n7 ,
         \SubCellInst3_LFInst_8_LFInst_3_n6 ,
         \SubCellInst3_LFInst_8_LFInst_3_n5 ,
         \SubCellInst3_LFInst_8_LFInst_3_n4 ,
         \SubCellInst3_LFInst_9_LFInst_0_n11 ,
         \SubCellInst3_LFInst_9_LFInst_0_n10 ,
         \SubCellInst3_LFInst_9_LFInst_0_n9 ,
         \SubCellInst3_LFInst_9_LFInst_0_n8 ,
         \SubCellInst3_LFInst_9_LFInst_0_n7 ,
         \SubCellInst3_LFInst_9_LFInst_1_n6 ,
         \SubCellInst3_LFInst_9_LFInst_1_n5 ,
         \SubCellInst3_LFInst_9_LFInst_1_n4 ,
         \SubCellInst3_LFInst_9_LFInst_2_n11 ,
         \SubCellInst3_LFInst_9_LFInst_2_n10 ,
         \SubCellInst3_LFInst_9_LFInst_2_n9 ,
         \SubCellInst3_LFInst_9_LFInst_2_n8 ,
         \SubCellInst3_LFInst_9_LFInst_2_n7 ,
         \SubCellInst3_LFInst_9_LFInst_3_n6 ,
         \SubCellInst3_LFInst_9_LFInst_3_n5 ,
         \SubCellInst3_LFInst_9_LFInst_3_n4 ,
         \SubCellInst3_LFInst_10_LFInst_0_n11 ,
         \SubCellInst3_LFInst_10_LFInst_0_n10 ,
         \SubCellInst3_LFInst_10_LFInst_0_n9 ,
         \SubCellInst3_LFInst_10_LFInst_0_n8 ,
         \SubCellInst3_LFInst_10_LFInst_0_n7 ,
         \SubCellInst3_LFInst_10_LFInst_1_n6 ,
         \SubCellInst3_LFInst_10_LFInst_1_n5 ,
         \SubCellInst3_LFInst_10_LFInst_1_n4 ,
         \SubCellInst3_LFInst_10_LFInst_2_n11 ,
         \SubCellInst3_LFInst_10_LFInst_2_n10 ,
         \SubCellInst3_LFInst_10_LFInst_2_n9 ,
         \SubCellInst3_LFInst_10_LFInst_2_n8 ,
         \SubCellInst3_LFInst_10_LFInst_2_n7 ,
         \SubCellInst3_LFInst_10_LFInst_3_n6 ,
         \SubCellInst3_LFInst_10_LFInst_3_n5 ,
         \SubCellInst3_LFInst_10_LFInst_3_n4 ,
         \SubCellInst3_LFInst_11_LFInst_0_n11 ,
         \SubCellInst3_LFInst_11_LFInst_0_n10 ,
         \SubCellInst3_LFInst_11_LFInst_0_n9 ,
         \SubCellInst3_LFInst_11_LFInst_0_n8 ,
         \SubCellInst3_LFInst_11_LFInst_0_n7 ,
         \SubCellInst3_LFInst_11_LFInst_1_n6 ,
         \SubCellInst3_LFInst_11_LFInst_1_n5 ,
         \SubCellInst3_LFInst_11_LFInst_1_n4 ,
         \SubCellInst3_LFInst_11_LFInst_2_n11 ,
         \SubCellInst3_LFInst_11_LFInst_2_n10 ,
         \SubCellInst3_LFInst_11_LFInst_2_n9 ,
         \SubCellInst3_LFInst_11_LFInst_2_n8 ,
         \SubCellInst3_LFInst_11_LFInst_2_n7 ,
         \SubCellInst3_LFInst_11_LFInst_3_n6 ,
         \SubCellInst3_LFInst_11_LFInst_3_n5 ,
         \SubCellInst3_LFInst_11_LFInst_3_n4 ,
         \SubCellInst3_LFInst_12_LFInst_0_n11 ,
         \SubCellInst3_LFInst_12_LFInst_0_n10 ,
         \SubCellInst3_LFInst_12_LFInst_0_n9 ,
         \SubCellInst3_LFInst_12_LFInst_0_n8 ,
         \SubCellInst3_LFInst_12_LFInst_0_n7 ,
         \SubCellInst3_LFInst_12_LFInst_1_n6 ,
         \SubCellInst3_LFInst_12_LFInst_1_n5 ,
         \SubCellInst3_LFInst_12_LFInst_1_n4 ,
         \SubCellInst3_LFInst_12_LFInst_2_n11 ,
         \SubCellInst3_LFInst_12_LFInst_2_n10 ,
         \SubCellInst3_LFInst_12_LFInst_2_n9 ,
         \SubCellInst3_LFInst_12_LFInst_2_n8 ,
         \SubCellInst3_LFInst_12_LFInst_2_n7 ,
         \SubCellInst3_LFInst_12_LFInst_3_n6 ,
         \SubCellInst3_LFInst_12_LFInst_3_n5 ,
         \SubCellInst3_LFInst_12_LFInst_3_n4 ,
         \SubCellInst3_LFInst_13_LFInst_0_n11 ,
         \SubCellInst3_LFInst_13_LFInst_0_n10 ,
         \SubCellInst3_LFInst_13_LFInst_0_n9 ,
         \SubCellInst3_LFInst_13_LFInst_0_n8 ,
         \SubCellInst3_LFInst_13_LFInst_0_n7 ,
         \SubCellInst3_LFInst_13_LFInst_1_n6 ,
         \SubCellInst3_LFInst_13_LFInst_1_n5 ,
         \SubCellInst3_LFInst_13_LFInst_1_n4 ,
         \SubCellInst3_LFInst_13_LFInst_2_n11 ,
         \SubCellInst3_LFInst_13_LFInst_2_n10 ,
         \SubCellInst3_LFInst_13_LFInst_2_n9 ,
         \SubCellInst3_LFInst_13_LFInst_2_n8 ,
         \SubCellInst3_LFInst_13_LFInst_2_n7 ,
         \SubCellInst3_LFInst_13_LFInst_3_n6 ,
         \SubCellInst3_LFInst_13_LFInst_3_n5 ,
         \SubCellInst3_LFInst_13_LFInst_3_n4 ,
         \SubCellInst3_LFInst_14_LFInst_0_n11 ,
         \SubCellInst3_LFInst_14_LFInst_0_n10 ,
         \SubCellInst3_LFInst_14_LFInst_0_n9 ,
         \SubCellInst3_LFInst_14_LFInst_0_n8 ,
         \SubCellInst3_LFInst_14_LFInst_0_n7 ,
         \SubCellInst3_LFInst_14_LFInst_1_n6 ,
         \SubCellInst3_LFInst_14_LFInst_1_n5 ,
         \SubCellInst3_LFInst_14_LFInst_1_n4 ,
         \SubCellInst3_LFInst_14_LFInst_2_n11 ,
         \SubCellInst3_LFInst_14_LFInst_2_n10 ,
         \SubCellInst3_LFInst_14_LFInst_2_n9 ,
         \SubCellInst3_LFInst_14_LFInst_2_n8 ,
         \SubCellInst3_LFInst_14_LFInst_2_n7 ,
         \SubCellInst3_LFInst_14_LFInst_3_n6 ,
         \SubCellInst3_LFInst_14_LFInst_3_n5 ,
         \SubCellInst3_LFInst_14_LFInst_3_n4 ,
         \SubCellInst3_LFInst_15_LFInst_0_n11 ,
         \SubCellInst3_LFInst_15_LFInst_0_n10 ,
         \SubCellInst3_LFInst_15_LFInst_0_n9 ,
         \SubCellInst3_LFInst_15_LFInst_0_n8 ,
         \SubCellInst3_LFInst_15_LFInst_0_n7 ,
         \SubCellInst3_LFInst_15_LFInst_1_n6 ,
         \SubCellInst3_LFInst_15_LFInst_1_n5 ,
         \SubCellInst3_LFInst_15_LFInst_1_n4 ,
         \SubCellInst3_LFInst_15_LFInst_2_n11 ,
         \SubCellInst3_LFInst_15_LFInst_2_n10 ,
         \SubCellInst3_LFInst_15_LFInst_2_n9 ,
         \SubCellInst3_LFInst_15_LFInst_2_n8 ,
         \SubCellInst3_LFInst_15_LFInst_2_n7 ,
         \SubCellInst3_LFInst_15_LFInst_3_n6 ,
         \SubCellInst3_LFInst_15_LFInst_3_n5 ,
         \SubCellInst3_LFInst_15_LFInst_3_n4 ,
         \Red_PlaintextInst_LFInst_0_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_0_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_0_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_0_LFInst_3_n2 ,
         \Red_PlaintextInst_LFInst_1_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_1_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_1_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_1_LFInst_3_n2 ,
         \Red_PlaintextInst_LFInst_2_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_2_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_2_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_2_LFInst_3_n2 ,
         \Red_PlaintextInst_LFInst_3_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_3_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_3_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_3_LFInst_3_n2 ,
         \Red_PlaintextInst_LFInst_4_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_4_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_4_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_4_LFInst_3_n2 ,
         \Red_PlaintextInst_LFInst_5_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_5_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_5_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_5_LFInst_3_n2 ,
         \Red_PlaintextInst_LFInst_6_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_6_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_6_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_6_LFInst_3_n2 ,
         \Red_PlaintextInst_LFInst_7_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_7_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_7_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_7_LFInst_3_n2 ,
         \Red_PlaintextInst_LFInst_8_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_8_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_8_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_8_LFInst_3_n2 ,
         \Red_PlaintextInst_LFInst_9_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_9_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_9_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_9_LFInst_3_n2 ,
         \Red_PlaintextInst_LFInst_10_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_10_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_10_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_10_LFInst_3_n2 ,
         \Red_PlaintextInst_LFInst_11_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_11_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_11_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_11_LFInst_3_n2 ,
         \Red_PlaintextInst_LFInst_12_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_12_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_12_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_12_LFInst_3_n2 ,
         \Red_PlaintextInst_LFInst_13_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_13_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_13_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_13_LFInst_3_n2 ,
         \Red_PlaintextInst_LFInst_14_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_14_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_14_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_14_LFInst_3_n2 ,
         \Red_PlaintextInst_LFInst_15_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_15_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_15_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_15_LFInst_3_n2 ,
         \Red_MCInst_XOR_r0_Inst_0_n3 , \Red_MCInst_XOR_r0_Inst_1_n3 ,
         \Red_MCInst_XOR_r0_Inst_2_n3 , \Red_MCInst_XOR_r0_Inst_3_n3 ,
         \Red_MCInst_XOR_r0_Inst_4_n3 , \Red_MCInst_XOR_r0_Inst_5_n3 ,
         \Red_MCInst_XOR_r0_Inst_6_n3 , \Red_MCInst_XOR_r0_Inst_7_n3 ,
         \Red_MCInst_XOR_r0_Inst_8_n3 , \Red_MCInst_XOR_r0_Inst_9_n3 ,
         \Red_MCInst_XOR_r0_Inst_10_n3 , \Red_MCInst_XOR_r0_Inst_11_n3 ,
         \Red_MCInst_XOR_r0_Inst_12_n3 , \Red_MCInst_XOR_r0_Inst_13_n3 ,
         \Red_MCInst_XOR_r0_Inst_14_n3 , \Red_MCInst_XOR_r0_Inst_15_n3 ,
         \Red_SubCellInst_LFInst_0_LFInst_0_n14 ,
         \Red_SubCellInst_LFInst_0_LFInst_0_n13 ,
         \Red_SubCellInst_LFInst_0_LFInst_0_n12 ,
         \Red_SubCellInst_LFInst_0_LFInst_0_n11 ,
         \Red_SubCellInst_LFInst_0_LFInst_0_n10 ,
         \Red_SubCellInst_LFInst_0_LFInst_0_n9 ,
         \Red_SubCellInst_LFInst_0_LFInst_0_n8 ,
         \Red_SubCellInst_LFInst_0_LFInst_1_n15 ,
         \Red_SubCellInst_LFInst_0_LFInst_1_n14 ,
         \Red_SubCellInst_LFInst_0_LFInst_1_n13 ,
         \Red_SubCellInst_LFInst_0_LFInst_1_n12 ,
         \Red_SubCellInst_LFInst_0_LFInst_1_n11 ,
         \Red_SubCellInst_LFInst_0_LFInst_2_n19 ,
         \Red_SubCellInst_LFInst_0_LFInst_2_n18 ,
         \Red_SubCellInst_LFInst_0_LFInst_2_n17 ,
         \Red_SubCellInst_LFInst_0_LFInst_2_n16 ,
         \Red_SubCellInst_LFInst_0_LFInst_2_n15 ,
         \Red_SubCellInst_LFInst_0_LFInst_2_n14 ,
         \Red_SubCellInst_LFInst_0_LFInst_2_n13 ,
         \Red_SubCellInst_LFInst_0_LFInst_3_n8 ,
         \Red_SubCellInst_LFInst_0_LFInst_3_n7 ,
         \Red_SubCellInst_LFInst_0_LFInst_3_n6 ,
         \Red_SubCellInst_LFInst_1_LFInst_0_n14 ,
         \Red_SubCellInst_LFInst_1_LFInst_0_n13 ,
         \Red_SubCellInst_LFInst_1_LFInst_0_n12 ,
         \Red_SubCellInst_LFInst_1_LFInst_0_n11 ,
         \Red_SubCellInst_LFInst_1_LFInst_0_n10 ,
         \Red_SubCellInst_LFInst_1_LFInst_0_n9 ,
         \Red_SubCellInst_LFInst_1_LFInst_0_n8 ,
         \Red_SubCellInst_LFInst_1_LFInst_1_n15 ,
         \Red_SubCellInst_LFInst_1_LFInst_1_n14 ,
         \Red_SubCellInst_LFInst_1_LFInst_1_n13 ,
         \Red_SubCellInst_LFInst_1_LFInst_1_n12 ,
         \Red_SubCellInst_LFInst_1_LFInst_1_n11 ,
         \Red_SubCellInst_LFInst_1_LFInst_2_n19 ,
         \Red_SubCellInst_LFInst_1_LFInst_2_n18 ,
         \Red_SubCellInst_LFInst_1_LFInst_2_n17 ,
         \Red_SubCellInst_LFInst_1_LFInst_2_n16 ,
         \Red_SubCellInst_LFInst_1_LFInst_2_n15 ,
         \Red_SubCellInst_LFInst_1_LFInst_2_n14 ,
         \Red_SubCellInst_LFInst_1_LFInst_2_n13 ,
         \Red_SubCellInst_LFInst_1_LFInst_3_n8 ,
         \Red_SubCellInst_LFInst_1_LFInst_3_n7 ,
         \Red_SubCellInst_LFInst_1_LFInst_3_n6 ,
         \Red_SubCellInst_LFInst_2_LFInst_0_n14 ,
         \Red_SubCellInst_LFInst_2_LFInst_0_n13 ,
         \Red_SubCellInst_LFInst_2_LFInst_0_n12 ,
         \Red_SubCellInst_LFInst_2_LFInst_0_n11 ,
         \Red_SubCellInst_LFInst_2_LFInst_0_n10 ,
         \Red_SubCellInst_LFInst_2_LFInst_0_n9 ,
         \Red_SubCellInst_LFInst_2_LFInst_0_n8 ,
         \Red_SubCellInst_LFInst_2_LFInst_1_n15 ,
         \Red_SubCellInst_LFInst_2_LFInst_1_n14 ,
         \Red_SubCellInst_LFInst_2_LFInst_1_n13 ,
         \Red_SubCellInst_LFInst_2_LFInst_1_n12 ,
         \Red_SubCellInst_LFInst_2_LFInst_1_n11 ,
         \Red_SubCellInst_LFInst_2_LFInst_2_n19 ,
         \Red_SubCellInst_LFInst_2_LFInst_2_n18 ,
         \Red_SubCellInst_LFInst_2_LFInst_2_n17 ,
         \Red_SubCellInst_LFInst_2_LFInst_2_n16 ,
         \Red_SubCellInst_LFInst_2_LFInst_2_n15 ,
         \Red_SubCellInst_LFInst_2_LFInst_2_n14 ,
         \Red_SubCellInst_LFInst_2_LFInst_2_n13 ,
         \Red_SubCellInst_LFInst_2_LFInst_3_n8 ,
         \Red_SubCellInst_LFInst_2_LFInst_3_n7 ,
         \Red_SubCellInst_LFInst_2_LFInst_3_n6 ,
         \Red_SubCellInst_LFInst_3_LFInst_0_n14 ,
         \Red_SubCellInst_LFInst_3_LFInst_0_n13 ,
         \Red_SubCellInst_LFInst_3_LFInst_0_n12 ,
         \Red_SubCellInst_LFInst_3_LFInst_0_n11 ,
         \Red_SubCellInst_LFInst_3_LFInst_0_n10 ,
         \Red_SubCellInst_LFInst_3_LFInst_0_n9 ,
         \Red_SubCellInst_LFInst_3_LFInst_0_n8 ,
         \Red_SubCellInst_LFInst_3_LFInst_1_n15 ,
         \Red_SubCellInst_LFInst_3_LFInst_1_n14 ,
         \Red_SubCellInst_LFInst_3_LFInst_1_n13 ,
         \Red_SubCellInst_LFInst_3_LFInst_1_n12 ,
         \Red_SubCellInst_LFInst_3_LFInst_1_n11 ,
         \Red_SubCellInst_LFInst_3_LFInst_2_n19 ,
         \Red_SubCellInst_LFInst_3_LFInst_2_n18 ,
         \Red_SubCellInst_LFInst_3_LFInst_2_n17 ,
         \Red_SubCellInst_LFInst_3_LFInst_2_n16 ,
         \Red_SubCellInst_LFInst_3_LFInst_2_n15 ,
         \Red_SubCellInst_LFInst_3_LFInst_2_n14 ,
         \Red_SubCellInst_LFInst_3_LFInst_2_n13 ,
         \Red_SubCellInst_LFInst_3_LFInst_3_n8 ,
         \Red_SubCellInst_LFInst_3_LFInst_3_n7 ,
         \Red_SubCellInst_LFInst_3_LFInst_3_n6 ,
         \Red_SubCellInst_LFInst_4_LFInst_0_n14 ,
         \Red_SubCellInst_LFInst_4_LFInst_0_n13 ,
         \Red_SubCellInst_LFInst_4_LFInst_0_n12 ,
         \Red_SubCellInst_LFInst_4_LFInst_0_n11 ,
         \Red_SubCellInst_LFInst_4_LFInst_0_n10 ,
         \Red_SubCellInst_LFInst_4_LFInst_0_n9 ,
         \Red_SubCellInst_LFInst_4_LFInst_0_n8 ,
         \Red_SubCellInst_LFInst_4_LFInst_1_n15 ,
         \Red_SubCellInst_LFInst_4_LFInst_1_n14 ,
         \Red_SubCellInst_LFInst_4_LFInst_1_n13 ,
         \Red_SubCellInst_LFInst_4_LFInst_1_n12 ,
         \Red_SubCellInst_LFInst_4_LFInst_1_n11 ,
         \Red_SubCellInst_LFInst_4_LFInst_2_n19 ,
         \Red_SubCellInst_LFInst_4_LFInst_2_n18 ,
         \Red_SubCellInst_LFInst_4_LFInst_2_n17 ,
         \Red_SubCellInst_LFInst_4_LFInst_2_n16 ,
         \Red_SubCellInst_LFInst_4_LFInst_2_n15 ,
         \Red_SubCellInst_LFInst_4_LFInst_2_n14 ,
         \Red_SubCellInst_LFInst_4_LFInst_2_n13 ,
         \Red_SubCellInst_LFInst_4_LFInst_3_n8 ,
         \Red_SubCellInst_LFInst_4_LFInst_3_n7 ,
         \Red_SubCellInst_LFInst_4_LFInst_3_n6 ,
         \Red_SubCellInst_LFInst_5_LFInst_0_n14 ,
         \Red_SubCellInst_LFInst_5_LFInst_0_n13 ,
         \Red_SubCellInst_LFInst_5_LFInst_0_n12 ,
         \Red_SubCellInst_LFInst_5_LFInst_0_n11 ,
         \Red_SubCellInst_LFInst_5_LFInst_0_n10 ,
         \Red_SubCellInst_LFInst_5_LFInst_0_n9 ,
         \Red_SubCellInst_LFInst_5_LFInst_0_n8 ,
         \Red_SubCellInst_LFInst_5_LFInst_1_n15 ,
         \Red_SubCellInst_LFInst_5_LFInst_1_n14 ,
         \Red_SubCellInst_LFInst_5_LFInst_1_n13 ,
         \Red_SubCellInst_LFInst_5_LFInst_1_n12 ,
         \Red_SubCellInst_LFInst_5_LFInst_1_n11 ,
         \Red_SubCellInst_LFInst_5_LFInst_2_n19 ,
         \Red_SubCellInst_LFInst_5_LFInst_2_n18 ,
         \Red_SubCellInst_LFInst_5_LFInst_2_n17 ,
         \Red_SubCellInst_LFInst_5_LFInst_2_n16 ,
         \Red_SubCellInst_LFInst_5_LFInst_2_n15 ,
         \Red_SubCellInst_LFInst_5_LFInst_2_n14 ,
         \Red_SubCellInst_LFInst_5_LFInst_2_n13 ,
         \Red_SubCellInst_LFInst_5_LFInst_3_n8 ,
         \Red_SubCellInst_LFInst_5_LFInst_3_n7 ,
         \Red_SubCellInst_LFInst_5_LFInst_3_n6 ,
         \Red_SubCellInst_LFInst_6_LFInst_0_n14 ,
         \Red_SubCellInst_LFInst_6_LFInst_0_n13 ,
         \Red_SubCellInst_LFInst_6_LFInst_0_n12 ,
         \Red_SubCellInst_LFInst_6_LFInst_0_n11 ,
         \Red_SubCellInst_LFInst_6_LFInst_0_n10 ,
         \Red_SubCellInst_LFInst_6_LFInst_0_n9 ,
         \Red_SubCellInst_LFInst_6_LFInst_0_n8 ,
         \Red_SubCellInst_LFInst_6_LFInst_1_n15 ,
         \Red_SubCellInst_LFInst_6_LFInst_1_n14 ,
         \Red_SubCellInst_LFInst_6_LFInst_1_n13 ,
         \Red_SubCellInst_LFInst_6_LFInst_1_n12 ,
         \Red_SubCellInst_LFInst_6_LFInst_1_n11 ,
         \Red_SubCellInst_LFInst_6_LFInst_2_n19 ,
         \Red_SubCellInst_LFInst_6_LFInst_2_n18 ,
         \Red_SubCellInst_LFInst_6_LFInst_2_n17 ,
         \Red_SubCellInst_LFInst_6_LFInst_2_n16 ,
         \Red_SubCellInst_LFInst_6_LFInst_2_n15 ,
         \Red_SubCellInst_LFInst_6_LFInst_2_n14 ,
         \Red_SubCellInst_LFInst_6_LFInst_2_n13 ,
         \Red_SubCellInst_LFInst_6_LFInst_3_n8 ,
         \Red_SubCellInst_LFInst_6_LFInst_3_n7 ,
         \Red_SubCellInst_LFInst_6_LFInst_3_n6 ,
         \Red_SubCellInst_LFInst_7_LFInst_0_n14 ,
         \Red_SubCellInst_LFInst_7_LFInst_0_n13 ,
         \Red_SubCellInst_LFInst_7_LFInst_0_n12 ,
         \Red_SubCellInst_LFInst_7_LFInst_0_n11 ,
         \Red_SubCellInst_LFInst_7_LFInst_0_n10 ,
         \Red_SubCellInst_LFInst_7_LFInst_0_n9 ,
         \Red_SubCellInst_LFInst_7_LFInst_0_n8 ,
         \Red_SubCellInst_LFInst_7_LFInst_1_n15 ,
         \Red_SubCellInst_LFInst_7_LFInst_1_n14 ,
         \Red_SubCellInst_LFInst_7_LFInst_1_n13 ,
         \Red_SubCellInst_LFInst_7_LFInst_1_n12 ,
         \Red_SubCellInst_LFInst_7_LFInst_1_n11 ,
         \Red_SubCellInst_LFInst_7_LFInst_2_n19 ,
         \Red_SubCellInst_LFInst_7_LFInst_2_n18 ,
         \Red_SubCellInst_LFInst_7_LFInst_2_n17 ,
         \Red_SubCellInst_LFInst_7_LFInst_2_n16 ,
         \Red_SubCellInst_LFInst_7_LFInst_2_n15 ,
         \Red_SubCellInst_LFInst_7_LFInst_2_n14 ,
         \Red_SubCellInst_LFInst_7_LFInst_2_n13 ,
         \Red_SubCellInst_LFInst_7_LFInst_3_n8 ,
         \Red_SubCellInst_LFInst_7_LFInst_3_n7 ,
         \Red_SubCellInst_LFInst_7_LFInst_3_n6 ,
         \Red_SubCellInst_LFInst_8_LFInst_0_n14 ,
         \Red_SubCellInst_LFInst_8_LFInst_0_n13 ,
         \Red_SubCellInst_LFInst_8_LFInst_0_n12 ,
         \Red_SubCellInst_LFInst_8_LFInst_0_n11 ,
         \Red_SubCellInst_LFInst_8_LFInst_0_n10 ,
         \Red_SubCellInst_LFInst_8_LFInst_0_n9 ,
         \Red_SubCellInst_LFInst_8_LFInst_0_n8 ,
         \Red_SubCellInst_LFInst_8_LFInst_1_n15 ,
         \Red_SubCellInst_LFInst_8_LFInst_1_n14 ,
         \Red_SubCellInst_LFInst_8_LFInst_1_n13 ,
         \Red_SubCellInst_LFInst_8_LFInst_1_n12 ,
         \Red_SubCellInst_LFInst_8_LFInst_1_n11 ,
         \Red_SubCellInst_LFInst_8_LFInst_2_n19 ,
         \Red_SubCellInst_LFInst_8_LFInst_2_n18 ,
         \Red_SubCellInst_LFInst_8_LFInst_2_n17 ,
         \Red_SubCellInst_LFInst_8_LFInst_2_n16 ,
         \Red_SubCellInst_LFInst_8_LFInst_2_n15 ,
         \Red_SubCellInst_LFInst_8_LFInst_2_n14 ,
         \Red_SubCellInst_LFInst_8_LFInst_2_n13 ,
         \Red_SubCellInst_LFInst_8_LFInst_3_n8 ,
         \Red_SubCellInst_LFInst_8_LFInst_3_n7 ,
         \Red_SubCellInst_LFInst_8_LFInst_3_n6 ,
         \Red_SubCellInst_LFInst_9_LFInst_0_n14 ,
         \Red_SubCellInst_LFInst_9_LFInst_0_n13 ,
         \Red_SubCellInst_LFInst_9_LFInst_0_n12 ,
         \Red_SubCellInst_LFInst_9_LFInst_0_n11 ,
         \Red_SubCellInst_LFInst_9_LFInst_0_n10 ,
         \Red_SubCellInst_LFInst_9_LFInst_0_n9 ,
         \Red_SubCellInst_LFInst_9_LFInst_0_n8 ,
         \Red_SubCellInst_LFInst_9_LFInst_1_n15 ,
         \Red_SubCellInst_LFInst_9_LFInst_1_n14 ,
         \Red_SubCellInst_LFInst_9_LFInst_1_n13 ,
         \Red_SubCellInst_LFInst_9_LFInst_1_n12 ,
         \Red_SubCellInst_LFInst_9_LFInst_1_n11 ,
         \Red_SubCellInst_LFInst_9_LFInst_2_n19 ,
         \Red_SubCellInst_LFInst_9_LFInst_2_n18 ,
         \Red_SubCellInst_LFInst_9_LFInst_2_n17 ,
         \Red_SubCellInst_LFInst_9_LFInst_2_n16 ,
         \Red_SubCellInst_LFInst_9_LFInst_2_n15 ,
         \Red_SubCellInst_LFInst_9_LFInst_2_n14 ,
         \Red_SubCellInst_LFInst_9_LFInst_2_n13 ,
         \Red_SubCellInst_LFInst_9_LFInst_3_n8 ,
         \Red_SubCellInst_LFInst_9_LFInst_3_n7 ,
         \Red_SubCellInst_LFInst_9_LFInst_3_n6 ,
         \Red_SubCellInst_LFInst_10_LFInst_0_n14 ,
         \Red_SubCellInst_LFInst_10_LFInst_0_n13 ,
         \Red_SubCellInst_LFInst_10_LFInst_0_n12 ,
         \Red_SubCellInst_LFInst_10_LFInst_0_n11 ,
         \Red_SubCellInst_LFInst_10_LFInst_0_n10 ,
         \Red_SubCellInst_LFInst_10_LFInst_0_n9 ,
         \Red_SubCellInst_LFInst_10_LFInst_0_n8 ,
         \Red_SubCellInst_LFInst_10_LFInst_1_n15 ,
         \Red_SubCellInst_LFInst_10_LFInst_1_n14 ,
         \Red_SubCellInst_LFInst_10_LFInst_1_n13 ,
         \Red_SubCellInst_LFInst_10_LFInst_1_n12 ,
         \Red_SubCellInst_LFInst_10_LFInst_1_n11 ,
         \Red_SubCellInst_LFInst_10_LFInst_2_n19 ,
         \Red_SubCellInst_LFInst_10_LFInst_2_n18 ,
         \Red_SubCellInst_LFInst_10_LFInst_2_n17 ,
         \Red_SubCellInst_LFInst_10_LFInst_2_n16 ,
         \Red_SubCellInst_LFInst_10_LFInst_2_n15 ,
         \Red_SubCellInst_LFInst_10_LFInst_2_n14 ,
         \Red_SubCellInst_LFInst_10_LFInst_2_n13 ,
         \Red_SubCellInst_LFInst_10_LFInst_3_n8 ,
         \Red_SubCellInst_LFInst_10_LFInst_3_n7 ,
         \Red_SubCellInst_LFInst_10_LFInst_3_n6 ,
         \Red_SubCellInst_LFInst_11_LFInst_0_n14 ,
         \Red_SubCellInst_LFInst_11_LFInst_0_n13 ,
         \Red_SubCellInst_LFInst_11_LFInst_0_n12 ,
         \Red_SubCellInst_LFInst_11_LFInst_0_n11 ,
         \Red_SubCellInst_LFInst_11_LFInst_0_n10 ,
         \Red_SubCellInst_LFInst_11_LFInst_0_n9 ,
         \Red_SubCellInst_LFInst_11_LFInst_0_n8 ,
         \Red_SubCellInst_LFInst_11_LFInst_1_n15 ,
         \Red_SubCellInst_LFInst_11_LFInst_1_n14 ,
         \Red_SubCellInst_LFInst_11_LFInst_1_n13 ,
         \Red_SubCellInst_LFInst_11_LFInst_1_n12 ,
         \Red_SubCellInst_LFInst_11_LFInst_1_n11 ,
         \Red_SubCellInst_LFInst_11_LFInst_2_n19 ,
         \Red_SubCellInst_LFInst_11_LFInst_2_n18 ,
         \Red_SubCellInst_LFInst_11_LFInst_2_n17 ,
         \Red_SubCellInst_LFInst_11_LFInst_2_n16 ,
         \Red_SubCellInst_LFInst_11_LFInst_2_n15 ,
         \Red_SubCellInst_LFInst_11_LFInst_2_n14 ,
         \Red_SubCellInst_LFInst_11_LFInst_2_n13 ,
         \Red_SubCellInst_LFInst_11_LFInst_3_n8 ,
         \Red_SubCellInst_LFInst_11_LFInst_3_n7 ,
         \Red_SubCellInst_LFInst_11_LFInst_3_n6 ,
         \Red_SubCellInst_LFInst_12_LFInst_0_n14 ,
         \Red_SubCellInst_LFInst_12_LFInst_0_n13 ,
         \Red_SubCellInst_LFInst_12_LFInst_0_n12 ,
         \Red_SubCellInst_LFInst_12_LFInst_0_n11 ,
         \Red_SubCellInst_LFInst_12_LFInst_0_n10 ,
         \Red_SubCellInst_LFInst_12_LFInst_0_n9 ,
         \Red_SubCellInst_LFInst_12_LFInst_0_n8 ,
         \Red_SubCellInst_LFInst_12_LFInst_1_n15 ,
         \Red_SubCellInst_LFInst_12_LFInst_1_n14 ,
         \Red_SubCellInst_LFInst_12_LFInst_1_n13 ,
         \Red_SubCellInst_LFInst_12_LFInst_1_n12 ,
         \Red_SubCellInst_LFInst_12_LFInst_1_n11 ,
         \Red_SubCellInst_LFInst_12_LFInst_2_n19 ,
         \Red_SubCellInst_LFInst_12_LFInst_2_n18 ,
         \Red_SubCellInst_LFInst_12_LFInst_2_n17 ,
         \Red_SubCellInst_LFInst_12_LFInst_2_n16 ,
         \Red_SubCellInst_LFInst_12_LFInst_2_n15 ,
         \Red_SubCellInst_LFInst_12_LFInst_2_n14 ,
         \Red_SubCellInst_LFInst_12_LFInst_2_n13 ,
         \Red_SubCellInst_LFInst_12_LFInst_3_n8 ,
         \Red_SubCellInst_LFInst_12_LFInst_3_n7 ,
         \Red_SubCellInst_LFInst_12_LFInst_3_n6 ,
         \Red_SubCellInst_LFInst_13_LFInst_0_n14 ,
         \Red_SubCellInst_LFInst_13_LFInst_0_n13 ,
         \Red_SubCellInst_LFInst_13_LFInst_0_n12 ,
         \Red_SubCellInst_LFInst_13_LFInst_0_n11 ,
         \Red_SubCellInst_LFInst_13_LFInst_0_n10 ,
         \Red_SubCellInst_LFInst_13_LFInst_0_n9 ,
         \Red_SubCellInst_LFInst_13_LFInst_0_n8 ,
         \Red_SubCellInst_LFInst_13_LFInst_1_n15 ,
         \Red_SubCellInst_LFInst_13_LFInst_1_n14 ,
         \Red_SubCellInst_LFInst_13_LFInst_1_n13 ,
         \Red_SubCellInst_LFInst_13_LFInst_1_n12 ,
         \Red_SubCellInst_LFInst_13_LFInst_1_n11 ,
         \Red_SubCellInst_LFInst_13_LFInst_2_n19 ,
         \Red_SubCellInst_LFInst_13_LFInst_2_n18 ,
         \Red_SubCellInst_LFInst_13_LFInst_2_n17 ,
         \Red_SubCellInst_LFInst_13_LFInst_2_n16 ,
         \Red_SubCellInst_LFInst_13_LFInst_2_n15 ,
         \Red_SubCellInst_LFInst_13_LFInst_2_n14 ,
         \Red_SubCellInst_LFInst_13_LFInst_2_n13 ,
         \Red_SubCellInst_LFInst_13_LFInst_3_n8 ,
         \Red_SubCellInst_LFInst_13_LFInst_3_n7 ,
         \Red_SubCellInst_LFInst_13_LFInst_3_n6 ,
         \Red_SubCellInst_LFInst_14_LFInst_0_n14 ,
         \Red_SubCellInst_LFInst_14_LFInst_0_n13 ,
         \Red_SubCellInst_LFInst_14_LFInst_0_n12 ,
         \Red_SubCellInst_LFInst_14_LFInst_0_n11 ,
         \Red_SubCellInst_LFInst_14_LFInst_0_n10 ,
         \Red_SubCellInst_LFInst_14_LFInst_0_n9 ,
         \Red_SubCellInst_LFInst_14_LFInst_0_n8 ,
         \Red_SubCellInst_LFInst_14_LFInst_1_n15 ,
         \Red_SubCellInst_LFInst_14_LFInst_1_n14 ,
         \Red_SubCellInst_LFInst_14_LFInst_1_n13 ,
         \Red_SubCellInst_LFInst_14_LFInst_1_n12 ,
         \Red_SubCellInst_LFInst_14_LFInst_1_n11 ,
         \Red_SubCellInst_LFInst_14_LFInst_2_n19 ,
         \Red_SubCellInst_LFInst_14_LFInst_2_n18 ,
         \Red_SubCellInst_LFInst_14_LFInst_2_n17 ,
         \Red_SubCellInst_LFInst_14_LFInst_2_n16 ,
         \Red_SubCellInst_LFInst_14_LFInst_2_n15 ,
         \Red_SubCellInst_LFInst_14_LFInst_2_n14 ,
         \Red_SubCellInst_LFInst_14_LFInst_2_n13 ,
         \Red_SubCellInst_LFInst_14_LFInst_3_n8 ,
         \Red_SubCellInst_LFInst_14_LFInst_3_n7 ,
         \Red_SubCellInst_LFInst_14_LFInst_3_n6 ,
         \Red_SubCellInst_LFInst_15_LFInst_0_n14 ,
         \Red_SubCellInst_LFInst_15_LFInst_0_n13 ,
         \Red_SubCellInst_LFInst_15_LFInst_0_n12 ,
         \Red_SubCellInst_LFInst_15_LFInst_0_n11 ,
         \Red_SubCellInst_LFInst_15_LFInst_0_n10 ,
         \Red_SubCellInst_LFInst_15_LFInst_0_n9 ,
         \Red_SubCellInst_LFInst_15_LFInst_0_n8 ,
         \Red_SubCellInst_LFInst_15_LFInst_1_n15 ,
         \Red_SubCellInst_LFInst_15_LFInst_1_n14 ,
         \Red_SubCellInst_LFInst_15_LFInst_1_n13 ,
         \Red_SubCellInst_LFInst_15_LFInst_1_n12 ,
         \Red_SubCellInst_LFInst_15_LFInst_1_n11 ,
         \Red_SubCellInst_LFInst_15_LFInst_2_n19 ,
         \Red_SubCellInst_LFInst_15_LFInst_2_n18 ,
         \Red_SubCellInst_LFInst_15_LFInst_2_n17 ,
         \Red_SubCellInst_LFInst_15_LFInst_2_n16 ,
         \Red_SubCellInst_LFInst_15_LFInst_2_n15 ,
         \Red_SubCellInst_LFInst_15_LFInst_2_n14 ,
         \Red_SubCellInst_LFInst_15_LFInst_2_n13 ,
         \Red_SubCellInst_LFInst_15_LFInst_3_n8 ,
         \Red_SubCellInst_LFInst_15_LFInst_3_n7 ,
         \Red_SubCellInst_LFInst_15_LFInst_3_n6 ,
         \Red_MCInst2_XOR_r0_Inst_0_n3 , \Red_MCInst2_XOR_r0_Inst_1_n3 ,
         \Red_MCInst2_XOR_r0_Inst_2_n3 , \Red_MCInst2_XOR_r0_Inst_3_n3 ,
         \Red_MCInst2_XOR_r0_Inst_4_n3 , \Red_MCInst2_XOR_r0_Inst_5_n3 ,
         \Red_MCInst2_XOR_r0_Inst_6_n3 , \Red_MCInst2_XOR_r0_Inst_7_n3 ,
         \Red_MCInst2_XOR_r0_Inst_8_n3 , \Red_MCInst2_XOR_r0_Inst_9_n3 ,
         \Red_MCInst2_XOR_r0_Inst_10_n3 , \Red_MCInst2_XOR_r0_Inst_11_n3 ,
         \Red_MCInst2_XOR_r0_Inst_12_n3 , \Red_MCInst2_XOR_r0_Inst_13_n3 ,
         \Red_MCInst2_XOR_r0_Inst_14_n3 , \Red_MCInst2_XOR_r0_Inst_15_n3 ,
         \Red_SubCellInst2_LFInst_0_LFInst_0_n14 ,
         \Red_SubCellInst2_LFInst_0_LFInst_0_n13 ,
         \Red_SubCellInst2_LFInst_0_LFInst_0_n12 ,
         \Red_SubCellInst2_LFInst_0_LFInst_0_n11 ,
         \Red_SubCellInst2_LFInst_0_LFInst_0_n10 ,
         \Red_SubCellInst2_LFInst_0_LFInst_0_n9 ,
         \Red_SubCellInst2_LFInst_0_LFInst_0_n8 ,
         \Red_SubCellInst2_LFInst_0_LFInst_1_n15 ,
         \Red_SubCellInst2_LFInst_0_LFInst_1_n14 ,
         \Red_SubCellInst2_LFInst_0_LFInst_1_n13 ,
         \Red_SubCellInst2_LFInst_0_LFInst_1_n12 ,
         \Red_SubCellInst2_LFInst_0_LFInst_1_n11 ,
         \Red_SubCellInst2_LFInst_0_LFInst_2_n19 ,
         \Red_SubCellInst2_LFInst_0_LFInst_2_n18 ,
         \Red_SubCellInst2_LFInst_0_LFInst_2_n17 ,
         \Red_SubCellInst2_LFInst_0_LFInst_2_n16 ,
         \Red_SubCellInst2_LFInst_0_LFInst_2_n15 ,
         \Red_SubCellInst2_LFInst_0_LFInst_2_n14 ,
         \Red_SubCellInst2_LFInst_0_LFInst_2_n13 ,
         \Red_SubCellInst2_LFInst_0_LFInst_3_n8 ,
         \Red_SubCellInst2_LFInst_0_LFInst_3_n7 ,
         \Red_SubCellInst2_LFInst_0_LFInst_3_n6 ,
         \Red_SubCellInst2_LFInst_1_LFInst_0_n14 ,
         \Red_SubCellInst2_LFInst_1_LFInst_0_n13 ,
         \Red_SubCellInst2_LFInst_1_LFInst_0_n12 ,
         \Red_SubCellInst2_LFInst_1_LFInst_0_n11 ,
         \Red_SubCellInst2_LFInst_1_LFInst_0_n10 ,
         \Red_SubCellInst2_LFInst_1_LFInst_0_n9 ,
         \Red_SubCellInst2_LFInst_1_LFInst_0_n8 ,
         \Red_SubCellInst2_LFInst_1_LFInst_1_n15 ,
         \Red_SubCellInst2_LFInst_1_LFInst_1_n14 ,
         \Red_SubCellInst2_LFInst_1_LFInst_1_n13 ,
         \Red_SubCellInst2_LFInst_1_LFInst_1_n12 ,
         \Red_SubCellInst2_LFInst_1_LFInst_1_n11 ,
         \Red_SubCellInst2_LFInst_1_LFInst_2_n19 ,
         \Red_SubCellInst2_LFInst_1_LFInst_2_n18 ,
         \Red_SubCellInst2_LFInst_1_LFInst_2_n17 ,
         \Red_SubCellInst2_LFInst_1_LFInst_2_n16 ,
         \Red_SubCellInst2_LFInst_1_LFInst_2_n15 ,
         \Red_SubCellInst2_LFInst_1_LFInst_2_n14 ,
         \Red_SubCellInst2_LFInst_1_LFInst_2_n13 ,
         \Red_SubCellInst2_LFInst_1_LFInst_3_n8 ,
         \Red_SubCellInst2_LFInst_1_LFInst_3_n7 ,
         \Red_SubCellInst2_LFInst_1_LFInst_3_n6 ,
         \Red_SubCellInst2_LFInst_2_LFInst_0_n14 ,
         \Red_SubCellInst2_LFInst_2_LFInst_0_n13 ,
         \Red_SubCellInst2_LFInst_2_LFInst_0_n12 ,
         \Red_SubCellInst2_LFInst_2_LFInst_0_n11 ,
         \Red_SubCellInst2_LFInst_2_LFInst_0_n10 ,
         \Red_SubCellInst2_LFInst_2_LFInst_0_n9 ,
         \Red_SubCellInst2_LFInst_2_LFInst_0_n8 ,
         \Red_SubCellInst2_LFInst_2_LFInst_1_n15 ,
         \Red_SubCellInst2_LFInst_2_LFInst_1_n14 ,
         \Red_SubCellInst2_LFInst_2_LFInst_1_n13 ,
         \Red_SubCellInst2_LFInst_2_LFInst_1_n12 ,
         \Red_SubCellInst2_LFInst_2_LFInst_1_n11 ,
         \Red_SubCellInst2_LFInst_2_LFInst_2_n19 ,
         \Red_SubCellInst2_LFInst_2_LFInst_2_n18 ,
         \Red_SubCellInst2_LFInst_2_LFInst_2_n17 ,
         \Red_SubCellInst2_LFInst_2_LFInst_2_n16 ,
         \Red_SubCellInst2_LFInst_2_LFInst_2_n15 ,
         \Red_SubCellInst2_LFInst_2_LFInst_2_n14 ,
         \Red_SubCellInst2_LFInst_2_LFInst_2_n13 ,
         \Red_SubCellInst2_LFInst_2_LFInst_3_n8 ,
         \Red_SubCellInst2_LFInst_2_LFInst_3_n7 ,
         \Red_SubCellInst2_LFInst_2_LFInst_3_n6 ,
         \Red_SubCellInst2_LFInst_3_LFInst_0_n14 ,
         \Red_SubCellInst2_LFInst_3_LFInst_0_n13 ,
         \Red_SubCellInst2_LFInst_3_LFInst_0_n12 ,
         \Red_SubCellInst2_LFInst_3_LFInst_0_n11 ,
         \Red_SubCellInst2_LFInst_3_LFInst_0_n10 ,
         \Red_SubCellInst2_LFInst_3_LFInst_0_n9 ,
         \Red_SubCellInst2_LFInst_3_LFInst_0_n8 ,
         \Red_SubCellInst2_LFInst_3_LFInst_1_n15 ,
         \Red_SubCellInst2_LFInst_3_LFInst_1_n14 ,
         \Red_SubCellInst2_LFInst_3_LFInst_1_n13 ,
         \Red_SubCellInst2_LFInst_3_LFInst_1_n12 ,
         \Red_SubCellInst2_LFInst_3_LFInst_1_n11 ,
         \Red_SubCellInst2_LFInst_3_LFInst_2_n19 ,
         \Red_SubCellInst2_LFInst_3_LFInst_2_n18 ,
         \Red_SubCellInst2_LFInst_3_LFInst_2_n17 ,
         \Red_SubCellInst2_LFInst_3_LFInst_2_n16 ,
         \Red_SubCellInst2_LFInst_3_LFInst_2_n15 ,
         \Red_SubCellInst2_LFInst_3_LFInst_2_n14 ,
         \Red_SubCellInst2_LFInst_3_LFInst_2_n13 ,
         \Red_SubCellInst2_LFInst_3_LFInst_3_n8 ,
         \Red_SubCellInst2_LFInst_3_LFInst_3_n7 ,
         \Red_SubCellInst2_LFInst_3_LFInst_3_n6 ,
         \Red_SubCellInst2_LFInst_4_LFInst_0_n14 ,
         \Red_SubCellInst2_LFInst_4_LFInst_0_n13 ,
         \Red_SubCellInst2_LFInst_4_LFInst_0_n12 ,
         \Red_SubCellInst2_LFInst_4_LFInst_0_n11 ,
         \Red_SubCellInst2_LFInst_4_LFInst_0_n10 ,
         \Red_SubCellInst2_LFInst_4_LFInst_0_n9 ,
         \Red_SubCellInst2_LFInst_4_LFInst_0_n8 ,
         \Red_SubCellInst2_LFInst_4_LFInst_1_n15 ,
         \Red_SubCellInst2_LFInst_4_LFInst_1_n14 ,
         \Red_SubCellInst2_LFInst_4_LFInst_1_n13 ,
         \Red_SubCellInst2_LFInst_4_LFInst_1_n12 ,
         \Red_SubCellInst2_LFInst_4_LFInst_1_n11 ,
         \Red_SubCellInst2_LFInst_4_LFInst_2_n19 ,
         \Red_SubCellInst2_LFInst_4_LFInst_2_n18 ,
         \Red_SubCellInst2_LFInst_4_LFInst_2_n17 ,
         \Red_SubCellInst2_LFInst_4_LFInst_2_n16 ,
         \Red_SubCellInst2_LFInst_4_LFInst_2_n15 ,
         \Red_SubCellInst2_LFInst_4_LFInst_2_n14 ,
         \Red_SubCellInst2_LFInst_4_LFInst_2_n13 ,
         \Red_SubCellInst2_LFInst_4_LFInst_3_n8 ,
         \Red_SubCellInst2_LFInst_4_LFInst_3_n7 ,
         \Red_SubCellInst2_LFInst_4_LFInst_3_n6 ,
         \Red_SubCellInst2_LFInst_5_LFInst_0_n14 ,
         \Red_SubCellInst2_LFInst_5_LFInst_0_n13 ,
         \Red_SubCellInst2_LFInst_5_LFInst_0_n12 ,
         \Red_SubCellInst2_LFInst_5_LFInst_0_n11 ,
         \Red_SubCellInst2_LFInst_5_LFInst_0_n10 ,
         \Red_SubCellInst2_LFInst_5_LFInst_0_n9 ,
         \Red_SubCellInst2_LFInst_5_LFInst_0_n8 ,
         \Red_SubCellInst2_LFInst_5_LFInst_1_n15 ,
         \Red_SubCellInst2_LFInst_5_LFInst_1_n14 ,
         \Red_SubCellInst2_LFInst_5_LFInst_1_n13 ,
         \Red_SubCellInst2_LFInst_5_LFInst_1_n12 ,
         \Red_SubCellInst2_LFInst_5_LFInst_1_n11 ,
         \Red_SubCellInst2_LFInst_5_LFInst_2_n19 ,
         \Red_SubCellInst2_LFInst_5_LFInst_2_n18 ,
         \Red_SubCellInst2_LFInst_5_LFInst_2_n17 ,
         \Red_SubCellInst2_LFInst_5_LFInst_2_n16 ,
         \Red_SubCellInst2_LFInst_5_LFInst_2_n15 ,
         \Red_SubCellInst2_LFInst_5_LFInst_2_n14 ,
         \Red_SubCellInst2_LFInst_5_LFInst_2_n13 ,
         \Red_SubCellInst2_LFInst_5_LFInst_3_n8 ,
         \Red_SubCellInst2_LFInst_5_LFInst_3_n7 ,
         \Red_SubCellInst2_LFInst_5_LFInst_3_n6 ,
         \Red_SubCellInst2_LFInst_6_LFInst_0_n14 ,
         \Red_SubCellInst2_LFInst_6_LFInst_0_n13 ,
         \Red_SubCellInst2_LFInst_6_LFInst_0_n12 ,
         \Red_SubCellInst2_LFInst_6_LFInst_0_n11 ,
         \Red_SubCellInst2_LFInst_6_LFInst_0_n10 ,
         \Red_SubCellInst2_LFInst_6_LFInst_0_n9 ,
         \Red_SubCellInst2_LFInst_6_LFInst_0_n8 ,
         \Red_SubCellInst2_LFInst_6_LFInst_1_n15 ,
         \Red_SubCellInst2_LFInst_6_LFInst_1_n14 ,
         \Red_SubCellInst2_LFInst_6_LFInst_1_n13 ,
         \Red_SubCellInst2_LFInst_6_LFInst_1_n12 ,
         \Red_SubCellInst2_LFInst_6_LFInst_1_n11 ,
         \Red_SubCellInst2_LFInst_6_LFInst_2_n19 ,
         \Red_SubCellInst2_LFInst_6_LFInst_2_n18 ,
         \Red_SubCellInst2_LFInst_6_LFInst_2_n17 ,
         \Red_SubCellInst2_LFInst_6_LFInst_2_n16 ,
         \Red_SubCellInst2_LFInst_6_LFInst_2_n15 ,
         \Red_SubCellInst2_LFInst_6_LFInst_2_n14 ,
         \Red_SubCellInst2_LFInst_6_LFInst_2_n13 ,
         \Red_SubCellInst2_LFInst_6_LFInst_3_n8 ,
         \Red_SubCellInst2_LFInst_6_LFInst_3_n7 ,
         \Red_SubCellInst2_LFInst_6_LFInst_3_n6 ,
         \Red_SubCellInst2_LFInst_7_LFInst_0_n14 ,
         \Red_SubCellInst2_LFInst_7_LFInst_0_n13 ,
         \Red_SubCellInst2_LFInst_7_LFInst_0_n12 ,
         \Red_SubCellInst2_LFInst_7_LFInst_0_n11 ,
         \Red_SubCellInst2_LFInst_7_LFInst_0_n10 ,
         \Red_SubCellInst2_LFInst_7_LFInst_0_n9 ,
         \Red_SubCellInst2_LFInst_7_LFInst_0_n8 ,
         \Red_SubCellInst2_LFInst_7_LFInst_1_n15 ,
         \Red_SubCellInst2_LFInst_7_LFInst_1_n14 ,
         \Red_SubCellInst2_LFInst_7_LFInst_1_n13 ,
         \Red_SubCellInst2_LFInst_7_LFInst_1_n12 ,
         \Red_SubCellInst2_LFInst_7_LFInst_1_n11 ,
         \Red_SubCellInst2_LFInst_7_LFInst_2_n19 ,
         \Red_SubCellInst2_LFInst_7_LFInst_2_n18 ,
         \Red_SubCellInst2_LFInst_7_LFInst_2_n17 ,
         \Red_SubCellInst2_LFInst_7_LFInst_2_n16 ,
         \Red_SubCellInst2_LFInst_7_LFInst_2_n15 ,
         \Red_SubCellInst2_LFInst_7_LFInst_2_n14 ,
         \Red_SubCellInst2_LFInst_7_LFInst_2_n13 ,
         \Red_SubCellInst2_LFInst_7_LFInst_3_n8 ,
         \Red_SubCellInst2_LFInst_7_LFInst_3_n7 ,
         \Red_SubCellInst2_LFInst_7_LFInst_3_n6 ,
         \Red_SubCellInst2_LFInst_8_LFInst_0_n14 ,
         \Red_SubCellInst2_LFInst_8_LFInst_0_n13 ,
         \Red_SubCellInst2_LFInst_8_LFInst_0_n12 ,
         \Red_SubCellInst2_LFInst_8_LFInst_0_n11 ,
         \Red_SubCellInst2_LFInst_8_LFInst_0_n10 ,
         \Red_SubCellInst2_LFInst_8_LFInst_0_n9 ,
         \Red_SubCellInst2_LFInst_8_LFInst_0_n8 ,
         \Red_SubCellInst2_LFInst_8_LFInst_1_n15 ,
         \Red_SubCellInst2_LFInst_8_LFInst_1_n14 ,
         \Red_SubCellInst2_LFInst_8_LFInst_1_n13 ,
         \Red_SubCellInst2_LFInst_8_LFInst_1_n12 ,
         \Red_SubCellInst2_LFInst_8_LFInst_1_n11 ,
         \Red_SubCellInst2_LFInst_8_LFInst_2_n19 ,
         \Red_SubCellInst2_LFInst_8_LFInst_2_n18 ,
         \Red_SubCellInst2_LFInst_8_LFInst_2_n17 ,
         \Red_SubCellInst2_LFInst_8_LFInst_2_n16 ,
         \Red_SubCellInst2_LFInst_8_LFInst_2_n15 ,
         \Red_SubCellInst2_LFInst_8_LFInst_2_n14 ,
         \Red_SubCellInst2_LFInst_8_LFInst_2_n13 ,
         \Red_SubCellInst2_LFInst_8_LFInst_3_n8 ,
         \Red_SubCellInst2_LFInst_8_LFInst_3_n7 ,
         \Red_SubCellInst2_LFInst_8_LFInst_3_n6 ,
         \Red_SubCellInst2_LFInst_9_LFInst_0_n14 ,
         \Red_SubCellInst2_LFInst_9_LFInst_0_n13 ,
         \Red_SubCellInst2_LFInst_9_LFInst_0_n12 ,
         \Red_SubCellInst2_LFInst_9_LFInst_0_n11 ,
         \Red_SubCellInst2_LFInst_9_LFInst_0_n10 ,
         \Red_SubCellInst2_LFInst_9_LFInst_0_n9 ,
         \Red_SubCellInst2_LFInst_9_LFInst_0_n8 ,
         \Red_SubCellInst2_LFInst_9_LFInst_1_n15 ,
         \Red_SubCellInst2_LFInst_9_LFInst_1_n14 ,
         \Red_SubCellInst2_LFInst_9_LFInst_1_n13 ,
         \Red_SubCellInst2_LFInst_9_LFInst_1_n12 ,
         \Red_SubCellInst2_LFInst_9_LFInst_1_n11 ,
         \Red_SubCellInst2_LFInst_9_LFInst_2_n19 ,
         \Red_SubCellInst2_LFInst_9_LFInst_2_n18 ,
         \Red_SubCellInst2_LFInst_9_LFInst_2_n17 ,
         \Red_SubCellInst2_LFInst_9_LFInst_2_n16 ,
         \Red_SubCellInst2_LFInst_9_LFInst_2_n15 ,
         \Red_SubCellInst2_LFInst_9_LFInst_2_n14 ,
         \Red_SubCellInst2_LFInst_9_LFInst_2_n13 ,
         \Red_SubCellInst2_LFInst_9_LFInst_3_n8 ,
         \Red_SubCellInst2_LFInst_9_LFInst_3_n7 ,
         \Red_SubCellInst2_LFInst_9_LFInst_3_n6 ,
         \Red_SubCellInst2_LFInst_10_LFInst_0_n14 ,
         \Red_SubCellInst2_LFInst_10_LFInst_0_n13 ,
         \Red_SubCellInst2_LFInst_10_LFInst_0_n12 ,
         \Red_SubCellInst2_LFInst_10_LFInst_0_n11 ,
         \Red_SubCellInst2_LFInst_10_LFInst_0_n10 ,
         \Red_SubCellInst2_LFInst_10_LFInst_0_n9 ,
         \Red_SubCellInst2_LFInst_10_LFInst_0_n8 ,
         \Red_SubCellInst2_LFInst_10_LFInst_1_n15 ,
         \Red_SubCellInst2_LFInst_10_LFInst_1_n14 ,
         \Red_SubCellInst2_LFInst_10_LFInst_1_n13 ,
         \Red_SubCellInst2_LFInst_10_LFInst_1_n12 ,
         \Red_SubCellInst2_LFInst_10_LFInst_1_n11 ,
         \Red_SubCellInst2_LFInst_10_LFInst_2_n19 ,
         \Red_SubCellInst2_LFInst_10_LFInst_2_n18 ,
         \Red_SubCellInst2_LFInst_10_LFInst_2_n17 ,
         \Red_SubCellInst2_LFInst_10_LFInst_2_n16 ,
         \Red_SubCellInst2_LFInst_10_LFInst_2_n15 ,
         \Red_SubCellInst2_LFInst_10_LFInst_2_n14 ,
         \Red_SubCellInst2_LFInst_10_LFInst_2_n13 ,
         \Red_SubCellInst2_LFInst_10_LFInst_3_n8 ,
         \Red_SubCellInst2_LFInst_10_LFInst_3_n7 ,
         \Red_SubCellInst2_LFInst_10_LFInst_3_n6 ,
         \Red_SubCellInst2_LFInst_11_LFInst_0_n14 ,
         \Red_SubCellInst2_LFInst_11_LFInst_0_n13 ,
         \Red_SubCellInst2_LFInst_11_LFInst_0_n12 ,
         \Red_SubCellInst2_LFInst_11_LFInst_0_n11 ,
         \Red_SubCellInst2_LFInst_11_LFInst_0_n10 ,
         \Red_SubCellInst2_LFInst_11_LFInst_0_n9 ,
         \Red_SubCellInst2_LFInst_11_LFInst_0_n8 ,
         \Red_SubCellInst2_LFInst_11_LFInst_1_n15 ,
         \Red_SubCellInst2_LFInst_11_LFInst_1_n14 ,
         \Red_SubCellInst2_LFInst_11_LFInst_1_n13 ,
         \Red_SubCellInst2_LFInst_11_LFInst_1_n12 ,
         \Red_SubCellInst2_LFInst_11_LFInst_1_n11 ,
         \Red_SubCellInst2_LFInst_11_LFInst_2_n19 ,
         \Red_SubCellInst2_LFInst_11_LFInst_2_n18 ,
         \Red_SubCellInst2_LFInst_11_LFInst_2_n17 ,
         \Red_SubCellInst2_LFInst_11_LFInst_2_n16 ,
         \Red_SubCellInst2_LFInst_11_LFInst_2_n15 ,
         \Red_SubCellInst2_LFInst_11_LFInst_2_n14 ,
         \Red_SubCellInst2_LFInst_11_LFInst_2_n13 ,
         \Red_SubCellInst2_LFInst_11_LFInst_3_n8 ,
         \Red_SubCellInst2_LFInst_11_LFInst_3_n7 ,
         \Red_SubCellInst2_LFInst_11_LFInst_3_n6 ,
         \Red_SubCellInst2_LFInst_12_LFInst_0_n14 ,
         \Red_SubCellInst2_LFInst_12_LFInst_0_n13 ,
         \Red_SubCellInst2_LFInst_12_LFInst_0_n12 ,
         \Red_SubCellInst2_LFInst_12_LFInst_0_n11 ,
         \Red_SubCellInst2_LFInst_12_LFInst_0_n10 ,
         \Red_SubCellInst2_LFInst_12_LFInst_0_n9 ,
         \Red_SubCellInst2_LFInst_12_LFInst_0_n8 ,
         \Red_SubCellInst2_LFInst_12_LFInst_1_n15 ,
         \Red_SubCellInst2_LFInst_12_LFInst_1_n14 ,
         \Red_SubCellInst2_LFInst_12_LFInst_1_n13 ,
         \Red_SubCellInst2_LFInst_12_LFInst_1_n12 ,
         \Red_SubCellInst2_LFInst_12_LFInst_1_n11 ,
         \Red_SubCellInst2_LFInst_12_LFInst_2_n19 ,
         \Red_SubCellInst2_LFInst_12_LFInst_2_n18 ,
         \Red_SubCellInst2_LFInst_12_LFInst_2_n17 ,
         \Red_SubCellInst2_LFInst_12_LFInst_2_n16 ,
         \Red_SubCellInst2_LFInst_12_LFInst_2_n15 ,
         \Red_SubCellInst2_LFInst_12_LFInst_2_n14 ,
         \Red_SubCellInst2_LFInst_12_LFInst_2_n13 ,
         \Red_SubCellInst2_LFInst_12_LFInst_3_n8 ,
         \Red_SubCellInst2_LFInst_12_LFInst_3_n7 ,
         \Red_SubCellInst2_LFInst_12_LFInst_3_n6 ,
         \Red_SubCellInst2_LFInst_13_LFInst_0_n14 ,
         \Red_SubCellInst2_LFInst_13_LFInst_0_n13 ,
         \Red_SubCellInst2_LFInst_13_LFInst_0_n12 ,
         \Red_SubCellInst2_LFInst_13_LFInst_0_n11 ,
         \Red_SubCellInst2_LFInst_13_LFInst_0_n10 ,
         \Red_SubCellInst2_LFInst_13_LFInst_0_n9 ,
         \Red_SubCellInst2_LFInst_13_LFInst_0_n8 ,
         \Red_SubCellInst2_LFInst_13_LFInst_1_n15 ,
         \Red_SubCellInst2_LFInst_13_LFInst_1_n14 ,
         \Red_SubCellInst2_LFInst_13_LFInst_1_n13 ,
         \Red_SubCellInst2_LFInst_13_LFInst_1_n12 ,
         \Red_SubCellInst2_LFInst_13_LFInst_1_n11 ,
         \Red_SubCellInst2_LFInst_13_LFInst_2_n19 ,
         \Red_SubCellInst2_LFInst_13_LFInst_2_n18 ,
         \Red_SubCellInst2_LFInst_13_LFInst_2_n17 ,
         \Red_SubCellInst2_LFInst_13_LFInst_2_n16 ,
         \Red_SubCellInst2_LFInst_13_LFInst_2_n15 ,
         \Red_SubCellInst2_LFInst_13_LFInst_2_n14 ,
         \Red_SubCellInst2_LFInst_13_LFInst_2_n13 ,
         \Red_SubCellInst2_LFInst_13_LFInst_3_n8 ,
         \Red_SubCellInst2_LFInst_13_LFInst_3_n7 ,
         \Red_SubCellInst2_LFInst_13_LFInst_3_n6 ,
         \Red_SubCellInst2_LFInst_14_LFInst_0_n14 ,
         \Red_SubCellInst2_LFInst_14_LFInst_0_n13 ,
         \Red_SubCellInst2_LFInst_14_LFInst_0_n12 ,
         \Red_SubCellInst2_LFInst_14_LFInst_0_n11 ,
         \Red_SubCellInst2_LFInst_14_LFInst_0_n10 ,
         \Red_SubCellInst2_LFInst_14_LFInst_0_n9 ,
         \Red_SubCellInst2_LFInst_14_LFInst_0_n8 ,
         \Red_SubCellInst2_LFInst_14_LFInst_1_n15 ,
         \Red_SubCellInst2_LFInst_14_LFInst_1_n14 ,
         \Red_SubCellInst2_LFInst_14_LFInst_1_n13 ,
         \Red_SubCellInst2_LFInst_14_LFInst_1_n12 ,
         \Red_SubCellInst2_LFInst_14_LFInst_1_n11 ,
         \Red_SubCellInst2_LFInst_14_LFInst_2_n19 ,
         \Red_SubCellInst2_LFInst_14_LFInst_2_n18 ,
         \Red_SubCellInst2_LFInst_14_LFInst_2_n17 ,
         \Red_SubCellInst2_LFInst_14_LFInst_2_n16 ,
         \Red_SubCellInst2_LFInst_14_LFInst_2_n15 ,
         \Red_SubCellInst2_LFInst_14_LFInst_2_n14 ,
         \Red_SubCellInst2_LFInst_14_LFInst_2_n13 ,
         \Red_SubCellInst2_LFInst_14_LFInst_3_n8 ,
         \Red_SubCellInst2_LFInst_14_LFInst_3_n7 ,
         \Red_SubCellInst2_LFInst_14_LFInst_3_n6 ,
         \Red_SubCellInst2_LFInst_15_LFInst_0_n14 ,
         \Red_SubCellInst2_LFInst_15_LFInst_0_n13 ,
         \Red_SubCellInst2_LFInst_15_LFInst_0_n12 ,
         \Red_SubCellInst2_LFInst_15_LFInst_0_n11 ,
         \Red_SubCellInst2_LFInst_15_LFInst_0_n10 ,
         \Red_SubCellInst2_LFInst_15_LFInst_0_n9 ,
         \Red_SubCellInst2_LFInst_15_LFInst_0_n8 ,
         \Red_SubCellInst2_LFInst_15_LFInst_1_n15 ,
         \Red_SubCellInst2_LFInst_15_LFInst_1_n14 ,
         \Red_SubCellInst2_LFInst_15_LFInst_1_n13 ,
         \Red_SubCellInst2_LFInst_15_LFInst_1_n12 ,
         \Red_SubCellInst2_LFInst_15_LFInst_1_n11 ,
         \Red_SubCellInst2_LFInst_15_LFInst_2_n19 ,
         \Red_SubCellInst2_LFInst_15_LFInst_2_n18 ,
         \Red_SubCellInst2_LFInst_15_LFInst_2_n17 ,
         \Red_SubCellInst2_LFInst_15_LFInst_2_n16 ,
         \Red_SubCellInst2_LFInst_15_LFInst_2_n15 ,
         \Red_SubCellInst2_LFInst_15_LFInst_2_n14 ,
         \Red_SubCellInst2_LFInst_15_LFInst_2_n13 ,
         \Red_SubCellInst2_LFInst_15_LFInst_3_n8 ,
         \Red_SubCellInst2_LFInst_15_LFInst_3_n7 ,
         \Red_SubCellInst2_LFInst_15_LFInst_3_n6 ,
         \Red_MCInst3_XOR_r0_Inst_0_n3 , \Red_MCInst3_XOR_r0_Inst_1_n3 ,
         \Red_MCInst3_XOR_r0_Inst_2_n3 , \Red_MCInst3_XOR_r0_Inst_3_n3 ,
         \Red_MCInst3_XOR_r0_Inst_4_n3 , \Red_MCInst3_XOR_r0_Inst_5_n3 ,
         \Red_MCInst3_XOR_r0_Inst_6_n3 , \Red_MCInst3_XOR_r0_Inst_7_n3 ,
         \Red_MCInst3_XOR_r0_Inst_8_n3 , \Red_MCInst3_XOR_r0_Inst_9_n3 ,
         \Red_MCInst3_XOR_r0_Inst_10_n3 , \Red_MCInst3_XOR_r0_Inst_11_n3 ,
         \Red_MCInst3_XOR_r0_Inst_12_n3 , \Red_MCInst3_XOR_r0_Inst_13_n3 ,
         \Red_MCInst3_XOR_r0_Inst_14_n3 , \Red_MCInst3_XOR_r0_Inst_15_n3 ,
         \Red_SubCellInst3_LFInst_0_LFInst_0_n14 ,
         \Red_SubCellInst3_LFInst_0_LFInst_0_n13 ,
         \Red_SubCellInst3_LFInst_0_LFInst_0_n12 ,
         \Red_SubCellInst3_LFInst_0_LFInst_0_n11 ,
         \Red_SubCellInst3_LFInst_0_LFInst_0_n10 ,
         \Red_SubCellInst3_LFInst_0_LFInst_0_n9 ,
         \Red_SubCellInst3_LFInst_0_LFInst_0_n8 ,
         \Red_SubCellInst3_LFInst_0_LFInst_1_n15 ,
         \Red_SubCellInst3_LFInst_0_LFInst_1_n14 ,
         \Red_SubCellInst3_LFInst_0_LFInst_1_n13 ,
         \Red_SubCellInst3_LFInst_0_LFInst_1_n12 ,
         \Red_SubCellInst3_LFInst_0_LFInst_1_n11 ,
         \Red_SubCellInst3_LFInst_0_LFInst_2_n19 ,
         \Red_SubCellInst3_LFInst_0_LFInst_2_n18 ,
         \Red_SubCellInst3_LFInst_0_LFInst_2_n17 ,
         \Red_SubCellInst3_LFInst_0_LFInst_2_n16 ,
         \Red_SubCellInst3_LFInst_0_LFInst_2_n15 ,
         \Red_SubCellInst3_LFInst_0_LFInst_2_n14 ,
         \Red_SubCellInst3_LFInst_0_LFInst_2_n13 ,
         \Red_SubCellInst3_LFInst_0_LFInst_3_n8 ,
         \Red_SubCellInst3_LFInst_0_LFInst_3_n7 ,
         \Red_SubCellInst3_LFInst_0_LFInst_3_n6 ,
         \Red_SubCellInst3_LFInst_1_LFInst_0_n14 ,
         \Red_SubCellInst3_LFInst_1_LFInst_0_n13 ,
         \Red_SubCellInst3_LFInst_1_LFInst_0_n12 ,
         \Red_SubCellInst3_LFInst_1_LFInst_0_n11 ,
         \Red_SubCellInst3_LFInst_1_LFInst_0_n10 ,
         \Red_SubCellInst3_LFInst_1_LFInst_0_n9 ,
         \Red_SubCellInst3_LFInst_1_LFInst_0_n8 ,
         \Red_SubCellInst3_LFInst_1_LFInst_1_n15 ,
         \Red_SubCellInst3_LFInst_1_LFInst_1_n14 ,
         \Red_SubCellInst3_LFInst_1_LFInst_1_n13 ,
         \Red_SubCellInst3_LFInst_1_LFInst_1_n12 ,
         \Red_SubCellInst3_LFInst_1_LFInst_1_n11 ,
         \Red_SubCellInst3_LFInst_1_LFInst_2_n19 ,
         \Red_SubCellInst3_LFInst_1_LFInst_2_n18 ,
         \Red_SubCellInst3_LFInst_1_LFInst_2_n17 ,
         \Red_SubCellInst3_LFInst_1_LFInst_2_n16 ,
         \Red_SubCellInst3_LFInst_1_LFInst_2_n15 ,
         \Red_SubCellInst3_LFInst_1_LFInst_2_n14 ,
         \Red_SubCellInst3_LFInst_1_LFInst_2_n13 ,
         \Red_SubCellInst3_LFInst_1_LFInst_3_n8 ,
         \Red_SubCellInst3_LFInst_1_LFInst_3_n7 ,
         \Red_SubCellInst3_LFInst_1_LFInst_3_n6 ,
         \Red_SubCellInst3_LFInst_2_LFInst_0_n14 ,
         \Red_SubCellInst3_LFInst_2_LFInst_0_n13 ,
         \Red_SubCellInst3_LFInst_2_LFInst_0_n12 ,
         \Red_SubCellInst3_LFInst_2_LFInst_0_n11 ,
         \Red_SubCellInst3_LFInst_2_LFInst_0_n10 ,
         \Red_SubCellInst3_LFInst_2_LFInst_0_n9 ,
         \Red_SubCellInst3_LFInst_2_LFInst_0_n8 ,
         \Red_SubCellInst3_LFInst_2_LFInst_1_n15 ,
         \Red_SubCellInst3_LFInst_2_LFInst_1_n14 ,
         \Red_SubCellInst3_LFInst_2_LFInst_1_n13 ,
         \Red_SubCellInst3_LFInst_2_LFInst_1_n12 ,
         \Red_SubCellInst3_LFInst_2_LFInst_1_n11 ,
         \Red_SubCellInst3_LFInst_2_LFInst_2_n19 ,
         \Red_SubCellInst3_LFInst_2_LFInst_2_n18 ,
         \Red_SubCellInst3_LFInst_2_LFInst_2_n17 ,
         \Red_SubCellInst3_LFInst_2_LFInst_2_n16 ,
         \Red_SubCellInst3_LFInst_2_LFInst_2_n15 ,
         \Red_SubCellInst3_LFInst_2_LFInst_2_n14 ,
         \Red_SubCellInst3_LFInst_2_LFInst_2_n13 ,
         \Red_SubCellInst3_LFInst_2_LFInst_3_n8 ,
         \Red_SubCellInst3_LFInst_2_LFInst_3_n7 ,
         \Red_SubCellInst3_LFInst_2_LFInst_3_n6 ,
         \Red_SubCellInst3_LFInst_3_LFInst_0_n14 ,
         \Red_SubCellInst3_LFInst_3_LFInst_0_n13 ,
         \Red_SubCellInst3_LFInst_3_LFInst_0_n12 ,
         \Red_SubCellInst3_LFInst_3_LFInst_0_n11 ,
         \Red_SubCellInst3_LFInst_3_LFInst_0_n10 ,
         \Red_SubCellInst3_LFInst_3_LFInst_0_n9 ,
         \Red_SubCellInst3_LFInst_3_LFInst_0_n8 ,
         \Red_SubCellInst3_LFInst_3_LFInst_1_n15 ,
         \Red_SubCellInst3_LFInst_3_LFInst_1_n14 ,
         \Red_SubCellInst3_LFInst_3_LFInst_1_n13 ,
         \Red_SubCellInst3_LFInst_3_LFInst_1_n12 ,
         \Red_SubCellInst3_LFInst_3_LFInst_1_n11 ,
         \Red_SubCellInst3_LFInst_3_LFInst_2_n19 ,
         \Red_SubCellInst3_LFInst_3_LFInst_2_n18 ,
         \Red_SubCellInst3_LFInst_3_LFInst_2_n17 ,
         \Red_SubCellInst3_LFInst_3_LFInst_2_n16 ,
         \Red_SubCellInst3_LFInst_3_LFInst_2_n15 ,
         \Red_SubCellInst3_LFInst_3_LFInst_2_n14 ,
         \Red_SubCellInst3_LFInst_3_LFInst_2_n13 ,
         \Red_SubCellInst3_LFInst_3_LFInst_3_n8 ,
         \Red_SubCellInst3_LFInst_3_LFInst_3_n7 ,
         \Red_SubCellInst3_LFInst_3_LFInst_3_n6 ,
         \Red_SubCellInst3_LFInst_4_LFInst_0_n14 ,
         \Red_SubCellInst3_LFInst_4_LFInst_0_n13 ,
         \Red_SubCellInst3_LFInst_4_LFInst_0_n12 ,
         \Red_SubCellInst3_LFInst_4_LFInst_0_n11 ,
         \Red_SubCellInst3_LFInst_4_LFInst_0_n10 ,
         \Red_SubCellInst3_LFInst_4_LFInst_0_n9 ,
         \Red_SubCellInst3_LFInst_4_LFInst_0_n8 ,
         \Red_SubCellInst3_LFInst_4_LFInst_1_n15 ,
         \Red_SubCellInst3_LFInst_4_LFInst_1_n14 ,
         \Red_SubCellInst3_LFInst_4_LFInst_1_n13 ,
         \Red_SubCellInst3_LFInst_4_LFInst_1_n12 ,
         \Red_SubCellInst3_LFInst_4_LFInst_1_n11 ,
         \Red_SubCellInst3_LFInst_4_LFInst_2_n19 ,
         \Red_SubCellInst3_LFInst_4_LFInst_2_n18 ,
         \Red_SubCellInst3_LFInst_4_LFInst_2_n17 ,
         \Red_SubCellInst3_LFInst_4_LFInst_2_n16 ,
         \Red_SubCellInst3_LFInst_4_LFInst_2_n15 ,
         \Red_SubCellInst3_LFInst_4_LFInst_2_n14 ,
         \Red_SubCellInst3_LFInst_4_LFInst_2_n13 ,
         \Red_SubCellInst3_LFInst_4_LFInst_3_n8 ,
         \Red_SubCellInst3_LFInst_4_LFInst_3_n7 ,
         \Red_SubCellInst3_LFInst_4_LFInst_3_n6 ,
         \Red_SubCellInst3_LFInst_5_LFInst_0_n14 ,
         \Red_SubCellInst3_LFInst_5_LFInst_0_n13 ,
         \Red_SubCellInst3_LFInst_5_LFInst_0_n12 ,
         \Red_SubCellInst3_LFInst_5_LFInst_0_n11 ,
         \Red_SubCellInst3_LFInst_5_LFInst_0_n10 ,
         \Red_SubCellInst3_LFInst_5_LFInst_0_n9 ,
         \Red_SubCellInst3_LFInst_5_LFInst_0_n8 ,
         \Red_SubCellInst3_LFInst_5_LFInst_1_n15 ,
         \Red_SubCellInst3_LFInst_5_LFInst_1_n14 ,
         \Red_SubCellInst3_LFInst_5_LFInst_1_n13 ,
         \Red_SubCellInst3_LFInst_5_LFInst_1_n12 ,
         \Red_SubCellInst3_LFInst_5_LFInst_1_n11 ,
         \Red_SubCellInst3_LFInst_5_LFInst_2_n19 ,
         \Red_SubCellInst3_LFInst_5_LFInst_2_n18 ,
         \Red_SubCellInst3_LFInst_5_LFInst_2_n17 ,
         \Red_SubCellInst3_LFInst_5_LFInst_2_n16 ,
         \Red_SubCellInst3_LFInst_5_LFInst_2_n15 ,
         \Red_SubCellInst3_LFInst_5_LFInst_2_n14 ,
         \Red_SubCellInst3_LFInst_5_LFInst_2_n13 ,
         \Red_SubCellInst3_LFInst_5_LFInst_3_n8 ,
         \Red_SubCellInst3_LFInst_5_LFInst_3_n7 ,
         \Red_SubCellInst3_LFInst_5_LFInst_3_n6 ,
         \Red_SubCellInst3_LFInst_6_LFInst_0_n14 ,
         \Red_SubCellInst3_LFInst_6_LFInst_0_n13 ,
         \Red_SubCellInst3_LFInst_6_LFInst_0_n12 ,
         \Red_SubCellInst3_LFInst_6_LFInst_0_n11 ,
         \Red_SubCellInst3_LFInst_6_LFInst_0_n10 ,
         \Red_SubCellInst3_LFInst_6_LFInst_0_n9 ,
         \Red_SubCellInst3_LFInst_6_LFInst_0_n8 ,
         \Red_SubCellInst3_LFInst_6_LFInst_1_n15 ,
         \Red_SubCellInst3_LFInst_6_LFInst_1_n14 ,
         \Red_SubCellInst3_LFInst_6_LFInst_1_n13 ,
         \Red_SubCellInst3_LFInst_6_LFInst_1_n12 ,
         \Red_SubCellInst3_LFInst_6_LFInst_1_n11 ,
         \Red_SubCellInst3_LFInst_6_LFInst_2_n19 ,
         \Red_SubCellInst3_LFInst_6_LFInst_2_n18 ,
         \Red_SubCellInst3_LFInst_6_LFInst_2_n17 ,
         \Red_SubCellInst3_LFInst_6_LFInst_2_n16 ,
         \Red_SubCellInst3_LFInst_6_LFInst_2_n15 ,
         \Red_SubCellInst3_LFInst_6_LFInst_2_n14 ,
         \Red_SubCellInst3_LFInst_6_LFInst_2_n13 ,
         \Red_SubCellInst3_LFInst_6_LFInst_3_n8 ,
         \Red_SubCellInst3_LFInst_6_LFInst_3_n7 ,
         \Red_SubCellInst3_LFInst_6_LFInst_3_n6 ,
         \Red_SubCellInst3_LFInst_7_LFInst_0_n14 ,
         \Red_SubCellInst3_LFInst_7_LFInst_0_n13 ,
         \Red_SubCellInst3_LFInst_7_LFInst_0_n12 ,
         \Red_SubCellInst3_LFInst_7_LFInst_0_n11 ,
         \Red_SubCellInst3_LFInst_7_LFInst_0_n10 ,
         \Red_SubCellInst3_LFInst_7_LFInst_0_n9 ,
         \Red_SubCellInst3_LFInst_7_LFInst_0_n8 ,
         \Red_SubCellInst3_LFInst_7_LFInst_1_n15 ,
         \Red_SubCellInst3_LFInst_7_LFInst_1_n14 ,
         \Red_SubCellInst3_LFInst_7_LFInst_1_n13 ,
         \Red_SubCellInst3_LFInst_7_LFInst_1_n12 ,
         \Red_SubCellInst3_LFInst_7_LFInst_1_n11 ,
         \Red_SubCellInst3_LFInst_7_LFInst_2_n19 ,
         \Red_SubCellInst3_LFInst_7_LFInst_2_n18 ,
         \Red_SubCellInst3_LFInst_7_LFInst_2_n17 ,
         \Red_SubCellInst3_LFInst_7_LFInst_2_n16 ,
         \Red_SubCellInst3_LFInst_7_LFInst_2_n15 ,
         \Red_SubCellInst3_LFInst_7_LFInst_2_n14 ,
         \Red_SubCellInst3_LFInst_7_LFInst_2_n13 ,
         \Red_SubCellInst3_LFInst_7_LFInst_3_n8 ,
         \Red_SubCellInst3_LFInst_7_LFInst_3_n7 ,
         \Red_SubCellInst3_LFInst_7_LFInst_3_n6 ,
         \Red_SubCellInst3_LFInst_8_LFInst_0_n14 ,
         \Red_SubCellInst3_LFInst_8_LFInst_0_n13 ,
         \Red_SubCellInst3_LFInst_8_LFInst_0_n12 ,
         \Red_SubCellInst3_LFInst_8_LFInst_0_n11 ,
         \Red_SubCellInst3_LFInst_8_LFInst_0_n10 ,
         \Red_SubCellInst3_LFInst_8_LFInst_0_n9 ,
         \Red_SubCellInst3_LFInst_8_LFInst_0_n8 ,
         \Red_SubCellInst3_LFInst_8_LFInst_1_n15 ,
         \Red_SubCellInst3_LFInst_8_LFInst_1_n14 ,
         \Red_SubCellInst3_LFInst_8_LFInst_1_n13 ,
         \Red_SubCellInst3_LFInst_8_LFInst_1_n12 ,
         \Red_SubCellInst3_LFInst_8_LFInst_1_n11 ,
         \Red_SubCellInst3_LFInst_8_LFInst_2_n19 ,
         \Red_SubCellInst3_LFInst_8_LFInst_2_n18 ,
         \Red_SubCellInst3_LFInst_8_LFInst_2_n17 ,
         \Red_SubCellInst3_LFInst_8_LFInst_2_n16 ,
         \Red_SubCellInst3_LFInst_8_LFInst_2_n15 ,
         \Red_SubCellInst3_LFInst_8_LFInst_2_n14 ,
         \Red_SubCellInst3_LFInst_8_LFInst_2_n13 ,
         \Red_SubCellInst3_LFInst_8_LFInst_3_n8 ,
         \Red_SubCellInst3_LFInst_8_LFInst_3_n7 ,
         \Red_SubCellInst3_LFInst_8_LFInst_3_n6 ,
         \Red_SubCellInst3_LFInst_9_LFInst_0_n14 ,
         \Red_SubCellInst3_LFInst_9_LFInst_0_n13 ,
         \Red_SubCellInst3_LFInst_9_LFInst_0_n12 ,
         \Red_SubCellInst3_LFInst_9_LFInst_0_n11 ,
         \Red_SubCellInst3_LFInst_9_LFInst_0_n10 ,
         \Red_SubCellInst3_LFInst_9_LFInst_0_n9 ,
         \Red_SubCellInst3_LFInst_9_LFInst_0_n8 ,
         \Red_SubCellInst3_LFInst_9_LFInst_1_n15 ,
         \Red_SubCellInst3_LFInst_9_LFInst_1_n14 ,
         \Red_SubCellInst3_LFInst_9_LFInst_1_n13 ,
         \Red_SubCellInst3_LFInst_9_LFInst_1_n12 ,
         \Red_SubCellInst3_LFInst_9_LFInst_1_n11 ,
         \Red_SubCellInst3_LFInst_9_LFInst_2_n19 ,
         \Red_SubCellInst3_LFInst_9_LFInst_2_n18 ,
         \Red_SubCellInst3_LFInst_9_LFInst_2_n17 ,
         \Red_SubCellInst3_LFInst_9_LFInst_2_n16 ,
         \Red_SubCellInst3_LFInst_9_LFInst_2_n15 ,
         \Red_SubCellInst3_LFInst_9_LFInst_2_n14 ,
         \Red_SubCellInst3_LFInst_9_LFInst_2_n13 ,
         \Red_SubCellInst3_LFInst_9_LFInst_3_n8 ,
         \Red_SubCellInst3_LFInst_9_LFInst_3_n7 ,
         \Red_SubCellInst3_LFInst_9_LFInst_3_n6 ,
         \Red_SubCellInst3_LFInst_10_LFInst_0_n14 ,
         \Red_SubCellInst3_LFInst_10_LFInst_0_n13 ,
         \Red_SubCellInst3_LFInst_10_LFInst_0_n12 ,
         \Red_SubCellInst3_LFInst_10_LFInst_0_n11 ,
         \Red_SubCellInst3_LFInst_10_LFInst_0_n10 ,
         \Red_SubCellInst3_LFInst_10_LFInst_0_n9 ,
         \Red_SubCellInst3_LFInst_10_LFInst_0_n8 ,
         \Red_SubCellInst3_LFInst_10_LFInst_1_n15 ,
         \Red_SubCellInst3_LFInst_10_LFInst_1_n14 ,
         \Red_SubCellInst3_LFInst_10_LFInst_1_n13 ,
         \Red_SubCellInst3_LFInst_10_LFInst_1_n12 ,
         \Red_SubCellInst3_LFInst_10_LFInst_1_n11 ,
         \Red_SubCellInst3_LFInst_10_LFInst_2_n19 ,
         \Red_SubCellInst3_LFInst_10_LFInst_2_n18 ,
         \Red_SubCellInst3_LFInst_10_LFInst_2_n17 ,
         \Red_SubCellInst3_LFInst_10_LFInst_2_n16 ,
         \Red_SubCellInst3_LFInst_10_LFInst_2_n15 ,
         \Red_SubCellInst3_LFInst_10_LFInst_2_n14 ,
         \Red_SubCellInst3_LFInst_10_LFInst_2_n13 ,
         \Red_SubCellInst3_LFInst_10_LFInst_3_n8 ,
         \Red_SubCellInst3_LFInst_10_LFInst_3_n7 ,
         \Red_SubCellInst3_LFInst_10_LFInst_3_n6 ,
         \Red_SubCellInst3_LFInst_11_LFInst_0_n14 ,
         \Red_SubCellInst3_LFInst_11_LFInst_0_n13 ,
         \Red_SubCellInst3_LFInst_11_LFInst_0_n12 ,
         \Red_SubCellInst3_LFInst_11_LFInst_0_n11 ,
         \Red_SubCellInst3_LFInst_11_LFInst_0_n10 ,
         \Red_SubCellInst3_LFInst_11_LFInst_0_n9 ,
         \Red_SubCellInst3_LFInst_11_LFInst_0_n8 ,
         \Red_SubCellInst3_LFInst_11_LFInst_1_n15 ,
         \Red_SubCellInst3_LFInst_11_LFInst_1_n14 ,
         \Red_SubCellInst3_LFInst_11_LFInst_1_n13 ,
         \Red_SubCellInst3_LFInst_11_LFInst_1_n12 ,
         \Red_SubCellInst3_LFInst_11_LFInst_1_n11 ,
         \Red_SubCellInst3_LFInst_11_LFInst_2_n19 ,
         \Red_SubCellInst3_LFInst_11_LFInst_2_n18 ,
         \Red_SubCellInst3_LFInst_11_LFInst_2_n17 ,
         \Red_SubCellInst3_LFInst_11_LFInst_2_n16 ,
         \Red_SubCellInst3_LFInst_11_LFInst_2_n15 ,
         \Red_SubCellInst3_LFInst_11_LFInst_2_n14 ,
         \Red_SubCellInst3_LFInst_11_LFInst_2_n13 ,
         \Red_SubCellInst3_LFInst_11_LFInst_3_n8 ,
         \Red_SubCellInst3_LFInst_11_LFInst_3_n7 ,
         \Red_SubCellInst3_LFInst_11_LFInst_3_n6 ,
         \Red_SubCellInst3_LFInst_12_LFInst_0_n14 ,
         \Red_SubCellInst3_LFInst_12_LFInst_0_n13 ,
         \Red_SubCellInst3_LFInst_12_LFInst_0_n12 ,
         \Red_SubCellInst3_LFInst_12_LFInst_0_n11 ,
         \Red_SubCellInst3_LFInst_12_LFInst_0_n10 ,
         \Red_SubCellInst3_LFInst_12_LFInst_0_n9 ,
         \Red_SubCellInst3_LFInst_12_LFInst_0_n8 ,
         \Red_SubCellInst3_LFInst_12_LFInst_1_n15 ,
         \Red_SubCellInst3_LFInst_12_LFInst_1_n14 ,
         \Red_SubCellInst3_LFInst_12_LFInst_1_n13 ,
         \Red_SubCellInst3_LFInst_12_LFInst_1_n12 ,
         \Red_SubCellInst3_LFInst_12_LFInst_1_n11 ,
         \Red_SubCellInst3_LFInst_12_LFInst_2_n19 ,
         \Red_SubCellInst3_LFInst_12_LFInst_2_n18 ,
         \Red_SubCellInst3_LFInst_12_LFInst_2_n17 ,
         \Red_SubCellInst3_LFInst_12_LFInst_2_n16 ,
         \Red_SubCellInst3_LFInst_12_LFInst_2_n15 ,
         \Red_SubCellInst3_LFInst_12_LFInst_2_n14 ,
         \Red_SubCellInst3_LFInst_12_LFInst_2_n13 ,
         \Red_SubCellInst3_LFInst_12_LFInst_3_n8 ,
         \Red_SubCellInst3_LFInst_12_LFInst_3_n7 ,
         \Red_SubCellInst3_LFInst_12_LFInst_3_n6 ,
         \Red_SubCellInst3_LFInst_13_LFInst_0_n14 ,
         \Red_SubCellInst3_LFInst_13_LFInst_0_n13 ,
         \Red_SubCellInst3_LFInst_13_LFInst_0_n12 ,
         \Red_SubCellInst3_LFInst_13_LFInst_0_n11 ,
         \Red_SubCellInst3_LFInst_13_LFInst_0_n10 ,
         \Red_SubCellInst3_LFInst_13_LFInst_0_n9 ,
         \Red_SubCellInst3_LFInst_13_LFInst_0_n8 ,
         \Red_SubCellInst3_LFInst_13_LFInst_1_n15 ,
         \Red_SubCellInst3_LFInst_13_LFInst_1_n14 ,
         \Red_SubCellInst3_LFInst_13_LFInst_1_n13 ,
         \Red_SubCellInst3_LFInst_13_LFInst_1_n12 ,
         \Red_SubCellInst3_LFInst_13_LFInst_1_n11 ,
         \Red_SubCellInst3_LFInst_13_LFInst_2_n19 ,
         \Red_SubCellInst3_LFInst_13_LFInst_2_n18 ,
         \Red_SubCellInst3_LFInst_13_LFInst_2_n17 ,
         \Red_SubCellInst3_LFInst_13_LFInst_2_n16 ,
         \Red_SubCellInst3_LFInst_13_LFInst_2_n15 ,
         \Red_SubCellInst3_LFInst_13_LFInst_2_n14 ,
         \Red_SubCellInst3_LFInst_13_LFInst_2_n13 ,
         \Red_SubCellInst3_LFInst_13_LFInst_3_n8 ,
         \Red_SubCellInst3_LFInst_13_LFInst_3_n7 ,
         \Red_SubCellInst3_LFInst_13_LFInst_3_n6 ,
         \Red_SubCellInst3_LFInst_14_LFInst_0_n14 ,
         \Red_SubCellInst3_LFInst_14_LFInst_0_n13 ,
         \Red_SubCellInst3_LFInst_14_LFInst_0_n12 ,
         \Red_SubCellInst3_LFInst_14_LFInst_0_n11 ,
         \Red_SubCellInst3_LFInst_14_LFInst_0_n10 ,
         \Red_SubCellInst3_LFInst_14_LFInst_0_n9 ,
         \Red_SubCellInst3_LFInst_14_LFInst_0_n8 ,
         \Red_SubCellInst3_LFInst_14_LFInst_1_n15 ,
         \Red_SubCellInst3_LFInst_14_LFInst_1_n14 ,
         \Red_SubCellInst3_LFInst_14_LFInst_1_n13 ,
         \Red_SubCellInst3_LFInst_14_LFInst_1_n12 ,
         \Red_SubCellInst3_LFInst_14_LFInst_1_n11 ,
         \Red_SubCellInst3_LFInst_14_LFInst_2_n19 ,
         \Red_SubCellInst3_LFInst_14_LFInst_2_n18 ,
         \Red_SubCellInst3_LFInst_14_LFInst_2_n17 ,
         \Red_SubCellInst3_LFInst_14_LFInst_2_n16 ,
         \Red_SubCellInst3_LFInst_14_LFInst_2_n15 ,
         \Red_SubCellInst3_LFInst_14_LFInst_2_n14 ,
         \Red_SubCellInst3_LFInst_14_LFInst_2_n13 ,
         \Red_SubCellInst3_LFInst_14_LFInst_3_n8 ,
         \Red_SubCellInst3_LFInst_14_LFInst_3_n7 ,
         \Red_SubCellInst3_LFInst_14_LFInst_3_n6 ,
         \Red_SubCellInst3_LFInst_15_LFInst_0_n14 ,
         \Red_SubCellInst3_LFInst_15_LFInst_0_n13 ,
         \Red_SubCellInst3_LFInst_15_LFInst_0_n12 ,
         \Red_SubCellInst3_LFInst_15_LFInst_0_n11 ,
         \Red_SubCellInst3_LFInst_15_LFInst_0_n10 ,
         \Red_SubCellInst3_LFInst_15_LFInst_0_n9 ,
         \Red_SubCellInst3_LFInst_15_LFInst_0_n8 ,
         \Red_SubCellInst3_LFInst_15_LFInst_1_n15 ,
         \Red_SubCellInst3_LFInst_15_LFInst_1_n14 ,
         \Red_SubCellInst3_LFInst_15_LFInst_1_n13 ,
         \Red_SubCellInst3_LFInst_15_LFInst_1_n12 ,
         \Red_SubCellInst3_LFInst_15_LFInst_1_n11 ,
         \Red_SubCellInst3_LFInst_15_LFInst_2_n19 ,
         \Red_SubCellInst3_LFInst_15_LFInst_2_n18 ,
         \Red_SubCellInst3_LFInst_15_LFInst_2_n17 ,
         \Red_SubCellInst3_LFInst_15_LFInst_2_n16 ,
         \Red_SubCellInst3_LFInst_15_LFInst_2_n15 ,
         \Red_SubCellInst3_LFInst_15_LFInst_2_n14 ,
         \Red_SubCellInst3_LFInst_15_LFInst_2_n13 ,
         \Red_SubCellInst3_LFInst_15_LFInst_3_n8 ,
         \Red_SubCellInst3_LFInst_15_LFInst_3_n7 ,
         \Red_SubCellInst3_LFInst_15_LFInst_3_n6 ,
         \Red_K0Inst_LFInst_0_LFInst_0_n2 , \Red_K0Inst_LFInst_0_LFInst_1_n2 ,
         \Red_K0Inst_LFInst_0_LFInst_2_n2 , \Red_K0Inst_LFInst_0_LFInst_3_n2 ,
         \Red_K0Inst_LFInst_1_LFInst_0_n2 , \Red_K0Inst_LFInst_1_LFInst_1_n2 ,
         \Red_K0Inst_LFInst_1_LFInst_2_n2 , \Red_K0Inst_LFInst_1_LFInst_3_n2 ,
         \Red_K0Inst_LFInst_2_LFInst_0_n2 , \Red_K0Inst_LFInst_2_LFInst_1_n2 ,
         \Red_K0Inst_LFInst_2_LFInst_2_n2 , \Red_K0Inst_LFInst_2_LFInst_3_n2 ,
         \Red_K0Inst_LFInst_3_LFInst_0_n2 , \Red_K0Inst_LFInst_3_LFInst_1_n2 ,
         \Red_K0Inst_LFInst_3_LFInst_2_n2 , \Red_K0Inst_LFInst_3_LFInst_3_n2 ,
         \Red_K0Inst_LFInst_4_LFInst_0_n2 , \Red_K0Inst_LFInst_4_LFInst_1_n2 ,
         \Red_K0Inst_LFInst_4_LFInst_2_n2 , \Red_K0Inst_LFInst_4_LFInst_3_n2 ,
         \Red_K0Inst_LFInst_5_LFInst_0_n2 , \Red_K0Inst_LFInst_5_LFInst_1_n2 ,
         \Red_K0Inst_LFInst_5_LFInst_2_n2 , \Red_K0Inst_LFInst_5_LFInst_3_n2 ,
         \Red_K0Inst_LFInst_6_LFInst_0_n2 , \Red_K0Inst_LFInst_6_LFInst_1_n2 ,
         \Red_K0Inst_LFInst_6_LFInst_2_n2 , \Red_K0Inst_LFInst_6_LFInst_3_n2 ,
         \Red_K0Inst_LFInst_7_LFInst_0_n2 , \Red_K0Inst_LFInst_7_LFInst_1_n2 ,
         \Red_K0Inst_LFInst_7_LFInst_2_n2 , \Red_K0Inst_LFInst_7_LFInst_3_n2 ,
         \Red_K0Inst_LFInst_8_LFInst_0_n2 , \Red_K0Inst_LFInst_8_LFInst_1_n2 ,
         \Red_K0Inst_LFInst_8_LFInst_2_n2 , \Red_K0Inst_LFInst_8_LFInst_3_n2 ,
         \Red_K0Inst_LFInst_9_LFInst_0_n2 , \Red_K0Inst_LFInst_9_LFInst_1_n2 ,
         \Red_K0Inst_LFInst_9_LFInst_2_n2 , \Red_K0Inst_LFInst_9_LFInst_3_n2 ,
         \Red_K0Inst_LFInst_10_LFInst_0_n2 ,
         \Red_K0Inst_LFInst_10_LFInst_1_n2 ,
         \Red_K0Inst_LFInst_10_LFInst_2_n2 ,
         \Red_K0Inst_LFInst_10_LFInst_3_n2 ,
         \Red_K0Inst_LFInst_11_LFInst_0_n2 ,
         \Red_K0Inst_LFInst_11_LFInst_1_n2 ,
         \Red_K0Inst_LFInst_11_LFInst_2_n2 ,
         \Red_K0Inst_LFInst_11_LFInst_3_n2 ,
         \Red_K0Inst_LFInst_12_LFInst_0_n2 ,
         \Red_K0Inst_LFInst_12_LFInst_1_n2 ,
         \Red_K0Inst_LFInst_12_LFInst_2_n2 ,
         \Red_K0Inst_LFInst_12_LFInst_3_n2 ,
         \Red_K0Inst_LFInst_13_LFInst_0_n2 ,
         \Red_K0Inst_LFInst_13_LFInst_1_n2 ,
         \Red_K0Inst_LFInst_13_LFInst_2_n2 ,
         \Red_K0Inst_LFInst_13_LFInst_3_n2 ,
         \Red_K0Inst_LFInst_14_LFInst_0_n2 ,
         \Red_K0Inst_LFInst_14_LFInst_1_n2 ,
         \Red_K0Inst_LFInst_14_LFInst_2_n2 ,
         \Red_K0Inst_LFInst_14_LFInst_3_n2 ,
         \Red_K0Inst_LFInst_15_LFInst_0_n2 ,
         \Red_K0Inst_LFInst_15_LFInst_1_n2 ,
         \Red_K0Inst_LFInst_15_LFInst_2_n2 ,
         \Red_K0Inst_LFInst_15_LFInst_3_n2 , \Red_K1Inst_LFInst_0_LFInst_0_n2 ,
         \Red_K1Inst_LFInst_0_LFInst_1_n2 , \Red_K1Inst_LFInst_0_LFInst_2_n2 ,
         \Red_K1Inst_LFInst_0_LFInst_3_n2 , \Red_K1Inst_LFInst_1_LFInst_0_n2 ,
         \Red_K1Inst_LFInst_1_LFInst_1_n2 , \Red_K1Inst_LFInst_1_LFInst_2_n2 ,
         \Red_K1Inst_LFInst_1_LFInst_3_n2 , \Red_K1Inst_LFInst_2_LFInst_0_n2 ,
         \Red_K1Inst_LFInst_2_LFInst_1_n2 , \Red_K1Inst_LFInst_2_LFInst_2_n2 ,
         \Red_K1Inst_LFInst_2_LFInst_3_n2 , \Red_K1Inst_LFInst_3_LFInst_0_n2 ,
         \Red_K1Inst_LFInst_3_LFInst_1_n2 , \Red_K1Inst_LFInst_3_LFInst_2_n2 ,
         \Red_K1Inst_LFInst_3_LFInst_3_n2 , \Red_K1Inst_LFInst_4_LFInst_0_n2 ,
         \Red_K1Inst_LFInst_4_LFInst_1_n2 , \Red_K1Inst_LFInst_4_LFInst_2_n2 ,
         \Red_K1Inst_LFInst_4_LFInst_3_n2 , \Red_K1Inst_LFInst_5_LFInst_0_n2 ,
         \Red_K1Inst_LFInst_5_LFInst_1_n2 , \Red_K1Inst_LFInst_5_LFInst_2_n2 ,
         \Red_K1Inst_LFInst_5_LFInst_3_n2 , \Red_K1Inst_LFInst_6_LFInst_0_n2 ,
         \Red_K1Inst_LFInst_6_LFInst_1_n2 , \Red_K1Inst_LFInst_6_LFInst_2_n2 ,
         \Red_K1Inst_LFInst_6_LFInst_3_n2 , \Red_K1Inst_LFInst_7_LFInst_0_n2 ,
         \Red_K1Inst_LFInst_7_LFInst_1_n2 , \Red_K1Inst_LFInst_7_LFInst_2_n2 ,
         \Red_K1Inst_LFInst_7_LFInst_3_n2 , \Red_K1Inst_LFInst_8_LFInst_0_n2 ,
         \Red_K1Inst_LFInst_8_LFInst_1_n2 , \Red_K1Inst_LFInst_8_LFInst_2_n2 ,
         \Red_K1Inst_LFInst_8_LFInst_3_n2 , \Red_K1Inst_LFInst_9_LFInst_0_n2 ,
         \Red_K1Inst_LFInst_9_LFInst_1_n2 , \Red_K1Inst_LFInst_9_LFInst_2_n2 ,
         \Red_K1Inst_LFInst_9_LFInst_3_n2 , \Red_K1Inst_LFInst_10_LFInst_0_n2 ,
         \Red_K1Inst_LFInst_10_LFInst_1_n2 ,
         \Red_K1Inst_LFInst_10_LFInst_2_n2 ,
         \Red_K1Inst_LFInst_10_LFInst_3_n2 ,
         \Red_K1Inst_LFInst_11_LFInst_0_n2 ,
         \Red_K1Inst_LFInst_11_LFInst_1_n2 ,
         \Red_K1Inst_LFInst_11_LFInst_2_n2 ,
         \Red_K1Inst_LFInst_11_LFInst_3_n2 ,
         \Red_K1Inst_LFInst_12_LFInst_0_n2 ,
         \Red_K1Inst_LFInst_12_LFInst_1_n2 ,
         \Red_K1Inst_LFInst_12_LFInst_2_n2 ,
         \Red_K1Inst_LFInst_12_LFInst_3_n2 ,
         \Red_K1Inst_LFInst_13_LFInst_0_n2 ,
         \Red_K1Inst_LFInst_13_LFInst_1_n2 ,
         \Red_K1Inst_LFInst_13_LFInst_2_n2 ,
         \Red_K1Inst_LFInst_13_LFInst_3_n2 ,
         \Red_K1Inst_LFInst_14_LFInst_0_n2 ,
         \Red_K1Inst_LFInst_14_LFInst_1_n2 ,
         \Red_K1Inst_LFInst_14_LFInst_2_n2 ,
         \Red_K1Inst_LFInst_14_LFInst_3_n2 ,
         \Red_K1Inst_LFInst_15_LFInst_0_n2 ,
         \Red_K1Inst_LFInst_15_LFInst_1_n2 ,
         \Red_K1Inst_LFInst_15_LFInst_2_n2 ,
         \Red_K1Inst_LFInst_15_LFInst_3_n2 , \Red_K2Inst_LFInst_0_LFInst_0_n2 ,
         \Red_K2Inst_LFInst_0_LFInst_1_n2 , \Red_K2Inst_LFInst_0_LFInst_2_n2 ,
         \Red_K2Inst_LFInst_0_LFInst_3_n2 , \Red_K2Inst_LFInst_1_LFInst_0_n2 ,
         \Red_K2Inst_LFInst_1_LFInst_1_n2 , \Red_K2Inst_LFInst_1_LFInst_2_n2 ,
         \Red_K2Inst_LFInst_1_LFInst_3_n2 , \Red_K2Inst_LFInst_2_LFInst_0_n2 ,
         \Red_K2Inst_LFInst_2_LFInst_1_n2 , \Red_K2Inst_LFInst_2_LFInst_2_n2 ,
         \Red_K2Inst_LFInst_2_LFInst_3_n2 , \Red_K2Inst_LFInst_3_LFInst_0_n2 ,
         \Red_K2Inst_LFInst_3_LFInst_1_n2 , \Red_K2Inst_LFInst_3_LFInst_2_n2 ,
         \Red_K2Inst_LFInst_3_LFInst_3_n2 , \Red_K2Inst_LFInst_4_LFInst_0_n2 ,
         \Red_K2Inst_LFInst_4_LFInst_1_n2 , \Red_K2Inst_LFInst_4_LFInst_2_n2 ,
         \Red_K2Inst_LFInst_4_LFInst_3_n2 , \Red_K2Inst_LFInst_5_LFInst_0_n2 ,
         \Red_K2Inst_LFInst_5_LFInst_1_n2 , \Red_K2Inst_LFInst_5_LFInst_2_n2 ,
         \Red_K2Inst_LFInst_5_LFInst_3_n2 , \Red_K2Inst_LFInst_6_LFInst_0_n2 ,
         \Red_K2Inst_LFInst_6_LFInst_1_n2 , \Red_K2Inst_LFInst_6_LFInst_2_n2 ,
         \Red_K2Inst_LFInst_6_LFInst_3_n2 , \Red_K2Inst_LFInst_7_LFInst_0_n2 ,
         \Red_K2Inst_LFInst_7_LFInst_1_n2 , \Red_K2Inst_LFInst_7_LFInst_2_n2 ,
         \Red_K2Inst_LFInst_7_LFInst_3_n2 , \Red_K2Inst_LFInst_8_LFInst_0_n2 ,
         \Red_K2Inst_LFInst_8_LFInst_1_n2 , \Red_K2Inst_LFInst_8_LFInst_2_n2 ,
         \Red_K2Inst_LFInst_8_LFInst_3_n2 , \Red_K2Inst_LFInst_9_LFInst_0_n2 ,
         \Red_K2Inst_LFInst_9_LFInst_1_n2 , \Red_K2Inst_LFInst_9_LFInst_2_n2 ,
         \Red_K2Inst_LFInst_9_LFInst_3_n2 , \Red_K2Inst_LFInst_10_LFInst_0_n2 ,
         \Red_K2Inst_LFInst_10_LFInst_1_n2 ,
         \Red_K2Inst_LFInst_10_LFInst_2_n2 ,
         \Red_K2Inst_LFInst_10_LFInst_3_n2 ,
         \Red_K2Inst_LFInst_11_LFInst_0_n2 ,
         \Red_K2Inst_LFInst_11_LFInst_1_n2 ,
         \Red_K2Inst_LFInst_11_LFInst_2_n2 ,
         \Red_K2Inst_LFInst_11_LFInst_3_n2 ,
         \Red_K2Inst_LFInst_12_LFInst_0_n2 ,
         \Red_K2Inst_LFInst_12_LFInst_1_n2 ,
         \Red_K2Inst_LFInst_12_LFInst_2_n2 ,
         \Red_K2Inst_LFInst_12_LFInst_3_n2 ,
         \Red_K2Inst_LFInst_13_LFInst_0_n2 ,
         \Red_K2Inst_LFInst_13_LFInst_1_n2 ,
         \Red_K2Inst_LFInst_13_LFInst_2_n2 ,
         \Red_K2Inst_LFInst_13_LFInst_3_n2 ,
         \Red_K2Inst_LFInst_14_LFInst_0_n2 ,
         \Red_K2Inst_LFInst_14_LFInst_1_n2 ,
         \Red_K2Inst_LFInst_14_LFInst_2_n2 ,
         \Red_K2Inst_LFInst_14_LFInst_3_n2 ,
         \Red_K2Inst_LFInst_15_LFInst_0_n2 ,
         \Red_K2Inst_LFInst_15_LFInst_1_n2 ,
         \Red_K2Inst_LFInst_15_LFInst_2_n2 ,
         \Red_K2Inst_LFInst_15_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_0_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_0_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_0_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_0_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_1_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_1_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_1_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_1_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_2_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_2_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_2_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_2_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_3_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_3_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_3_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_3_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_4_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_4_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_4_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_4_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_5_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_5_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_5_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_5_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_6_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_6_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_6_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_6_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_7_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_7_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_7_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_7_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_8_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_8_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_8_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_8_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_9_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_9_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_9_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_9_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_10_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_10_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_10_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_10_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_11_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_11_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_11_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_11_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_12_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_12_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_12_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_12_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_13_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_13_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_13_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_13_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_14_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_14_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_14_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_14_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_15_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_15_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_15_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_15_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_16_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_16_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_16_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_16_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_17_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_17_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_17_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_17_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_18_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_18_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_18_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_18_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_19_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_19_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_19_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_19_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_20_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_20_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_20_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_20_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_21_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_21_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_21_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_21_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_22_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_22_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_22_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_22_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_23_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_23_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_23_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_23_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_24_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_24_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_24_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_24_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_25_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_25_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_25_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_25_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_26_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_26_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_26_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_26_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_27_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_27_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_27_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_27_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_28_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_28_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_28_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_28_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_29_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_29_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_29_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_29_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_30_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_30_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_30_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_30_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_31_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_31_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_31_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_31_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_32_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_32_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_32_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_32_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_33_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_33_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_33_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_33_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_34_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_34_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_34_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_34_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_35_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_35_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_35_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_35_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_36_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_36_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_36_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_36_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_37_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_37_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_37_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_37_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_38_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_38_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_38_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_38_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_39_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_39_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_39_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_39_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_40_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_40_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_40_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_40_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_41_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_41_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_41_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_41_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_42_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_42_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_42_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_42_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_43_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_43_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_43_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_43_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_44_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_44_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_44_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_44_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_45_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_45_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_45_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_45_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_46_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_46_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_46_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_46_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_47_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_47_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_47_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_47_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_48_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_48_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_48_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_48_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_49_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_49_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_49_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_49_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_50_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_50_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_50_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_50_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_51_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_51_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_51_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_51_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_52_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_52_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_52_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_52_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_53_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_53_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_53_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_53_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_54_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_54_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_54_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_54_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_55_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_55_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_55_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_55_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_56_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_56_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_56_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_56_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_57_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_57_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_57_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_57_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_58_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_58_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_58_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_58_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_59_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_59_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_59_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_59_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_60_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_60_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_60_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_60_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_61_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_61_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_61_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_61_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_62_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_62_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_62_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_62_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_63_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_63_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_63_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_63_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_64_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_64_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_64_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_64_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_65_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_65_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_65_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_65_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_66_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_66_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_66_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_66_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_67_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_67_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_67_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_67_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_68_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_68_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_68_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_68_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_69_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_69_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_69_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_69_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_70_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_70_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_70_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_70_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_71_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_71_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_71_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_71_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_72_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_72_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_72_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_72_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_73_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_73_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_73_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_73_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_74_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_74_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_74_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_74_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_75_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_75_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_75_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_75_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_76_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_76_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_76_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_76_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_77_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_77_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_77_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_77_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_78_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_78_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_78_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_78_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_79_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_79_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_79_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_79_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_80_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_80_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_80_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_80_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_81_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_81_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_81_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_81_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_82_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_82_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_82_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_82_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_83_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_83_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_83_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_83_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_84_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_84_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_84_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_84_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_85_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_85_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_85_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_85_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_86_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_86_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_86_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_86_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_87_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_87_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_87_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_87_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_88_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_88_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_88_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_88_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_89_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_89_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_89_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_89_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_90_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_90_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_90_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_90_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_91_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_91_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_91_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_91_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_92_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_92_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_92_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_92_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_93_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_93_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_93_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_93_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_94_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_94_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_94_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_94_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_95_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_95_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_95_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_95_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_96_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_96_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_96_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_96_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_97_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_97_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_97_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_97_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_98_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_98_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_98_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_98_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_99_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_99_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_99_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_99_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_100_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_100_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_100_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_100_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_101_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_101_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_101_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_101_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_102_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_102_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_102_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_102_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_103_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_103_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_103_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_103_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_104_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_104_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_104_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_104_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_105_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_105_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_105_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_105_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_106_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_106_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_106_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_106_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_107_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_107_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_107_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_107_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_108_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_108_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_108_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_108_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_109_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_109_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_109_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_109_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_110_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_110_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_110_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_110_LFInst_3_n2 ,
         \Red_ToCheckInst_LFInst_111_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_111_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_111_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_111_LFInst_3_n2 , \Check1_CheckInst_0_n222 ,
         \Check1_CheckInst_0_n221 , \Check1_CheckInst_0_n220 ,
         \Check1_CheckInst_0_n219 , \Check1_CheckInst_0_n218 ,
         \Check1_CheckInst_0_n217 , \Check1_CheckInst_0_n216 ,
         \Check1_CheckInst_0_n215 , \Check1_CheckInst_0_n214 ,
         \Check1_CheckInst_0_n213 , \Check1_CheckInst_0_n212 ,
         \Check1_CheckInst_0_n211 , \Check1_CheckInst_0_n210 ,
         \Check1_CheckInst_0_n209 , \Check1_CheckInst_0_n208 ,
         \Check1_CheckInst_0_n207 , \Check1_CheckInst_0_n206 ,
         \Check1_CheckInst_0_n205 , \Check1_CheckInst_0_n204 ,
         \Check1_CheckInst_0_n203 , \Check1_CheckInst_0_n202 ,
         \Check1_CheckInst_0_n201 , \Check1_CheckInst_0_n200 ,
         \Check1_CheckInst_0_n199 , \Check1_CheckInst_0_n198 ,
         \Check1_CheckInst_0_n197 , \Check1_CheckInst_0_n196 ,
         \Check1_CheckInst_0_n195 , \Check1_CheckInst_0_n194 ,
         \Check1_CheckInst_0_n193 , \Check1_CheckInst_0_n192 ,
         \Check1_CheckInst_0_n191 , \Check1_CheckInst_0_n190 ,
         \Check1_CheckInst_0_n189 , \Check1_CheckInst_0_n188 ,
         \Check1_CheckInst_0_n187 , \Check1_CheckInst_0_n186 ,
         \Check1_CheckInst_0_n185 , \Check1_CheckInst_0_n184 ,
         \Check1_CheckInst_0_n183 , \Check1_CheckInst_0_n182 ,
         \Check1_CheckInst_0_n181 , \Check1_CheckInst_0_n180 ,
         \Check1_CheckInst_0_n179 , \Check1_CheckInst_0_n178 ,
         \Check1_CheckInst_0_n177 , \Check1_CheckInst_0_n176 ,
         \Check1_CheckInst_0_n175 , \Check1_CheckInst_0_n174 ,
         \Check1_CheckInst_0_n173 , \Check1_CheckInst_0_n172 ,
         \Check1_CheckInst_0_n171 , \Check1_CheckInst_0_n170 ,
         \Check1_CheckInst_0_n169 , \Check1_CheckInst_0_n168 ,
         \Check1_CheckInst_0_n167 , \Check1_CheckInst_0_n166 ,
         \Check1_CheckInst_0_n165 , \Check1_CheckInst_0_n164 ,
         \Check1_CheckInst_0_n163 , \Check1_CheckInst_0_n162 ,
         \Check1_CheckInst_0_n161 , \Check1_CheckInst_0_n160 ,
         \Check1_CheckInst_0_n159 , \Check1_CheckInst_0_n158 ,
         \Check1_CheckInst_0_n157 , \Check1_CheckInst_0_n156 ,
         \Check1_CheckInst_0_n155 , \Check1_CheckInst_0_n154 ,
         \Check1_CheckInst_0_n153 , \Check1_CheckInst_0_n152 ,
         \Check1_CheckInst_0_n151 , \Check1_CheckInst_0_n150 ,
         \Check1_CheckInst_0_n149 , \Check1_CheckInst_0_n148 ,
         \Check1_CheckInst_0_n147 , \Check1_CheckInst_0_n146 ,
         \Check1_CheckInst_0_n145 , \Check1_CheckInst_0_n144 ,
         \Check1_CheckInst_0_n143 , \Check1_CheckInst_0_n142 ,
         \Check1_CheckInst_0_n141 , \Check1_CheckInst_0_n140 ,
         \Check1_CheckInst_0_n139 , \Check1_CheckInst_0_n138 ,
         \Check1_CheckInst_0_n137 , \Check1_CheckInst_0_n136 ,
         \Check1_CheckInst_0_n135 , \Check1_CheckInst_0_n134 ,
         \Check1_CheckInst_0_n133 , \Check1_CheckInst_0_n132 ,
         \Check1_CheckInst_0_n131 , \Check1_CheckInst_0_n130 ,
         \Check1_CheckInst_0_n129 , \Check1_CheckInst_0_n128 ,
         \Check1_CheckInst_0_n127 , \Check1_CheckInst_0_n126 ,
         \Check1_CheckInst_0_n125 , \Check1_CheckInst_0_n124 ,
         \Check1_CheckInst_0_n123 , \Check1_CheckInst_0_n122 ,
         \Check1_CheckInst_0_n121 , \Check1_CheckInst_0_n120 ,
         \Check1_CheckInst_0_n119 , \Check1_CheckInst_0_n118 ,
         \Check1_CheckInst_0_n117 , \Check1_CheckInst_0_n116 ,
         \Check1_CheckInst_0_n115 , \Check1_CheckInst_0_n114 ,
         \Check1_CheckInst_0_n113 , \Check1_CheckInst_0_n112 ,
         \Check1_CheckInst_0_n111 , \Check1_CheckInst_0_n110 ,
         \Check1_CheckInst_0_n109 , \Check1_CheckInst_0_n108 ,
         \Check1_CheckInst_0_n107 , \Check1_CheckInst_0_n106 ,
         \Check1_CheckInst_0_n105 , \Check1_CheckInst_0_n104 ,
         \Check1_CheckInst_0_n103 , \Check1_CheckInst_0_n102 ,
         \Check1_CheckInst_0_n101 , \Check1_CheckInst_0_n100 ,
         \Check1_CheckInst_0_n99 , \Check1_CheckInst_0_n98 ,
         \Check1_CheckInst_0_n97 , \Check1_CheckInst_0_n96 ,
         \Check1_CheckInst_0_n95 , \Check1_CheckInst_0_n94 ,
         \Check1_CheckInst_0_n93 , \Check1_CheckInst_0_n92 ,
         \Check1_CheckInst_0_n91 , \Check1_CheckInst_0_n90 ,
         \Check1_CheckInst_0_n89 , \Check1_CheckInst_0_n88 ,
         \Check1_CheckInst_0_n87 , \Check1_CheckInst_0_n86 ,
         \Check1_CheckInst_0_n85 , \Check1_CheckInst_0_n84 ,
         \Check1_CheckInst_0_n83 , \Check1_CheckInst_0_n82 ,
         \Check1_CheckInst_0_n81 , \Check1_CheckInst_0_n80 ,
         \Check1_CheckInst_0_n79 , \Check1_CheckInst_0_n78 ,
         \Check1_CheckInst_0_n77 , \Check1_CheckInst_0_n76 ,
         \Check1_CheckInst_0_n75 , \Check1_CheckInst_0_n74 ,
         \Check1_CheckInst_0_n73 , \Check1_CheckInst_0_n72 ,
         \Check1_CheckInst_0_n71 , \Check1_CheckInst_0_n70 ,
         \Check1_CheckInst_0_n69 , \Check1_CheckInst_0_n68 ,
         \Check1_CheckInst_0_n67 , \Check1_CheckInst_0_n66 ,
         \Check1_CheckInst_0_n65 , \Check1_CheckInst_0_n64 ,
         \Check1_CheckInst_0_n63 , \Check1_CheckInst_0_n62 ,
         \Check1_CheckInst_0_n61 , \Check1_CheckInst_0_n60 ,
         \Check1_CheckInst_0_n59 , \Check1_CheckInst_0_n58 ,
         \Check1_CheckInst_0_n57 , \Check1_CheckInst_0_n56 ,
         \Check1_CheckInst_0_n55 , \Check1_CheckInst_0_n54 ,
         \Check1_CheckInst_0_n53 , \Check1_CheckInst_0_n52 ,
         \Check1_CheckInst_0_n51 , \Check1_CheckInst_0_n50 ,
         \Check1_CheckInst_0_n49 , \Check1_CheckInst_0_n48 ,
         \Check1_CheckInst_0_n47 , \Check1_CheckInst_0_n46 ,
         \Check1_CheckInst_0_n45 , \Check1_CheckInst_0_n44 ,
         \Check1_CheckInst_0_n43 , \Check1_CheckInst_0_n42 ,
         \Check1_CheckInst_0_n41 , \Check1_CheckInst_0_n40 ,
         \Check1_CheckInst_0_n39 , \Check1_CheckInst_0_n38 ,
         \Check1_CheckInst_0_n37 , \Check1_CheckInst_0_n36 ,
         \Check1_CheckInst_0_n35 , \Check1_CheckInst_0_n34 ,
         \Check1_CheckInst_0_n33 , \Check1_CheckInst_0_n32 ,
         \Check1_CheckInst_0_n31 , \Check1_CheckInst_0_n30 ,
         \Check1_CheckInst_0_n29 , \Check1_CheckInst_0_n28 ,
         \Check1_CheckInst_0_n27 , \Check1_CheckInst_0_n26 ,
         \Check1_CheckInst_0_n25 , \Check1_CheckInst_0_n24 ,
         \Check1_CheckInst_0_n23 , \Check1_CheckInst_0_n22 ,
         \Check1_CheckInst_0_n21 , \Check1_CheckInst_0_n20 ,
         \Check1_CheckInst_0_n19 , \Check1_CheckInst_0_n18 ,
         \Check1_CheckInst_0_n17 , \Check1_CheckInst_0_n16 ,
         \Check1_CheckInst_0_n15 , \Check1_CheckInst_0_n14 ,
         \Check1_CheckInst_0_n13 , \Check1_CheckInst_0_n12 ,
         \Check1_CheckInst_0_n11 , \Check1_CheckInst_0_n10 ,
         \Check1_CheckInst_0_n9 , \Check1_CheckInst_0_n8 ,
         \Check1_CheckInst_0_n7 , \Check1_CheckInst_0_n6 ,
         \Check1_CheckInst_0_n5 , \Check1_CheckInst_0_n4 ,
         \Check1_CheckInst_0_n3 , \Check1_CheckInst_0_n2 ,
         \Check1_CheckInst_0_n1 , \Check1_CheckInst_1_n224 ,
         \Check1_CheckInst_1_n223 , \Check1_CheckInst_1_n222 ,
         \Check1_CheckInst_1_n221 , \Check1_CheckInst_1_n220 ,
         \Check1_CheckInst_1_n219 , \Check1_CheckInst_1_n218 ,
         \Check1_CheckInst_1_n217 , \Check1_CheckInst_1_n216 ,
         \Check1_CheckInst_1_n215 , \Check1_CheckInst_1_n214 ,
         \Check1_CheckInst_1_n213 , \Check1_CheckInst_1_n212 ,
         \Check1_CheckInst_1_n211 , \Check1_CheckInst_1_n210 ,
         \Check1_CheckInst_1_n209 , \Check1_CheckInst_1_n208 ,
         \Check1_CheckInst_1_n207 , \Check1_CheckInst_1_n206 ,
         \Check1_CheckInst_1_n205 , \Check1_CheckInst_1_n204 ,
         \Check1_CheckInst_1_n203 , \Check1_CheckInst_1_n202 ,
         \Check1_CheckInst_1_n201 , \Check1_CheckInst_1_n200 ,
         \Check1_CheckInst_1_n199 , \Check1_CheckInst_1_n198 ,
         \Check1_CheckInst_1_n197 , \Check1_CheckInst_1_n196 ,
         \Check1_CheckInst_1_n195 , \Check1_CheckInst_1_n194 ,
         \Check1_CheckInst_1_n193 , \Check1_CheckInst_1_n192 ,
         \Check1_CheckInst_1_n191 , \Check1_CheckInst_1_n190 ,
         \Check1_CheckInst_1_n189 , \Check1_CheckInst_1_n188 ,
         \Check1_CheckInst_1_n187 , \Check1_CheckInst_1_n186 ,
         \Check1_CheckInst_1_n185 , \Check1_CheckInst_1_n184 ,
         \Check1_CheckInst_1_n183 , \Check1_CheckInst_1_n182 ,
         \Check1_CheckInst_1_n181 , \Check1_CheckInst_1_n180 ,
         \Check1_CheckInst_1_n179 , \Check1_CheckInst_1_n178 ,
         \Check1_CheckInst_1_n177 , \Check1_CheckInst_1_n176 ,
         \Check1_CheckInst_1_n175 , \Check1_CheckInst_1_n174 ,
         \Check1_CheckInst_1_n173 , \Check1_CheckInst_1_n172 ,
         \Check1_CheckInst_1_n171 , \Check1_CheckInst_1_n170 ,
         \Check1_CheckInst_1_n169 , \Check1_CheckInst_1_n168 ,
         \Check1_CheckInst_1_n167 , \Check1_CheckInst_1_n166 ,
         \Check1_CheckInst_1_n165 , \Check1_CheckInst_1_n164 ,
         \Check1_CheckInst_1_n163 , \Check1_CheckInst_1_n162 ,
         \Check1_CheckInst_1_n161 , \Check1_CheckInst_1_n160 ,
         \Check1_CheckInst_1_n159 , \Check1_CheckInst_1_n158 ,
         \Check1_CheckInst_1_n157 , \Check1_CheckInst_1_n156 ,
         \Check1_CheckInst_1_n155 , \Check1_CheckInst_1_n154 ,
         \Check1_CheckInst_1_n153 , \Check1_CheckInst_1_n152 ,
         \Check1_CheckInst_1_n151 , \Check1_CheckInst_1_n150 ,
         \Check1_CheckInst_1_n149 , \Check1_CheckInst_1_n148 ,
         \Check1_CheckInst_1_n147 , \Check1_CheckInst_1_n146 ,
         \Check1_CheckInst_1_n145 , \Check1_CheckInst_1_n144 ,
         \Check1_CheckInst_1_n143 , \Check1_CheckInst_1_n142 ,
         \Check1_CheckInst_1_n141 , \Check1_CheckInst_1_n140 ,
         \Check1_CheckInst_1_n139 , \Check1_CheckInst_1_n138 ,
         \Check1_CheckInst_1_n137 , \Check1_CheckInst_1_n136 ,
         \Check1_CheckInst_1_n135 , \Check1_CheckInst_1_n134 ,
         \Check1_CheckInst_1_n133 , \Check1_CheckInst_1_n132 ,
         \Check1_CheckInst_1_n131 , \Check1_CheckInst_1_n130 ,
         \Check1_CheckInst_1_n129 , \Check1_CheckInst_1_n128 ,
         \Check1_CheckInst_1_n127 , \Check1_CheckInst_1_n126 ,
         \Check1_CheckInst_1_n125 , \Check1_CheckInst_1_n124 ,
         \Check1_CheckInst_1_n123 , \Check1_CheckInst_1_n122 ,
         \Check1_CheckInst_1_n121 , \Check1_CheckInst_1_n120 ,
         \Check1_CheckInst_1_n119 , \Check1_CheckInst_1_n118 ,
         \Check1_CheckInst_1_n117 , \Check1_CheckInst_1_n116 ,
         \Check1_CheckInst_1_n115 , \Check1_CheckInst_1_n114 ,
         \Check1_CheckInst_1_n113 , \Check1_CheckInst_1_n112 ,
         \Check1_CheckInst_1_n111 , \Check1_CheckInst_1_n110 ,
         \Check1_CheckInst_1_n109 , \Check1_CheckInst_1_n108 ,
         \Check1_CheckInst_1_n107 , \Check1_CheckInst_1_n106 ,
         \Check1_CheckInst_1_n105 , \Check1_CheckInst_1_n104 ,
         \Check1_CheckInst_1_n103 , \Check1_CheckInst_1_n102 ,
         \Check1_CheckInst_1_n101 , \Check1_CheckInst_1_n100 ,
         \Check1_CheckInst_1_n99 , \Check1_CheckInst_1_n98 ,
         \Check1_CheckInst_1_n97 , \Check1_CheckInst_1_n96 ,
         \Check1_CheckInst_1_n95 , \Check1_CheckInst_1_n94 ,
         \Check1_CheckInst_1_n93 , \Check1_CheckInst_1_n92 ,
         \Check1_CheckInst_1_n91 , \Check1_CheckInst_1_n90 ,
         \Check1_CheckInst_1_n89 , \Check1_CheckInst_1_n88 ,
         \Check1_CheckInst_1_n87 , \Check1_CheckInst_1_n86 ,
         \Check1_CheckInst_1_n85 , \Check1_CheckInst_1_n84 ,
         \Check1_CheckInst_1_n83 , \Check1_CheckInst_1_n82 ,
         \Check1_CheckInst_1_n81 , \Check1_CheckInst_1_n80 ,
         \Check1_CheckInst_1_n79 , \Check1_CheckInst_1_n78 ,
         \Check1_CheckInst_1_n77 , \Check1_CheckInst_1_n76 ,
         \Check1_CheckInst_1_n75 , \Check1_CheckInst_1_n74 ,
         \Check1_CheckInst_1_n73 , \Check1_CheckInst_1_n72 ,
         \Check1_CheckInst_1_n71 , \Check1_CheckInst_1_n70 ,
         \Check1_CheckInst_1_n69 , \Check1_CheckInst_1_n68 ,
         \Check1_CheckInst_1_n67 , \Check1_CheckInst_1_n66 ,
         \Check1_CheckInst_1_n65 , \Check1_CheckInst_1_n64 ,
         \Check1_CheckInst_1_n63 , \Check1_CheckInst_1_n62 ,
         \Check1_CheckInst_1_n61 , \Check1_CheckInst_1_n60 ,
         \Check1_CheckInst_1_n59 , \Check1_CheckInst_1_n58 ,
         \Check1_CheckInst_1_n57 , \Check1_CheckInst_1_n56 ,
         \Check1_CheckInst_1_n55 , \Check1_CheckInst_1_n54 ,
         \Check1_CheckInst_1_n53 , \Check1_CheckInst_1_n52 ,
         \Check1_CheckInst_1_n51 , \Check1_CheckInst_1_n50 ,
         \Check1_CheckInst_1_n49 , \Check1_CheckInst_1_n48 ,
         \Check1_CheckInst_1_n47 , \Check1_CheckInst_1_n46 ,
         \Check1_CheckInst_1_n45 , \Check1_CheckInst_1_n44 ,
         \Check1_CheckInst_1_n43 , \Check1_CheckInst_1_n42 ,
         \Check1_CheckInst_1_n41 , \Check1_CheckInst_1_n40 ,
         \Check1_CheckInst_1_n39 , \Check1_CheckInst_1_n38 ,
         \Check1_CheckInst_1_n37 , \Check1_CheckInst_1_n36 ,
         \Check1_CheckInst_1_n35 , \Check1_CheckInst_1_n34 ,
         \Check1_CheckInst_1_n33 , \Check1_CheckInst_1_n32 ,
         \Check1_CheckInst_1_n31 , \Check1_CheckInst_1_n30 ,
         \Check1_CheckInst_1_n29 , \Check1_CheckInst_1_n28 ,
         \Check1_CheckInst_1_n27 , \Check1_CheckInst_1_n26 ,
         \Check1_CheckInst_1_n25 , \Check1_CheckInst_1_n24 ,
         \Check1_CheckInst_1_n23 , \Check1_CheckInst_1_n22 ,
         \Check1_CheckInst_1_n21 , \Check1_CheckInst_1_n20 ,
         \Check1_CheckInst_1_n19 , \Check1_CheckInst_1_n18 ,
         \Check1_CheckInst_1_n17 , \Check1_CheckInst_1_n16 ,
         \Check1_CheckInst_1_n15 , \Check1_CheckInst_1_n14 ,
         \Check1_CheckInst_1_n13 , \Check1_CheckInst_1_n12 ,
         \Check1_CheckInst_1_n11 , \Check1_CheckInst_1_n10 ,
         \Check1_CheckInst_1_n9 , \Check1_CheckInst_1_n8 ,
         \Check1_CheckInst_1_n7 , \Check1_CheckInst_1_n6 ,
         \Check1_CheckInst_1_n5 , \Check1_CheckInst_1_n4 ,
         \Check1_CheckInst_1_n3 , \Check1_CheckInst_2_n224 ,
         \Check1_CheckInst_2_n223 , \Check1_CheckInst_2_n222 ,
         \Check1_CheckInst_2_n221 , \Check1_CheckInst_2_n220 ,
         \Check1_CheckInst_2_n219 , \Check1_CheckInst_2_n218 ,
         \Check1_CheckInst_2_n217 , \Check1_CheckInst_2_n216 ,
         \Check1_CheckInst_2_n215 , \Check1_CheckInst_2_n214 ,
         \Check1_CheckInst_2_n213 , \Check1_CheckInst_2_n212 ,
         \Check1_CheckInst_2_n211 , \Check1_CheckInst_2_n210 ,
         \Check1_CheckInst_2_n209 , \Check1_CheckInst_2_n208 ,
         \Check1_CheckInst_2_n207 , \Check1_CheckInst_2_n206 ,
         \Check1_CheckInst_2_n205 , \Check1_CheckInst_2_n204 ,
         \Check1_CheckInst_2_n203 , \Check1_CheckInst_2_n202 ,
         \Check1_CheckInst_2_n201 , \Check1_CheckInst_2_n200 ,
         \Check1_CheckInst_2_n199 , \Check1_CheckInst_2_n198 ,
         \Check1_CheckInst_2_n197 , \Check1_CheckInst_2_n196 ,
         \Check1_CheckInst_2_n195 , \Check1_CheckInst_2_n194 ,
         \Check1_CheckInst_2_n193 , \Check1_CheckInst_2_n192 ,
         \Check1_CheckInst_2_n191 , \Check1_CheckInst_2_n190 ,
         \Check1_CheckInst_2_n189 , \Check1_CheckInst_2_n188 ,
         \Check1_CheckInst_2_n187 , \Check1_CheckInst_2_n186 ,
         \Check1_CheckInst_2_n185 , \Check1_CheckInst_2_n184 ,
         \Check1_CheckInst_2_n183 , \Check1_CheckInst_2_n182 ,
         \Check1_CheckInst_2_n181 , \Check1_CheckInst_2_n180 ,
         \Check1_CheckInst_2_n179 , \Check1_CheckInst_2_n178 ,
         \Check1_CheckInst_2_n177 , \Check1_CheckInst_2_n176 ,
         \Check1_CheckInst_2_n175 , \Check1_CheckInst_2_n174 ,
         \Check1_CheckInst_2_n173 , \Check1_CheckInst_2_n172 ,
         \Check1_CheckInst_2_n171 , \Check1_CheckInst_2_n170 ,
         \Check1_CheckInst_2_n169 , \Check1_CheckInst_2_n168 ,
         \Check1_CheckInst_2_n167 , \Check1_CheckInst_2_n166 ,
         \Check1_CheckInst_2_n165 , \Check1_CheckInst_2_n164 ,
         \Check1_CheckInst_2_n163 , \Check1_CheckInst_2_n162 ,
         \Check1_CheckInst_2_n161 , \Check1_CheckInst_2_n160 ,
         \Check1_CheckInst_2_n159 , \Check1_CheckInst_2_n158 ,
         \Check1_CheckInst_2_n157 , \Check1_CheckInst_2_n156 ,
         \Check1_CheckInst_2_n155 , \Check1_CheckInst_2_n154 ,
         \Check1_CheckInst_2_n153 , \Check1_CheckInst_2_n152 ,
         \Check1_CheckInst_2_n151 , \Check1_CheckInst_2_n150 ,
         \Check1_CheckInst_2_n149 , \Check1_CheckInst_2_n148 ,
         \Check1_CheckInst_2_n147 , \Check1_CheckInst_2_n146 ,
         \Check1_CheckInst_2_n145 , \Check1_CheckInst_2_n144 ,
         \Check1_CheckInst_2_n143 , \Check1_CheckInst_2_n142 ,
         \Check1_CheckInst_2_n141 , \Check1_CheckInst_2_n140 ,
         \Check1_CheckInst_2_n139 , \Check1_CheckInst_2_n138 ,
         \Check1_CheckInst_2_n137 , \Check1_CheckInst_2_n136 ,
         \Check1_CheckInst_2_n135 , \Check1_CheckInst_2_n134 ,
         \Check1_CheckInst_2_n133 , \Check1_CheckInst_2_n132 ,
         \Check1_CheckInst_2_n131 , \Check1_CheckInst_2_n130 ,
         \Check1_CheckInst_2_n129 , \Check1_CheckInst_2_n128 ,
         \Check1_CheckInst_2_n127 , \Check1_CheckInst_2_n126 ,
         \Check1_CheckInst_2_n125 , \Check1_CheckInst_2_n124 ,
         \Check1_CheckInst_2_n123 , \Check1_CheckInst_2_n122 ,
         \Check1_CheckInst_2_n121 , \Check1_CheckInst_2_n120 ,
         \Check1_CheckInst_2_n119 , \Check1_CheckInst_2_n118 ,
         \Check1_CheckInst_2_n117 , \Check1_CheckInst_2_n116 ,
         \Check1_CheckInst_2_n115 , \Check1_CheckInst_2_n114 ,
         \Check1_CheckInst_2_n113 , \Check1_CheckInst_2_n112 ,
         \Check1_CheckInst_2_n111 , \Check1_CheckInst_2_n110 ,
         \Check1_CheckInst_2_n109 , \Check1_CheckInst_2_n108 ,
         \Check1_CheckInst_2_n107 , \Check1_CheckInst_2_n106 ,
         \Check1_CheckInst_2_n105 , \Check1_CheckInst_2_n104 ,
         \Check1_CheckInst_2_n103 , \Check1_CheckInst_2_n102 ,
         \Check1_CheckInst_2_n101 , \Check1_CheckInst_2_n100 ,
         \Check1_CheckInst_2_n99 , \Check1_CheckInst_2_n98 ,
         \Check1_CheckInst_2_n97 , \Check1_CheckInst_2_n96 ,
         \Check1_CheckInst_2_n95 , \Check1_CheckInst_2_n94 ,
         \Check1_CheckInst_2_n93 , \Check1_CheckInst_2_n92 ,
         \Check1_CheckInst_2_n91 , \Check1_CheckInst_2_n90 ,
         \Check1_CheckInst_2_n89 , \Check1_CheckInst_2_n88 ,
         \Check1_CheckInst_2_n87 , \Check1_CheckInst_2_n86 ,
         \Check1_CheckInst_2_n85 , \Check1_CheckInst_2_n84 ,
         \Check1_CheckInst_2_n83 , \Check1_CheckInst_2_n82 ,
         \Check1_CheckInst_2_n81 , \Check1_CheckInst_2_n80 ,
         \Check1_CheckInst_2_n79 , \Check1_CheckInst_2_n78 ,
         \Check1_CheckInst_2_n77 , \Check1_CheckInst_2_n76 ,
         \Check1_CheckInst_2_n75 , \Check1_CheckInst_2_n74 ,
         \Check1_CheckInst_2_n73 , \Check1_CheckInst_2_n72 ,
         \Check1_CheckInst_2_n71 , \Check1_CheckInst_2_n70 ,
         \Check1_CheckInst_2_n69 , \Check1_CheckInst_2_n68 ,
         \Check1_CheckInst_2_n67 , \Check1_CheckInst_2_n66 ,
         \Check1_CheckInst_2_n65 , \Check1_CheckInst_2_n64 ,
         \Check1_CheckInst_2_n63 , \Check1_CheckInst_2_n62 ,
         \Check1_CheckInst_2_n61 , \Check1_CheckInst_2_n60 ,
         \Check1_CheckInst_2_n59 , \Check1_CheckInst_2_n58 ,
         \Check1_CheckInst_2_n57 , \Check1_CheckInst_2_n56 ,
         \Check1_CheckInst_2_n55 , \Check1_CheckInst_2_n54 ,
         \Check1_CheckInst_2_n53 , \Check1_CheckInst_2_n52 ,
         \Check1_CheckInst_2_n51 , \Check1_CheckInst_2_n50 ,
         \Check1_CheckInst_2_n49 , \Check1_CheckInst_2_n48 ,
         \Check1_CheckInst_2_n47 , \Check1_CheckInst_2_n46 ,
         \Check1_CheckInst_2_n45 , \Check1_CheckInst_2_n44 ,
         \Check1_CheckInst_2_n43 , \Check1_CheckInst_2_n42 ,
         \Check1_CheckInst_2_n41 , \Check1_CheckInst_2_n40 ,
         \Check1_CheckInst_2_n39 , \Check1_CheckInst_2_n38 ,
         \Check1_CheckInst_2_n37 , \Check1_CheckInst_2_n36 ,
         \Check1_CheckInst_2_n35 , \Check1_CheckInst_2_n34 ,
         \Check1_CheckInst_2_n33 , \Check1_CheckInst_2_n32 ,
         \Check1_CheckInst_2_n31 , \Check1_CheckInst_2_n30 ,
         \Check1_CheckInst_2_n29 , \Check1_CheckInst_2_n28 ,
         \Check1_CheckInst_2_n27 , \Check1_CheckInst_2_n26 ,
         \Check1_CheckInst_2_n25 , \Check1_CheckInst_2_n24 ,
         \Check1_CheckInst_2_n23 , \Check1_CheckInst_2_n22 ,
         \Check1_CheckInst_2_n21 , \Check1_CheckInst_2_n20 ,
         \Check1_CheckInst_2_n19 , \Check1_CheckInst_2_n18 ,
         \Check1_CheckInst_2_n17 , \Check1_CheckInst_2_n16 ,
         \Check1_CheckInst_2_n15 , \Check1_CheckInst_2_n14 ,
         \Check1_CheckInst_2_n13 , \Check1_CheckInst_2_n12 ,
         \Check1_CheckInst_2_n11 , \Check1_CheckInst_2_n10 ,
         \Check1_CheckInst_2_n9 , \Check1_CheckInst_2_n8 ,
         \Check1_CheckInst_2_n7 , \Check1_CheckInst_2_n6 ,
         \Check1_CheckInst_2_n5 , \Check1_CheckInst_2_n4 ,
         \Check1_CheckInst_2_n3 , \Check1_CheckInst_3_n224 ,
         \Check1_CheckInst_3_n223 , \Check1_CheckInst_3_n222 ,
         \Check1_CheckInst_3_n221 , \Check1_CheckInst_3_n220 ,
         \Check1_CheckInst_3_n219 , \Check1_CheckInst_3_n218 ,
         \Check1_CheckInst_3_n217 , \Check1_CheckInst_3_n216 ,
         \Check1_CheckInst_3_n215 , \Check1_CheckInst_3_n214 ,
         \Check1_CheckInst_3_n213 , \Check1_CheckInst_3_n212 ,
         \Check1_CheckInst_3_n211 , \Check1_CheckInst_3_n210 ,
         \Check1_CheckInst_3_n209 , \Check1_CheckInst_3_n208 ,
         \Check1_CheckInst_3_n207 , \Check1_CheckInst_3_n206 ,
         \Check1_CheckInst_3_n205 , \Check1_CheckInst_3_n204 ,
         \Check1_CheckInst_3_n203 , \Check1_CheckInst_3_n202 ,
         \Check1_CheckInst_3_n201 , \Check1_CheckInst_3_n200 ,
         \Check1_CheckInst_3_n199 , \Check1_CheckInst_3_n198 ,
         \Check1_CheckInst_3_n197 , \Check1_CheckInst_3_n196 ,
         \Check1_CheckInst_3_n195 , \Check1_CheckInst_3_n194 ,
         \Check1_CheckInst_3_n193 , \Check1_CheckInst_3_n192 ,
         \Check1_CheckInst_3_n191 , \Check1_CheckInst_3_n190 ,
         \Check1_CheckInst_3_n189 , \Check1_CheckInst_3_n188 ,
         \Check1_CheckInst_3_n187 , \Check1_CheckInst_3_n186 ,
         \Check1_CheckInst_3_n185 , \Check1_CheckInst_3_n184 ,
         \Check1_CheckInst_3_n183 , \Check1_CheckInst_3_n182 ,
         \Check1_CheckInst_3_n181 , \Check1_CheckInst_3_n180 ,
         \Check1_CheckInst_3_n179 , \Check1_CheckInst_3_n178 ,
         \Check1_CheckInst_3_n177 , \Check1_CheckInst_3_n176 ,
         \Check1_CheckInst_3_n175 , \Check1_CheckInst_3_n174 ,
         \Check1_CheckInst_3_n173 , \Check1_CheckInst_3_n172 ,
         \Check1_CheckInst_3_n171 , \Check1_CheckInst_3_n170 ,
         \Check1_CheckInst_3_n169 , \Check1_CheckInst_3_n168 ,
         \Check1_CheckInst_3_n167 , \Check1_CheckInst_3_n166 ,
         \Check1_CheckInst_3_n165 , \Check1_CheckInst_3_n164 ,
         \Check1_CheckInst_3_n163 , \Check1_CheckInst_3_n162 ,
         \Check1_CheckInst_3_n161 , \Check1_CheckInst_3_n160 ,
         \Check1_CheckInst_3_n159 , \Check1_CheckInst_3_n158 ,
         \Check1_CheckInst_3_n157 , \Check1_CheckInst_3_n156 ,
         \Check1_CheckInst_3_n155 , \Check1_CheckInst_3_n154 ,
         \Check1_CheckInst_3_n153 , \Check1_CheckInst_3_n152 ,
         \Check1_CheckInst_3_n151 , \Check1_CheckInst_3_n150 ,
         \Check1_CheckInst_3_n149 , \Check1_CheckInst_3_n148 ,
         \Check1_CheckInst_3_n147 , \Check1_CheckInst_3_n146 ,
         \Check1_CheckInst_3_n145 , \Check1_CheckInst_3_n144 ,
         \Check1_CheckInst_3_n143 , \Check1_CheckInst_3_n142 ,
         \Check1_CheckInst_3_n141 , \Check1_CheckInst_3_n140 ,
         \Check1_CheckInst_3_n139 , \Check1_CheckInst_3_n138 ,
         \Check1_CheckInst_3_n137 , \Check1_CheckInst_3_n136 ,
         \Check1_CheckInst_3_n135 , \Check1_CheckInst_3_n134 ,
         \Check1_CheckInst_3_n133 , \Check1_CheckInst_3_n132 ,
         \Check1_CheckInst_3_n131 , \Check1_CheckInst_3_n130 ,
         \Check1_CheckInst_3_n129 , \Check1_CheckInst_3_n128 ,
         \Check1_CheckInst_3_n127 , \Check1_CheckInst_3_n126 ,
         \Check1_CheckInst_3_n125 , \Check1_CheckInst_3_n124 ,
         \Check1_CheckInst_3_n123 , \Check1_CheckInst_3_n122 ,
         \Check1_CheckInst_3_n121 , \Check1_CheckInst_3_n120 ,
         \Check1_CheckInst_3_n119 , \Check1_CheckInst_3_n118 ,
         \Check1_CheckInst_3_n117 , \Check1_CheckInst_3_n116 ,
         \Check1_CheckInst_3_n115 , \Check1_CheckInst_3_n114 ,
         \Check1_CheckInst_3_n113 , \Check1_CheckInst_3_n112 ,
         \Check1_CheckInst_3_n111 , \Check1_CheckInst_3_n110 ,
         \Check1_CheckInst_3_n109 , \Check1_CheckInst_3_n108 ,
         \Check1_CheckInst_3_n107 , \Check1_CheckInst_3_n106 ,
         \Check1_CheckInst_3_n105 , \Check1_CheckInst_3_n104 ,
         \Check1_CheckInst_3_n103 , \Check1_CheckInst_3_n102 ,
         \Check1_CheckInst_3_n101 , \Check1_CheckInst_3_n100 ,
         \Check1_CheckInst_3_n99 , \Check1_CheckInst_3_n98 ,
         \Check1_CheckInst_3_n97 , \Check1_CheckInst_3_n96 ,
         \Check1_CheckInst_3_n95 , \Check1_CheckInst_3_n94 ,
         \Check1_CheckInst_3_n93 , \Check1_CheckInst_3_n92 ,
         \Check1_CheckInst_3_n91 , \Check1_CheckInst_3_n90 ,
         \Check1_CheckInst_3_n89 , \Check1_CheckInst_3_n88 ,
         \Check1_CheckInst_3_n87 , \Check1_CheckInst_3_n86 ,
         \Check1_CheckInst_3_n85 , \Check1_CheckInst_3_n84 ,
         \Check1_CheckInst_3_n83 , \Check1_CheckInst_3_n82 ,
         \Check1_CheckInst_3_n81 , \Check1_CheckInst_3_n80 ,
         \Check1_CheckInst_3_n79 , \Check1_CheckInst_3_n78 ,
         \Check1_CheckInst_3_n77 , \Check1_CheckInst_3_n76 ,
         \Check1_CheckInst_3_n75 , \Check1_CheckInst_3_n74 ,
         \Check1_CheckInst_3_n73 , \Check1_CheckInst_3_n72 ,
         \Check1_CheckInst_3_n71 , \Check1_CheckInst_3_n70 ,
         \Check1_CheckInst_3_n69 , \Check1_CheckInst_3_n68 ,
         \Check1_CheckInst_3_n67 , \Check1_CheckInst_3_n66 ,
         \Check1_CheckInst_3_n65 , \Check1_CheckInst_3_n64 ,
         \Check1_CheckInst_3_n63 , \Check1_CheckInst_3_n62 ,
         \Check1_CheckInst_3_n61 , \Check1_CheckInst_3_n60 ,
         \Check1_CheckInst_3_n59 , \Check1_CheckInst_3_n58 ,
         \Check1_CheckInst_3_n57 , \Check1_CheckInst_3_n56 ,
         \Check1_CheckInst_3_n55 , \Check1_CheckInst_3_n54 ,
         \Check1_CheckInst_3_n53 , \Check1_CheckInst_3_n52 ,
         \Check1_CheckInst_3_n51 , \Check1_CheckInst_3_n50 ,
         \Check1_CheckInst_3_n49 , \Check1_CheckInst_3_n48 ,
         \Check1_CheckInst_3_n47 , \Check1_CheckInst_3_n46 ,
         \Check1_CheckInst_3_n45 , \Check1_CheckInst_3_n44 ,
         \Check1_CheckInst_3_n43 , \Check1_CheckInst_3_n42 ,
         \Check1_CheckInst_3_n41 , \Check1_CheckInst_3_n40 ,
         \Check1_CheckInst_3_n39 , \Check1_CheckInst_3_n38 ,
         \Check1_CheckInst_3_n37 , \Check1_CheckInst_3_n36 ,
         \Check1_CheckInst_3_n35 , \Check1_CheckInst_3_n34 ,
         \Check1_CheckInst_3_n33 , \Check1_CheckInst_3_n32 ,
         \Check1_CheckInst_3_n31 , \Check1_CheckInst_3_n30 ,
         \Check1_CheckInst_3_n29 , \Check1_CheckInst_3_n28 ,
         \Check1_CheckInst_3_n27 , \Check1_CheckInst_3_n26 ,
         \Check1_CheckInst_3_n25 , \Check1_CheckInst_3_n24 ,
         \Check1_CheckInst_3_n23 , \Check1_CheckInst_3_n22 ,
         \Check1_CheckInst_3_n21 , \Check1_CheckInst_3_n20 ,
         \Check1_CheckInst_3_n19 , \Check1_CheckInst_3_n18 ,
         \Check1_CheckInst_3_n17 , \Check1_CheckInst_3_n16 ,
         \Check1_CheckInst_3_n15 , \Check1_CheckInst_3_n14 ,
         \Check1_CheckInst_3_n13 , \Check1_CheckInst_3_n12 ,
         \Check1_CheckInst_3_n11 , \Check1_CheckInst_3_n10 ,
         \Check1_CheckInst_3_n9 , \Check1_CheckInst_3_n8 ,
         \Check1_CheckInst_3_n7 , \Check1_CheckInst_3_n6 ,
         \Check1_CheckInst_3_n5 , \Check1_CheckInst_3_n4 ,
         \Check1_CheckInst_3_n3 ;
  wire   [63:0] MCOutput;
  wire   [63:0] AddRoundKeyOutput;
  wire   [63:0] PermutationOutput;
  wire   [63:0] Feedback;
  wire   [63:0] MCOutput2;
  wire   [63:0] AddRoundKeyOutput2;
  wire   [63:0] PermutationOutput2;
  wire   [63:0] Feedback2;
  wire   [63:0] MCOutput3;
  wire   [63:0] AddRoundKeyOutput3;
  wire   [63:0] PermutationOutput3;
  wire   [63:0] Red_Input;
  wire   [63:0] Red_MCOutput;
  wire   [63:0] Red_K0;
  wire   [63:0] Red_AddRoundKeyOutput;
  wire   [63:0] Red_StateRegOutput;
  wire   [63:0] Red_Feedback;
  wire   [63:0] Red_MCOutput2;
  wire   [63:0] Red_K1;
  wire   [63:0] Red_AddRoundKeyOutput2;
  wire   [63:0] Red_StateRegOutput2;
  wire   [63:0] Red_Feedback2;
  wire   [63:0] Red_MCOutput3;
  wire   [63:0] Red_K2;
  wire   [63:0] Red_AddRoundKeyOutput3;
  wire   [63:0] Red_StateRegOutput3;
  wire   [63:0] Red_Feedback3;
  wire   [447:0] Red_SignaltoCheck;
  wire   [3:0] Error;

  NAND2_X1 U9 ( .A1(Error[2]), .A2(Error[3]), .ZN(n9) );
  NAND2_X1 U10 ( .A1(Error[0]), .A2(Error[1]), .ZN(n8) );
  OR2_X1 U11 ( .A1(n9), .A2(n8), .ZN(ErrorFlag) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_0_U2  ( .A(\MCInst_XOR_r0_Inst_0_n3 ), .B(
        Input[0]), .ZN(MCOutput[48]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_0_U1  ( .A(Input[48]), .B(Input[16]), .ZN(
        \MCInst_XOR_r0_Inst_0_n3 ) );
  XOR2_X1 \MCInst_XOR_r1_Inst_0_U1  ( .A(Input[32]), .B(Input[0]), .Z(
        MCOutput[32]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_1_U2  ( .A(\MCInst_XOR_r0_Inst_1_n3 ), .B(
        Input[1]), .ZN(MCOutput[49]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_1_U1  ( .A(Input[49]), .B(Input[17]), .ZN(
        \MCInst_XOR_r0_Inst_1_n3 ) );
  XOR2_X1 \MCInst_XOR_r1_Inst_1_U1  ( .A(Input[33]), .B(Input[1]), .Z(
        MCOutput[33]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_2_U2  ( .A(\MCInst_XOR_r0_Inst_2_n3 ), .B(
        Input[2]), .ZN(MCOutput[50]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_2_U1  ( .A(Input[50]), .B(Input[18]), .ZN(
        \MCInst_XOR_r0_Inst_2_n3 ) );
  XOR2_X1 \MCInst_XOR_r1_Inst_2_U1  ( .A(Input[34]), .B(Input[2]), .Z(
        MCOutput[34]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_3_U2  ( .A(\MCInst_XOR_r0_Inst_3_n3 ), .B(
        Input[3]), .ZN(MCOutput[51]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_3_U1  ( .A(Input[51]), .B(Input[19]), .ZN(
        \MCInst_XOR_r0_Inst_3_n3 ) );
  XOR2_X1 \MCInst_XOR_r1_Inst_3_U1  ( .A(Input[35]), .B(Input[3]), .Z(
        MCOutput[35]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_4_U2  ( .A(\MCInst_XOR_r0_Inst_4_n3 ), .B(
        Input[4]), .ZN(MCOutput[52]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_4_U1  ( .A(Input[52]), .B(Input[20]), .ZN(
        \MCInst_XOR_r0_Inst_4_n3 ) );
  XOR2_X1 \MCInst_XOR_r1_Inst_4_U1  ( .A(Input[36]), .B(Input[4]), .Z(
        MCOutput[36]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_5_U2  ( .A(\MCInst_XOR_r0_Inst_5_n3 ), .B(
        Input[5]), .ZN(MCOutput[53]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_5_U1  ( .A(Input[53]), .B(Input[21]), .ZN(
        \MCInst_XOR_r0_Inst_5_n3 ) );
  XOR2_X1 \MCInst_XOR_r1_Inst_5_U1  ( .A(Input[37]), .B(Input[5]), .Z(
        MCOutput[37]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_6_U2  ( .A(\MCInst_XOR_r0_Inst_6_n3 ), .B(
        Input[6]), .ZN(MCOutput[54]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_6_U1  ( .A(Input[54]), .B(Input[22]), .ZN(
        \MCInst_XOR_r0_Inst_6_n3 ) );
  XOR2_X1 \MCInst_XOR_r1_Inst_6_U1  ( .A(Input[38]), .B(Input[6]), .Z(
        MCOutput[38]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_7_U2  ( .A(\MCInst_XOR_r0_Inst_7_n3 ), .B(
        Input[7]), .ZN(MCOutput[55]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_7_U1  ( .A(Input[55]), .B(Input[23]), .ZN(
        \MCInst_XOR_r0_Inst_7_n3 ) );
  XOR2_X1 \MCInst_XOR_r1_Inst_7_U1  ( .A(Input[39]), .B(Input[7]), .Z(
        MCOutput[39]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_8_U2  ( .A(\MCInst_XOR_r0_Inst_8_n3 ), .B(
        Input[8]), .ZN(MCOutput[56]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_8_U1  ( .A(Input[56]), .B(Input[24]), .ZN(
        \MCInst_XOR_r0_Inst_8_n3 ) );
  XOR2_X1 \MCInst_XOR_r1_Inst_8_U1  ( .A(Input[40]), .B(Input[8]), .Z(
        MCOutput[40]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_9_U2  ( .A(\MCInst_XOR_r0_Inst_9_n3 ), .B(
        Input[9]), .ZN(MCOutput[57]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_9_U1  ( .A(Input[57]), .B(Input[25]), .ZN(
        \MCInst_XOR_r0_Inst_9_n3 ) );
  XOR2_X1 \MCInst_XOR_r1_Inst_9_U1  ( .A(Input[41]), .B(Input[9]), .Z(
        MCOutput[41]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_10_U2  ( .A(\MCInst_XOR_r0_Inst_10_n3 ), .B(
        Input[10]), .ZN(MCOutput[58]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_10_U1  ( .A(Input[58]), .B(Input[26]), .ZN(
        \MCInst_XOR_r0_Inst_10_n3 ) );
  XOR2_X1 \MCInst_XOR_r1_Inst_10_U1  ( .A(Input[42]), .B(Input[10]), .Z(
        MCOutput[42]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_11_U2  ( .A(\MCInst_XOR_r0_Inst_11_n3 ), .B(
        Input[11]), .ZN(MCOutput[59]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_11_U1  ( .A(Input[59]), .B(Input[27]), .ZN(
        \MCInst_XOR_r0_Inst_11_n3 ) );
  XOR2_X1 \MCInst_XOR_r1_Inst_11_U1  ( .A(Input[43]), .B(Input[11]), .Z(
        MCOutput[43]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_12_U2  ( .A(\MCInst_XOR_r0_Inst_12_n3 ), .B(
        Input[12]), .ZN(MCOutput[60]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_12_U1  ( .A(Input[60]), .B(Input[28]), .ZN(
        \MCInst_XOR_r0_Inst_12_n3 ) );
  XOR2_X1 \MCInst_XOR_r1_Inst_12_U1  ( .A(Input[44]), .B(Input[12]), .Z(
        MCOutput[44]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_13_U2  ( .A(\MCInst_XOR_r0_Inst_13_n3 ), .B(
        Input[13]), .ZN(MCOutput[61]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_13_U1  ( .A(Input[61]), .B(Input[29]), .ZN(
        \MCInst_XOR_r0_Inst_13_n3 ) );
  XOR2_X1 \MCInst_XOR_r1_Inst_13_U1  ( .A(Input[45]), .B(Input[13]), .Z(
        MCOutput[45]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_14_U2  ( .A(\MCInst_XOR_r0_Inst_14_n3 ), .B(
        Input[14]), .ZN(MCOutput[62]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_14_U1  ( .A(Input[62]), .B(Input[30]), .ZN(
        \MCInst_XOR_r0_Inst_14_n3 ) );
  XOR2_X1 \MCInst_XOR_r1_Inst_14_U1  ( .A(Input[46]), .B(Input[14]), .Z(
        MCOutput[46]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_15_U2  ( .A(\MCInst_XOR_r0_Inst_15_n3 ), .B(
        Input[15]), .ZN(MCOutput[63]) );
  XNOR2_X1 \MCInst_XOR_r0_Inst_15_U1  ( .A(Input[63]), .B(Input[31]), .ZN(
        \MCInst_XOR_r0_Inst_15_n3 ) );
  XOR2_X1 \MCInst_XOR_r1_Inst_15_U1  ( .A(Input[47]), .B(Input[15]), .Z(
        MCOutput[47]) );
  XOR2_X1 \AddKeyXOR1_XORInst_0_0_U1  ( .A(MCOutput[48]), .B(Key[176]), .Z(
        AddRoundKeyOutput[48]) );
  XOR2_X1 \AddKeyXOR1_XORInst_0_1_U1  ( .A(MCOutput[49]), .B(Key[177]), .Z(
        AddRoundKeyOutput[49]) );
  XOR2_X1 \AddKeyXOR1_XORInst_0_2_U1  ( .A(MCOutput[50]), .B(Key[178]), .Z(
        AddRoundKeyOutput[50]) );
  XOR2_X1 \AddKeyXOR1_XORInst_0_3_U1  ( .A(MCOutput[51]), .B(Key[179]), .Z(
        AddRoundKeyOutput[51]) );
  XOR2_X1 \AddKeyXOR1_XORInst_1_0_U1  ( .A(MCOutput[52]), .B(Key[180]), .Z(
        AddRoundKeyOutput[52]) );
  XOR2_X1 \AddKeyXOR1_XORInst_1_1_U1  ( .A(MCOutput[53]), .B(Key[181]), .Z(
        AddRoundKeyOutput[53]) );
  XOR2_X1 \AddKeyXOR1_XORInst_1_2_U1  ( .A(MCOutput[54]), .B(Key[182]), .Z(
        AddRoundKeyOutput[54]) );
  XOR2_X1 \AddKeyXOR1_XORInst_1_3_U1  ( .A(MCOutput[55]), .B(Key[183]), .Z(
        AddRoundKeyOutput[55]) );
  XOR2_X1 \AddKeyXOR1_XORInst_2_0_U1  ( .A(MCOutput[56]), .B(Key[184]), .Z(
        AddRoundKeyOutput[56]) );
  XOR2_X1 \AddKeyXOR1_XORInst_2_1_U1  ( .A(MCOutput[57]), .B(Key[185]), .Z(
        AddRoundKeyOutput[57]) );
  XOR2_X1 \AddKeyXOR1_XORInst_2_2_U1  ( .A(MCOutput[58]), .B(Key[186]), .Z(
        AddRoundKeyOutput[58]) );
  XOR2_X1 \AddKeyXOR1_XORInst_2_3_U1  ( .A(MCOutput[59]), .B(Key[187]), .Z(
        AddRoundKeyOutput[59]) );
  XOR2_X1 \AddKeyXOR1_XORInst_3_0_U1  ( .A(MCOutput[60]), .B(Key[188]), .Z(
        AddRoundKeyOutput[60]) );
  XOR2_X1 \AddKeyXOR1_XORInst_3_1_U1  ( .A(MCOutput[61]), .B(Key[189]), .Z(
        AddRoundKeyOutput[61]) );
  XOR2_X1 \AddKeyXOR1_XORInst_3_2_U1  ( .A(MCOutput[62]), .B(Key[190]), .Z(
        AddRoundKeyOutput[62]) );
  XOR2_X1 \AddKeyXOR1_XORInst_3_3_U1  ( .A(MCOutput[63]), .B(Key[191]), .Z(
        AddRoundKeyOutput[63]) );
  XOR2_X1 \AddKeyConstXOR_XORInst_0_0_U1  ( .A(Key[168]), .B(MCOutput[40]), 
        .Z(AddRoundKeyOutput[40]) );
  XOR2_X1 \AddKeyConstXOR_XORInst_0_1_U1  ( .A(Key[169]), .B(MCOutput[41]), 
        .Z(AddRoundKeyOutput[41]) );
  XOR2_X1 \AddKeyConstXOR_XORInst_0_2_U1  ( .A(Key[170]), .B(MCOutput[42]), 
        .Z(AddRoundKeyOutput[42]) );
  XOR2_X1 \AddKeyConstXOR_XORInst_0_3_U1  ( .A(Key[171]), .B(MCOutput[43]), 
        .Z(AddRoundKeyOutput[43]) );
  XOR2_X1 \AddKeyConstXOR_XORInst_1_0_U1  ( .A(Key[172]), .B(MCOutput[44]), 
        .Z(AddRoundKeyOutput[44]) );
  XOR2_X1 \AddKeyConstXOR_XORInst_1_1_U1  ( .A(Key[173]), .B(MCOutput[45]), 
        .Z(AddRoundKeyOutput[45]) );
  XOR2_X1 \AddKeyConstXOR_XORInst_1_2_U1  ( .A(Key[174]), .B(MCOutput[46]), 
        .Z(AddRoundKeyOutput[46]) );
  XOR2_X1 \AddKeyConstXOR_XORInst_1_3_U1  ( .A(Key[175]), .B(MCOutput[47]), 
        .Z(AddRoundKeyOutput[47]) );
  XOR2_X1 \AddKeyXOR2_XORInst_0_0_U1  ( .A(Input[0]), .B(Key[128]), .Z(
        AddRoundKeyOutput[0]) );
  XOR2_X1 \AddKeyXOR2_XORInst_0_1_U1  ( .A(Input[1]), .B(Key[129]), .Z(
        AddRoundKeyOutput[1]) );
  XOR2_X1 \AddKeyXOR2_XORInst_0_2_U1  ( .A(Input[2]), .B(Key[130]), .Z(
        AddRoundKeyOutput[2]) );
  XOR2_X1 \AddKeyXOR2_XORInst_0_3_U1  ( .A(Input[3]), .B(Key[131]), .Z(
        AddRoundKeyOutput[3]) );
  XOR2_X1 \AddKeyXOR2_XORInst_1_0_U1  ( .A(Input[4]), .B(Key[132]), .Z(
        AddRoundKeyOutput[4]) );
  XOR2_X1 \AddKeyXOR2_XORInst_1_1_U1  ( .A(Input[5]), .B(Key[133]), .Z(
        AddRoundKeyOutput[5]) );
  XOR2_X1 \AddKeyXOR2_XORInst_1_2_U1  ( .A(Input[6]), .B(Key[134]), .Z(
        AddRoundKeyOutput[6]) );
  XOR2_X1 \AddKeyXOR2_XORInst_1_3_U1  ( .A(Input[7]), .B(Key[135]), .Z(
        AddRoundKeyOutput[7]) );
  XOR2_X1 \AddKeyXOR2_XORInst_2_0_U1  ( .A(Input[8]), .B(Key[136]), .Z(
        AddRoundKeyOutput[8]) );
  XOR2_X1 \AddKeyXOR2_XORInst_2_1_U1  ( .A(Input[9]), .B(Key[137]), .Z(
        AddRoundKeyOutput[9]) );
  XOR2_X1 \AddKeyXOR2_XORInst_2_2_U1  ( .A(Input[10]), .B(Key[138]), .Z(
        AddRoundKeyOutput[10]) );
  XOR2_X1 \AddKeyXOR2_XORInst_2_3_U1  ( .A(Input[11]), .B(Key[139]), .Z(
        AddRoundKeyOutput[11]) );
  XOR2_X1 \AddKeyXOR2_XORInst_3_0_U1  ( .A(Input[12]), .B(Key[140]), .Z(
        AddRoundKeyOutput[12]) );
  XOR2_X1 \AddKeyXOR2_XORInst_3_1_U1  ( .A(Input[13]), .B(Key[141]), .Z(
        AddRoundKeyOutput[13]) );
  XOR2_X1 \AddKeyXOR2_XORInst_3_2_U1  ( .A(Input[14]), .B(Key[142]), .Z(
        AddRoundKeyOutput[14]) );
  XOR2_X1 \AddKeyXOR2_XORInst_3_3_U1  ( .A(Input[15]), .B(Key[143]), .Z(
        AddRoundKeyOutput[15]) );
  XOR2_X1 \AddKeyXOR2_XORInst_4_0_U1  ( .A(Input[16]), .B(Key[144]), .Z(
        AddRoundKeyOutput[16]) );
  XOR2_X1 \AddKeyXOR2_XORInst_4_1_U1  ( .A(Input[17]), .B(Key[145]), .Z(
        AddRoundKeyOutput[17]) );
  XOR2_X1 \AddKeyXOR2_XORInst_4_2_U1  ( .A(Input[18]), .B(Key[146]), .Z(
        AddRoundKeyOutput[18]) );
  XOR2_X1 \AddKeyXOR2_XORInst_4_3_U1  ( .A(Input[19]), .B(Key[147]), .Z(
        AddRoundKeyOutput[19]) );
  XOR2_X1 \AddKeyXOR2_XORInst_5_0_U1  ( .A(Input[20]), .B(Key[148]), .Z(
        AddRoundKeyOutput[20]) );
  XOR2_X1 \AddKeyXOR2_XORInst_5_1_U1  ( .A(Input[21]), .B(Key[149]), .Z(
        AddRoundKeyOutput[21]) );
  XOR2_X1 \AddKeyXOR2_XORInst_5_2_U1  ( .A(Input[22]), .B(Key[150]), .Z(
        AddRoundKeyOutput[22]) );
  XOR2_X1 \AddKeyXOR2_XORInst_5_3_U1  ( .A(Input[23]), .B(Key[151]), .Z(
        AddRoundKeyOutput[23]) );
  XOR2_X1 \AddKeyXOR2_XORInst_6_0_U1  ( .A(Input[24]), .B(Key[152]), .Z(
        AddRoundKeyOutput[24]) );
  XOR2_X1 \AddKeyXOR2_XORInst_6_1_U1  ( .A(Input[25]), .B(Key[153]), .Z(
        AddRoundKeyOutput[25]) );
  XOR2_X1 \AddKeyXOR2_XORInst_6_2_U1  ( .A(Input[26]), .B(Key[154]), .Z(
        AddRoundKeyOutput[26]) );
  XOR2_X1 \AddKeyXOR2_XORInst_6_3_U1  ( .A(Input[27]), .B(Key[155]), .Z(
        AddRoundKeyOutput[27]) );
  XOR2_X1 \AddKeyXOR2_XORInst_7_0_U1  ( .A(Input[28]), .B(Key[156]), .Z(
        AddRoundKeyOutput[28]) );
  XOR2_X1 \AddKeyXOR2_XORInst_7_1_U1  ( .A(Input[29]), .B(Key[157]), .Z(
        AddRoundKeyOutput[29]) );
  XOR2_X1 \AddKeyXOR2_XORInst_7_2_U1  ( .A(Input[30]), .B(Key[158]), .Z(
        AddRoundKeyOutput[30]) );
  XOR2_X1 \AddKeyXOR2_XORInst_7_3_U1  ( .A(Input[31]), .B(Key[159]), .Z(
        AddRoundKeyOutput[31]) );
  XOR2_X1 \AddKeyXOR2_XORInst_8_0_U1  ( .A(MCOutput[32]), .B(Key[160]), .Z(
        AddRoundKeyOutput[32]) );
  XOR2_X1 \AddKeyXOR2_XORInst_8_1_U1  ( .A(MCOutput[33]), .B(Key[161]), .Z(
        AddRoundKeyOutput[33]) );
  XOR2_X1 \AddKeyXOR2_XORInst_8_2_U1  ( .A(MCOutput[34]), .B(Key[162]), .Z(
        AddRoundKeyOutput[34]) );
  XOR2_X1 \AddKeyXOR2_XORInst_8_3_U1  ( .A(MCOutput[35]), .B(Key[163]), .Z(
        AddRoundKeyOutput[35]) );
  XOR2_X1 \AddKeyXOR2_XORInst_9_0_U1  ( .A(MCOutput[36]), .B(Key[164]), .Z(
        AddRoundKeyOutput[36]) );
  XOR2_X1 \AddKeyXOR2_XORInst_9_1_U1  ( .A(MCOutput[37]), .B(Key[165]), .Z(
        AddRoundKeyOutput[37]) );
  XOR2_X1 \AddKeyXOR2_XORInst_9_2_U1  ( .A(MCOutput[38]), .B(Key[166]), .Z(
        AddRoundKeyOutput[38]) );
  XOR2_X1 \AddKeyXOR2_XORInst_9_3_U1  ( .A(MCOutput[39]), .B(Key[167]), .Z(
        AddRoundKeyOutput[39]) );
  DFF_X1 \StateReg_s_current_state_reg[0]  ( .D(AddRoundKeyOutput[0]), .CK(clk), .Q(PermutationOutput[60]) );
  DFF_X1 \StateReg_s_current_state_reg[1]  ( .D(AddRoundKeyOutput[1]), .CK(clk), .Q(PermutationOutput[61]) );
  DFF_X1 \StateReg_s_current_state_reg[2]  ( .D(AddRoundKeyOutput[2]), .CK(clk), .Q(PermutationOutput[62]) );
  DFF_X1 \StateReg_s_current_state_reg[3]  ( .D(AddRoundKeyOutput[3]), .CK(clk), .Q(PermutationOutput[63]) );
  DFF_X1 \StateReg_s_current_state_reg[4]  ( .D(AddRoundKeyOutput[4]), .CK(clk), .Q(PermutationOutput[48]) );
  DFF_X1 \StateReg_s_current_state_reg[5]  ( .D(AddRoundKeyOutput[5]), .CK(clk), .Q(PermutationOutput[49]) );
  DFF_X1 \StateReg_s_current_state_reg[6]  ( .D(AddRoundKeyOutput[6]), .CK(clk), .Q(PermutationOutput[50]) );
  DFF_X1 \StateReg_s_current_state_reg[7]  ( .D(AddRoundKeyOutput[7]), .CK(clk), .Q(PermutationOutput[51]) );
  DFF_X1 \StateReg_s_current_state_reg[8]  ( .D(AddRoundKeyOutput[8]), .CK(clk), .Q(PermutationOutput[52]) );
  DFF_X1 \StateReg_s_current_state_reg[9]  ( .D(AddRoundKeyOutput[9]), .CK(clk), .Q(PermutationOutput[53]) );
  DFF_X1 \StateReg_s_current_state_reg[10]  ( .D(AddRoundKeyOutput[10]), .CK(
        clk), .Q(PermutationOutput[54]) );
  DFF_X1 \StateReg_s_current_state_reg[11]  ( .D(AddRoundKeyOutput[11]), .CK(
        clk), .Q(PermutationOutput[55]) );
  DFF_X1 \StateReg_s_current_state_reg[12]  ( .D(AddRoundKeyOutput[12]), .CK(
        clk), .Q(PermutationOutput[56]) );
  DFF_X1 \StateReg_s_current_state_reg[13]  ( .D(AddRoundKeyOutput[13]), .CK(
        clk), .Q(PermutationOutput[57]) );
  DFF_X1 \StateReg_s_current_state_reg[14]  ( .D(AddRoundKeyOutput[14]), .CK(
        clk), .Q(PermutationOutput[58]) );
  DFF_X1 \StateReg_s_current_state_reg[15]  ( .D(AddRoundKeyOutput[15]), .CK(
        clk), .Q(PermutationOutput[59]) );
  DFF_X1 \StateReg_s_current_state_reg[16]  ( .D(AddRoundKeyOutput[16]), .CK(
        clk), .Q(PermutationOutput[32]) );
  DFF_X1 \StateReg_s_current_state_reg[17]  ( .D(AddRoundKeyOutput[17]), .CK(
        clk), .Q(PermutationOutput[33]) );
  DFF_X1 \StateReg_s_current_state_reg[18]  ( .D(AddRoundKeyOutput[18]), .CK(
        clk), .Q(PermutationOutput[34]) );
  DFF_X1 \StateReg_s_current_state_reg[19]  ( .D(AddRoundKeyOutput[19]), .CK(
        clk), .Q(PermutationOutput[35]) );
  DFF_X1 \StateReg_s_current_state_reg[20]  ( .D(AddRoundKeyOutput[20]), .CK(
        clk), .Q(PermutationOutput[44]) );
  DFF_X1 \StateReg_s_current_state_reg[21]  ( .D(AddRoundKeyOutput[21]), .CK(
        clk), .Q(PermutationOutput[45]) );
  DFF_X1 \StateReg_s_current_state_reg[22]  ( .D(AddRoundKeyOutput[22]), .CK(
        clk), .Q(PermutationOutput[46]) );
  DFF_X1 \StateReg_s_current_state_reg[23]  ( .D(AddRoundKeyOutput[23]), .CK(
        clk), .Q(PermutationOutput[47]) );
  DFF_X1 \StateReg_s_current_state_reg[24]  ( .D(AddRoundKeyOutput[24]), .CK(
        clk), .Q(PermutationOutput[40]) );
  DFF_X1 \StateReg_s_current_state_reg[25]  ( .D(AddRoundKeyOutput[25]), .CK(
        clk), .Q(PermutationOutput[41]) );
  DFF_X1 \StateReg_s_current_state_reg[26]  ( .D(AddRoundKeyOutput[26]), .CK(
        clk), .Q(PermutationOutput[42]) );
  DFF_X1 \StateReg_s_current_state_reg[27]  ( .D(AddRoundKeyOutput[27]), .CK(
        clk), .Q(PermutationOutput[43]) );
  DFF_X1 \StateReg_s_current_state_reg[28]  ( .D(AddRoundKeyOutput[28]), .CK(
        clk), .Q(PermutationOutput[36]) );
  DFF_X1 \StateReg_s_current_state_reg[29]  ( .D(AddRoundKeyOutput[29]), .CK(
        clk), .Q(PermutationOutput[37]) );
  DFF_X1 \StateReg_s_current_state_reg[30]  ( .D(AddRoundKeyOutput[30]), .CK(
        clk), .Q(PermutationOutput[38]) );
  DFF_X1 \StateReg_s_current_state_reg[31]  ( .D(AddRoundKeyOutput[31]), .CK(
        clk), .Q(PermutationOutput[39]) );
  DFF_X1 \StateReg_s_current_state_reg[32]  ( .D(AddRoundKeyOutput[32]), .CK(
        clk), .Q(PermutationOutput[16]) );
  DFF_X1 \StateReg_s_current_state_reg[33]  ( .D(AddRoundKeyOutput[33]), .CK(
        clk), .Q(PermutationOutput[17]) );
  DFF_X1 \StateReg_s_current_state_reg[34]  ( .D(AddRoundKeyOutput[34]), .CK(
        clk), .Q(PermutationOutput[18]) );
  DFF_X1 \StateReg_s_current_state_reg[35]  ( .D(AddRoundKeyOutput[35]), .CK(
        clk), .Q(PermutationOutput[19]) );
  DFF_X1 \StateReg_s_current_state_reg[36]  ( .D(AddRoundKeyOutput[36]), .CK(
        clk), .Q(PermutationOutput[28]) );
  DFF_X1 \StateReg_s_current_state_reg[37]  ( .D(AddRoundKeyOutput[37]), .CK(
        clk), .Q(PermutationOutput[29]) );
  DFF_X1 \StateReg_s_current_state_reg[38]  ( .D(AddRoundKeyOutput[38]), .CK(
        clk), .Q(PermutationOutput[30]) );
  DFF_X1 \StateReg_s_current_state_reg[39]  ( .D(AddRoundKeyOutput[39]), .CK(
        clk), .Q(PermutationOutput[31]) );
  DFF_X1 \StateReg_s_current_state_reg[40]  ( .D(AddRoundKeyOutput[40]), .CK(
        clk), .Q(PermutationOutput[24]) );
  DFF_X1 \StateReg_s_current_state_reg[41]  ( .D(AddRoundKeyOutput[41]), .CK(
        clk), .Q(PermutationOutput[25]) );
  DFF_X1 \StateReg_s_current_state_reg[42]  ( .D(AddRoundKeyOutput[42]), .CK(
        clk), .Q(PermutationOutput[26]) );
  DFF_X1 \StateReg_s_current_state_reg[43]  ( .D(AddRoundKeyOutput[43]), .CK(
        clk), .Q(PermutationOutput[27]) );
  DFF_X1 \StateReg_s_current_state_reg[44]  ( .D(AddRoundKeyOutput[44]), .CK(
        clk), .Q(PermutationOutput[20]) );
  DFF_X1 \StateReg_s_current_state_reg[45]  ( .D(AddRoundKeyOutput[45]), .CK(
        clk), .Q(PermutationOutput[21]) );
  DFF_X1 \StateReg_s_current_state_reg[46]  ( .D(AddRoundKeyOutput[46]), .CK(
        clk), .Q(PermutationOutput[22]) );
  DFF_X1 \StateReg_s_current_state_reg[47]  ( .D(AddRoundKeyOutput[47]), .CK(
        clk), .Q(PermutationOutput[23]) );
  DFF_X1 \StateReg_s_current_state_reg[48]  ( .D(AddRoundKeyOutput[48]), .CK(
        clk), .Q(PermutationOutput[4]) );
  DFF_X1 \StateReg_s_current_state_reg[49]  ( .D(AddRoundKeyOutput[49]), .CK(
        clk), .Q(PermutationOutput[5]) );
  DFF_X1 \StateReg_s_current_state_reg[50]  ( .D(AddRoundKeyOutput[50]), .CK(
        clk), .Q(PermutationOutput[6]) );
  DFF_X1 \StateReg_s_current_state_reg[51]  ( .D(AddRoundKeyOutput[51]), .CK(
        clk), .Q(PermutationOutput[7]) );
  DFF_X1 \StateReg_s_current_state_reg[52]  ( .D(AddRoundKeyOutput[52]), .CK(
        clk), .Q(PermutationOutput[8]) );
  DFF_X1 \StateReg_s_current_state_reg[53]  ( .D(AddRoundKeyOutput[53]), .CK(
        clk), .Q(PermutationOutput[9]) );
  DFF_X1 \StateReg_s_current_state_reg[54]  ( .D(AddRoundKeyOutput[54]), .CK(
        clk), .Q(PermutationOutput[10]) );
  DFF_X1 \StateReg_s_current_state_reg[55]  ( .D(AddRoundKeyOutput[55]), .CK(
        clk), .Q(PermutationOutput[11]) );
  DFF_X1 \StateReg_s_current_state_reg[56]  ( .D(AddRoundKeyOutput[56]), .CK(
        clk), .Q(PermutationOutput[12]) );
  DFF_X1 \StateReg_s_current_state_reg[57]  ( .D(AddRoundKeyOutput[57]), .CK(
        clk), .Q(PermutationOutput[13]) );
  DFF_X1 \StateReg_s_current_state_reg[58]  ( .D(AddRoundKeyOutput[58]), .CK(
        clk), .Q(PermutationOutput[14]) );
  DFF_X1 \StateReg_s_current_state_reg[59]  ( .D(AddRoundKeyOutput[59]), .CK(
        clk), .Q(PermutationOutput[15]) );
  DFF_X1 \StateReg_s_current_state_reg[60]  ( .D(AddRoundKeyOutput[60]), .CK(
        clk), .Q(PermutationOutput[0]) );
  DFF_X1 \StateReg_s_current_state_reg[61]  ( .D(AddRoundKeyOutput[61]), .CK(
        clk), .Q(PermutationOutput[1]) );
  DFF_X1 \StateReg_s_current_state_reg[62]  ( .D(AddRoundKeyOutput[62]), .CK(
        clk), .Q(PermutationOutput[2]) );
  DFF_X1 \StateReg_s_current_state_reg[63]  ( .D(AddRoundKeyOutput[63]), .CK(
        clk), .Q(PermutationOutput[3]) );
  NOR2_X1 \SubCellInst_LFInst_0_LFInst_0_U8  ( .A1(
        \SubCellInst_LFInst_0_LFInst_0_n11 ), .A2(
        \SubCellInst_LFInst_0_LFInst_0_n10 ), .ZN(MCOutput2[0]) );
  AND2_X1 \SubCellInst_LFInst_0_LFInst_0_U7  ( .A1(PermutationOutput[3]), .A2(
        PermutationOutput[2]), .ZN(\SubCellInst_LFInst_0_LFInst_0_n10 ) );
  NOR2_X1 \SubCellInst_LFInst_0_LFInst_0_U6  ( .A1(PermutationOutput[1]), .A2(
        \SubCellInst_LFInst_0_LFInst_0_n9 ), .ZN(
        \SubCellInst_LFInst_0_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst_LFInst_0_LFInst_0_U5  ( .A1(
        \SubCellInst_LFInst_0_LFInst_0_n8 ), .A2(
        \SubCellInst_LFInst_0_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_0_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst_LFInst_0_LFInst_0_U4  ( .A1(PermutationOutput[3]), .A2(
        PermutationOutput[2]), .ZN(\SubCellInst_LFInst_0_LFInst_0_n7 ) );
  INV_X1 \SubCellInst_LFInst_0_LFInst_0_U3  ( .A(PermutationOutput[0]), .ZN(
        \SubCellInst_LFInst_0_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst_LFInst_0_LFInst_1_U6  ( .A1(
        \SubCellInst_LFInst_0_LFInst_1_n6 ), .A2(
        \SubCellInst_LFInst_0_LFInst_1_n5 ), .ZN(MCOutput2[1]) );
  NAND2_X1 \SubCellInst_LFInst_0_LFInst_1_U5  ( .A1(PermutationOutput[2]), 
        .A2(PermutationOutput[0]), .ZN(\SubCellInst_LFInst_0_LFInst_1_n5 ) );
  OR2_X1 \SubCellInst_LFInst_0_LFInst_1_U4  ( .A1(PermutationOutput[3]), .A2(
        \SubCellInst_LFInst_0_LFInst_1_n4 ), .ZN(
        \SubCellInst_LFInst_0_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst_LFInst_0_LFInst_1_U3  ( .A1(PermutationOutput[2]), .A2(
        PermutationOutput[0]), .ZN(\SubCellInst_LFInst_0_LFInst_1_n4 ) );
  NAND2_X1 \SubCellInst_LFInst_0_LFInst_2_U8  ( .A1(
        \SubCellInst_LFInst_0_LFInst_2_n11 ), .A2(
        \SubCellInst_LFInst_0_LFInst_2_n10 ), .ZN(MCOutput2[2]) );
  OR2_X1 \SubCellInst_LFInst_0_LFInst_2_U7  ( .A1(PermutationOutput[0]), .A2(
        PermutationOutput[3]), .ZN(\SubCellInst_LFInst_0_LFInst_2_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_0_LFInst_2_U6  ( .A1(PermutationOutput[1]), 
        .A2(\SubCellInst_LFInst_0_LFInst_2_n9 ), .ZN(
        \SubCellInst_LFInst_0_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_0_LFInst_2_U5  ( .A1(
        \SubCellInst_LFInst_0_LFInst_2_n8 ), .A2(
        \SubCellInst_LFInst_0_LFInst_2_n7 ), .ZN(
        \SubCellInst_LFInst_0_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst_LFInst_0_LFInst_2_U4  ( .A1(PermutationOutput[0]), 
        .A2(PermutationOutput[3]), .ZN(\SubCellInst_LFInst_0_LFInst_2_n7 ) );
  INV_X1 \SubCellInst_LFInst_0_LFInst_2_U3  ( .A(PermutationOutput[2]), .ZN(
        \SubCellInst_LFInst_0_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst_LFInst_0_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_0_LFInst_3_n6 ), .A2(
        \SubCellInst_LFInst_0_LFInst_3_n5 ), .ZN(MCOutput2[3]) );
  NOR2_X1 \SubCellInst_LFInst_0_LFInst_3_U5  ( .A1(PermutationOutput[3]), .A2(
        PermutationOutput[0]), .ZN(\SubCellInst_LFInst_0_LFInst_3_n5 ) );
  NOR2_X1 \SubCellInst_LFInst_0_LFInst_3_U4  ( .A1(PermutationOutput[1]), .A2(
        \SubCellInst_LFInst_0_LFInst_3_n4 ), .ZN(
        \SubCellInst_LFInst_0_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst_LFInst_0_LFInst_3_U3  ( .A1(PermutationOutput[3]), .A2(
        PermutationOutput[2]), .ZN(\SubCellInst_LFInst_0_LFInst_3_n4 ) );
  NOR2_X1 \SubCellInst_LFInst_1_LFInst_0_U8  ( .A1(
        \SubCellInst_LFInst_1_LFInst_0_n11 ), .A2(
        \SubCellInst_LFInst_1_LFInst_0_n10 ), .ZN(MCOutput2[4]) );
  AND2_X1 \SubCellInst_LFInst_1_LFInst_0_U7  ( .A1(PermutationOutput[7]), .A2(
        PermutationOutput[6]), .ZN(\SubCellInst_LFInst_1_LFInst_0_n10 ) );
  NOR2_X1 \SubCellInst_LFInst_1_LFInst_0_U6  ( .A1(PermutationOutput[5]), .A2(
        \SubCellInst_LFInst_1_LFInst_0_n9 ), .ZN(
        \SubCellInst_LFInst_1_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst_LFInst_1_LFInst_0_U5  ( .A1(
        \SubCellInst_LFInst_1_LFInst_0_n8 ), .A2(
        \SubCellInst_LFInst_1_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_1_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst_LFInst_1_LFInst_0_U4  ( .A1(PermutationOutput[7]), .A2(
        PermutationOutput[6]), .ZN(\SubCellInst_LFInst_1_LFInst_0_n7 ) );
  INV_X1 \SubCellInst_LFInst_1_LFInst_0_U3  ( .A(PermutationOutput[4]), .ZN(
        \SubCellInst_LFInst_1_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst_LFInst_1_LFInst_1_U6  ( .A1(
        \SubCellInst_LFInst_1_LFInst_1_n6 ), .A2(
        \SubCellInst_LFInst_1_LFInst_1_n5 ), .ZN(MCOutput2[5]) );
  NAND2_X1 \SubCellInst_LFInst_1_LFInst_1_U5  ( .A1(PermutationOutput[6]), 
        .A2(PermutationOutput[4]), .ZN(\SubCellInst_LFInst_1_LFInst_1_n5 ) );
  OR2_X1 \SubCellInst_LFInst_1_LFInst_1_U4  ( .A1(PermutationOutput[7]), .A2(
        \SubCellInst_LFInst_1_LFInst_1_n4 ), .ZN(
        \SubCellInst_LFInst_1_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst_LFInst_1_LFInst_1_U3  ( .A1(PermutationOutput[6]), .A2(
        PermutationOutput[4]), .ZN(\SubCellInst_LFInst_1_LFInst_1_n4 ) );
  NAND2_X1 \SubCellInst_LFInst_1_LFInst_2_U8  ( .A1(
        \SubCellInst_LFInst_1_LFInst_2_n11 ), .A2(
        \SubCellInst_LFInst_1_LFInst_2_n10 ), .ZN(MCOutput2[6]) );
  OR2_X1 \SubCellInst_LFInst_1_LFInst_2_U7  ( .A1(PermutationOutput[4]), .A2(
        PermutationOutput[7]), .ZN(\SubCellInst_LFInst_1_LFInst_2_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_1_LFInst_2_U6  ( .A1(PermutationOutput[5]), 
        .A2(\SubCellInst_LFInst_1_LFInst_2_n9 ), .ZN(
        \SubCellInst_LFInst_1_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_1_LFInst_2_U5  ( .A1(
        \SubCellInst_LFInst_1_LFInst_2_n8 ), .A2(
        \SubCellInst_LFInst_1_LFInst_2_n7 ), .ZN(
        \SubCellInst_LFInst_1_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst_LFInst_1_LFInst_2_U4  ( .A1(PermutationOutput[4]), 
        .A2(PermutationOutput[7]), .ZN(\SubCellInst_LFInst_1_LFInst_2_n7 ) );
  INV_X1 \SubCellInst_LFInst_1_LFInst_2_U3  ( .A(PermutationOutput[6]), .ZN(
        \SubCellInst_LFInst_1_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst_LFInst_1_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_1_LFInst_3_n6 ), .A2(
        \SubCellInst_LFInst_1_LFInst_3_n5 ), .ZN(MCOutput2[7]) );
  NOR2_X1 \SubCellInst_LFInst_1_LFInst_3_U5  ( .A1(PermutationOutput[7]), .A2(
        PermutationOutput[4]), .ZN(\SubCellInst_LFInst_1_LFInst_3_n5 ) );
  NOR2_X1 \SubCellInst_LFInst_1_LFInst_3_U4  ( .A1(PermutationOutput[5]), .A2(
        \SubCellInst_LFInst_1_LFInst_3_n4 ), .ZN(
        \SubCellInst_LFInst_1_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst_LFInst_1_LFInst_3_U3  ( .A1(PermutationOutput[7]), .A2(
        PermutationOutput[6]), .ZN(\SubCellInst_LFInst_1_LFInst_3_n4 ) );
  NOR2_X1 \SubCellInst_LFInst_2_LFInst_0_U8  ( .A1(
        \SubCellInst_LFInst_2_LFInst_0_n11 ), .A2(
        \SubCellInst_LFInst_2_LFInst_0_n10 ), .ZN(MCOutput2[8]) );
  AND2_X1 \SubCellInst_LFInst_2_LFInst_0_U7  ( .A1(PermutationOutput[11]), 
        .A2(PermutationOutput[10]), .ZN(\SubCellInst_LFInst_2_LFInst_0_n10 )
         );
  NOR2_X1 \SubCellInst_LFInst_2_LFInst_0_U6  ( .A1(PermutationOutput[9]), .A2(
        \SubCellInst_LFInst_2_LFInst_0_n9 ), .ZN(
        \SubCellInst_LFInst_2_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst_LFInst_2_LFInst_0_U5  ( .A1(
        \SubCellInst_LFInst_2_LFInst_0_n8 ), .A2(
        \SubCellInst_LFInst_2_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_2_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst_LFInst_2_LFInst_0_U4  ( .A1(PermutationOutput[11]), 
        .A2(PermutationOutput[10]), .ZN(\SubCellInst_LFInst_2_LFInst_0_n7 ) );
  INV_X1 \SubCellInst_LFInst_2_LFInst_0_U3  ( .A(PermutationOutput[8]), .ZN(
        \SubCellInst_LFInst_2_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst_LFInst_2_LFInst_1_U6  ( .A1(
        \SubCellInst_LFInst_2_LFInst_1_n6 ), .A2(
        \SubCellInst_LFInst_2_LFInst_1_n5 ), .ZN(MCOutput2[9]) );
  NAND2_X1 \SubCellInst_LFInst_2_LFInst_1_U5  ( .A1(PermutationOutput[10]), 
        .A2(PermutationOutput[8]), .ZN(\SubCellInst_LFInst_2_LFInst_1_n5 ) );
  OR2_X1 \SubCellInst_LFInst_2_LFInst_1_U4  ( .A1(PermutationOutput[11]), .A2(
        \SubCellInst_LFInst_2_LFInst_1_n4 ), .ZN(
        \SubCellInst_LFInst_2_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst_LFInst_2_LFInst_1_U3  ( .A1(PermutationOutput[10]), 
        .A2(PermutationOutput[8]), .ZN(\SubCellInst_LFInst_2_LFInst_1_n4 ) );
  NAND2_X1 \SubCellInst_LFInst_2_LFInst_2_U8  ( .A1(
        \SubCellInst_LFInst_2_LFInst_2_n11 ), .A2(
        \SubCellInst_LFInst_2_LFInst_2_n10 ), .ZN(MCOutput2[10]) );
  OR2_X1 \SubCellInst_LFInst_2_LFInst_2_U7  ( .A1(PermutationOutput[8]), .A2(
        PermutationOutput[11]), .ZN(\SubCellInst_LFInst_2_LFInst_2_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_2_LFInst_2_U6  ( .A1(PermutationOutput[9]), 
        .A2(\SubCellInst_LFInst_2_LFInst_2_n9 ), .ZN(
        \SubCellInst_LFInst_2_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_2_LFInst_2_U5  ( .A1(
        \SubCellInst_LFInst_2_LFInst_2_n8 ), .A2(
        \SubCellInst_LFInst_2_LFInst_2_n7 ), .ZN(
        \SubCellInst_LFInst_2_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst_LFInst_2_LFInst_2_U4  ( .A1(PermutationOutput[8]), 
        .A2(PermutationOutput[11]), .ZN(\SubCellInst_LFInst_2_LFInst_2_n7 ) );
  INV_X1 \SubCellInst_LFInst_2_LFInst_2_U3  ( .A(PermutationOutput[10]), .ZN(
        \SubCellInst_LFInst_2_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst_LFInst_2_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_2_LFInst_3_n6 ), .A2(
        \SubCellInst_LFInst_2_LFInst_3_n5 ), .ZN(MCOutput2[11]) );
  NOR2_X1 \SubCellInst_LFInst_2_LFInst_3_U5  ( .A1(PermutationOutput[11]), 
        .A2(PermutationOutput[8]), .ZN(\SubCellInst_LFInst_2_LFInst_3_n5 ) );
  NOR2_X1 \SubCellInst_LFInst_2_LFInst_3_U4  ( .A1(PermutationOutput[9]), .A2(
        \SubCellInst_LFInst_2_LFInst_3_n4 ), .ZN(
        \SubCellInst_LFInst_2_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst_LFInst_2_LFInst_3_U3  ( .A1(PermutationOutput[11]), 
        .A2(PermutationOutput[10]), .ZN(\SubCellInst_LFInst_2_LFInst_3_n4 ) );
  NOR2_X1 \SubCellInst_LFInst_3_LFInst_0_U8  ( .A1(
        \SubCellInst_LFInst_3_LFInst_0_n11 ), .A2(
        \SubCellInst_LFInst_3_LFInst_0_n10 ), .ZN(MCOutput2[12]) );
  AND2_X1 \SubCellInst_LFInst_3_LFInst_0_U7  ( .A1(PermutationOutput[15]), 
        .A2(PermutationOutput[14]), .ZN(\SubCellInst_LFInst_3_LFInst_0_n10 )
         );
  NOR2_X1 \SubCellInst_LFInst_3_LFInst_0_U6  ( .A1(PermutationOutput[13]), 
        .A2(\SubCellInst_LFInst_3_LFInst_0_n9 ), .ZN(
        \SubCellInst_LFInst_3_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst_LFInst_3_LFInst_0_U5  ( .A1(
        \SubCellInst_LFInst_3_LFInst_0_n8 ), .A2(
        \SubCellInst_LFInst_3_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_3_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst_LFInst_3_LFInst_0_U4  ( .A1(PermutationOutput[15]), 
        .A2(PermutationOutput[14]), .ZN(\SubCellInst_LFInst_3_LFInst_0_n7 ) );
  INV_X1 \SubCellInst_LFInst_3_LFInst_0_U3  ( .A(PermutationOutput[12]), .ZN(
        \SubCellInst_LFInst_3_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst_LFInst_3_LFInst_1_U6  ( .A1(
        \SubCellInst_LFInst_3_LFInst_1_n6 ), .A2(
        \SubCellInst_LFInst_3_LFInst_1_n5 ), .ZN(MCOutput2[13]) );
  NAND2_X1 \SubCellInst_LFInst_3_LFInst_1_U5  ( .A1(PermutationOutput[14]), 
        .A2(PermutationOutput[12]), .ZN(\SubCellInst_LFInst_3_LFInst_1_n5 ) );
  OR2_X1 \SubCellInst_LFInst_3_LFInst_1_U4  ( .A1(PermutationOutput[15]), .A2(
        \SubCellInst_LFInst_3_LFInst_1_n4 ), .ZN(
        \SubCellInst_LFInst_3_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst_LFInst_3_LFInst_1_U3  ( .A1(PermutationOutput[14]), 
        .A2(PermutationOutput[12]), .ZN(\SubCellInst_LFInst_3_LFInst_1_n4 ) );
  NAND2_X1 \SubCellInst_LFInst_3_LFInst_2_U8  ( .A1(
        \SubCellInst_LFInst_3_LFInst_2_n11 ), .A2(
        \SubCellInst_LFInst_3_LFInst_2_n10 ), .ZN(MCOutput2[14]) );
  OR2_X1 \SubCellInst_LFInst_3_LFInst_2_U7  ( .A1(PermutationOutput[12]), .A2(
        PermutationOutput[15]), .ZN(\SubCellInst_LFInst_3_LFInst_2_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_3_LFInst_2_U6  ( .A1(PermutationOutput[13]), 
        .A2(\SubCellInst_LFInst_3_LFInst_2_n9 ), .ZN(
        \SubCellInst_LFInst_3_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_3_LFInst_2_U5  ( .A1(
        \SubCellInst_LFInst_3_LFInst_2_n8 ), .A2(
        \SubCellInst_LFInst_3_LFInst_2_n7 ), .ZN(
        \SubCellInst_LFInst_3_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst_LFInst_3_LFInst_2_U4  ( .A1(PermutationOutput[12]), 
        .A2(PermutationOutput[15]), .ZN(\SubCellInst_LFInst_3_LFInst_2_n7 ) );
  INV_X1 \SubCellInst_LFInst_3_LFInst_2_U3  ( .A(PermutationOutput[14]), .ZN(
        \SubCellInst_LFInst_3_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst_LFInst_3_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_3_LFInst_3_n6 ), .A2(
        \SubCellInst_LFInst_3_LFInst_3_n5 ), .ZN(MCOutput2[15]) );
  NOR2_X1 \SubCellInst_LFInst_3_LFInst_3_U5  ( .A1(PermutationOutput[15]), 
        .A2(PermutationOutput[12]), .ZN(\SubCellInst_LFInst_3_LFInst_3_n5 ) );
  NOR2_X1 \SubCellInst_LFInst_3_LFInst_3_U4  ( .A1(PermutationOutput[13]), 
        .A2(\SubCellInst_LFInst_3_LFInst_3_n4 ), .ZN(
        \SubCellInst_LFInst_3_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst_LFInst_3_LFInst_3_U3  ( .A1(PermutationOutput[15]), 
        .A2(PermutationOutput[14]), .ZN(\SubCellInst_LFInst_3_LFInst_3_n4 ) );
  NOR2_X1 \SubCellInst_LFInst_4_LFInst_0_U8  ( .A1(
        \SubCellInst_LFInst_4_LFInst_0_n11 ), .A2(
        \SubCellInst_LFInst_4_LFInst_0_n10 ), .ZN(MCOutput2[16]) );
  AND2_X1 \SubCellInst_LFInst_4_LFInst_0_U7  ( .A1(PermutationOutput[19]), 
        .A2(PermutationOutput[18]), .ZN(\SubCellInst_LFInst_4_LFInst_0_n10 )
         );
  NOR2_X1 \SubCellInst_LFInst_4_LFInst_0_U6  ( .A1(PermutationOutput[17]), 
        .A2(\SubCellInst_LFInst_4_LFInst_0_n9 ), .ZN(
        \SubCellInst_LFInst_4_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst_LFInst_4_LFInst_0_U5  ( .A1(
        \SubCellInst_LFInst_4_LFInst_0_n8 ), .A2(
        \SubCellInst_LFInst_4_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_4_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst_LFInst_4_LFInst_0_U4  ( .A1(PermutationOutput[19]), 
        .A2(PermutationOutput[18]), .ZN(\SubCellInst_LFInst_4_LFInst_0_n7 ) );
  INV_X1 \SubCellInst_LFInst_4_LFInst_0_U3  ( .A(PermutationOutput[16]), .ZN(
        \SubCellInst_LFInst_4_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst_LFInst_4_LFInst_1_U6  ( .A1(
        \SubCellInst_LFInst_4_LFInst_1_n6 ), .A2(
        \SubCellInst_LFInst_4_LFInst_1_n5 ), .ZN(MCOutput2[17]) );
  NAND2_X1 \SubCellInst_LFInst_4_LFInst_1_U5  ( .A1(PermutationOutput[18]), 
        .A2(PermutationOutput[16]), .ZN(\SubCellInst_LFInst_4_LFInst_1_n5 ) );
  OR2_X1 \SubCellInst_LFInst_4_LFInst_1_U4  ( .A1(PermutationOutput[19]), .A2(
        \SubCellInst_LFInst_4_LFInst_1_n4 ), .ZN(
        \SubCellInst_LFInst_4_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst_LFInst_4_LFInst_1_U3  ( .A1(PermutationOutput[18]), 
        .A2(PermutationOutput[16]), .ZN(\SubCellInst_LFInst_4_LFInst_1_n4 ) );
  NAND2_X1 \SubCellInst_LFInst_4_LFInst_2_U8  ( .A1(
        \SubCellInst_LFInst_4_LFInst_2_n11 ), .A2(
        \SubCellInst_LFInst_4_LFInst_2_n10 ), .ZN(MCOutput2[18]) );
  OR2_X1 \SubCellInst_LFInst_4_LFInst_2_U7  ( .A1(PermutationOutput[16]), .A2(
        PermutationOutput[19]), .ZN(\SubCellInst_LFInst_4_LFInst_2_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_4_LFInst_2_U6  ( .A1(PermutationOutput[17]), 
        .A2(\SubCellInst_LFInst_4_LFInst_2_n9 ), .ZN(
        \SubCellInst_LFInst_4_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_4_LFInst_2_U5  ( .A1(
        \SubCellInst_LFInst_4_LFInst_2_n8 ), .A2(
        \SubCellInst_LFInst_4_LFInst_2_n7 ), .ZN(
        \SubCellInst_LFInst_4_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst_LFInst_4_LFInst_2_U4  ( .A1(PermutationOutput[16]), 
        .A2(PermutationOutput[19]), .ZN(\SubCellInst_LFInst_4_LFInst_2_n7 ) );
  INV_X1 \SubCellInst_LFInst_4_LFInst_2_U3  ( .A(PermutationOutput[18]), .ZN(
        \SubCellInst_LFInst_4_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst_LFInst_4_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_4_LFInst_3_n6 ), .A2(
        \SubCellInst_LFInst_4_LFInst_3_n5 ), .ZN(MCOutput2[19]) );
  NOR2_X1 \SubCellInst_LFInst_4_LFInst_3_U5  ( .A1(PermutationOutput[19]), 
        .A2(PermutationOutput[16]), .ZN(\SubCellInst_LFInst_4_LFInst_3_n5 ) );
  NOR2_X1 \SubCellInst_LFInst_4_LFInst_3_U4  ( .A1(PermutationOutput[17]), 
        .A2(\SubCellInst_LFInst_4_LFInst_3_n4 ), .ZN(
        \SubCellInst_LFInst_4_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst_LFInst_4_LFInst_3_U3  ( .A1(PermutationOutput[19]), 
        .A2(PermutationOutput[18]), .ZN(\SubCellInst_LFInst_4_LFInst_3_n4 ) );
  NOR2_X1 \SubCellInst_LFInst_5_LFInst_0_U8  ( .A1(
        \SubCellInst_LFInst_5_LFInst_0_n11 ), .A2(
        \SubCellInst_LFInst_5_LFInst_0_n10 ), .ZN(MCOutput2[20]) );
  AND2_X1 \SubCellInst_LFInst_5_LFInst_0_U7  ( .A1(PermutationOutput[23]), 
        .A2(PermutationOutput[22]), .ZN(\SubCellInst_LFInst_5_LFInst_0_n10 )
         );
  NOR2_X1 \SubCellInst_LFInst_5_LFInst_0_U6  ( .A1(PermutationOutput[21]), 
        .A2(\SubCellInst_LFInst_5_LFInst_0_n9 ), .ZN(
        \SubCellInst_LFInst_5_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst_LFInst_5_LFInst_0_U5  ( .A1(
        \SubCellInst_LFInst_5_LFInst_0_n8 ), .A2(
        \SubCellInst_LFInst_5_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_5_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst_LFInst_5_LFInst_0_U4  ( .A1(PermutationOutput[23]), 
        .A2(PermutationOutput[22]), .ZN(\SubCellInst_LFInst_5_LFInst_0_n7 ) );
  INV_X1 \SubCellInst_LFInst_5_LFInst_0_U3  ( .A(PermutationOutput[20]), .ZN(
        \SubCellInst_LFInst_5_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst_LFInst_5_LFInst_1_U6  ( .A1(
        \SubCellInst_LFInst_5_LFInst_1_n6 ), .A2(
        \SubCellInst_LFInst_5_LFInst_1_n5 ), .ZN(MCOutput2[21]) );
  NAND2_X1 \SubCellInst_LFInst_5_LFInst_1_U5  ( .A1(PermutationOutput[22]), 
        .A2(PermutationOutput[20]), .ZN(\SubCellInst_LFInst_5_LFInst_1_n5 ) );
  OR2_X1 \SubCellInst_LFInst_5_LFInst_1_U4  ( .A1(PermutationOutput[23]), .A2(
        \SubCellInst_LFInst_5_LFInst_1_n4 ), .ZN(
        \SubCellInst_LFInst_5_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst_LFInst_5_LFInst_1_U3  ( .A1(PermutationOutput[22]), 
        .A2(PermutationOutput[20]), .ZN(\SubCellInst_LFInst_5_LFInst_1_n4 ) );
  NAND2_X1 \SubCellInst_LFInst_5_LFInst_2_U8  ( .A1(
        \SubCellInst_LFInst_5_LFInst_2_n11 ), .A2(
        \SubCellInst_LFInst_5_LFInst_2_n10 ), .ZN(MCOutput2[22]) );
  OR2_X1 \SubCellInst_LFInst_5_LFInst_2_U7  ( .A1(PermutationOutput[20]), .A2(
        PermutationOutput[23]), .ZN(\SubCellInst_LFInst_5_LFInst_2_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_5_LFInst_2_U6  ( .A1(PermutationOutput[21]), 
        .A2(\SubCellInst_LFInst_5_LFInst_2_n9 ), .ZN(
        \SubCellInst_LFInst_5_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_5_LFInst_2_U5  ( .A1(
        \SubCellInst_LFInst_5_LFInst_2_n8 ), .A2(
        \SubCellInst_LFInst_5_LFInst_2_n7 ), .ZN(
        \SubCellInst_LFInst_5_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst_LFInst_5_LFInst_2_U4  ( .A1(PermutationOutput[20]), 
        .A2(PermutationOutput[23]), .ZN(\SubCellInst_LFInst_5_LFInst_2_n7 ) );
  INV_X1 \SubCellInst_LFInst_5_LFInst_2_U3  ( .A(PermutationOutput[22]), .ZN(
        \SubCellInst_LFInst_5_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst_LFInst_5_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_5_LFInst_3_n6 ), .A2(
        \SubCellInst_LFInst_5_LFInst_3_n5 ), .ZN(MCOutput2[23]) );
  NOR2_X1 \SubCellInst_LFInst_5_LFInst_3_U5  ( .A1(PermutationOutput[23]), 
        .A2(PermutationOutput[20]), .ZN(\SubCellInst_LFInst_5_LFInst_3_n5 ) );
  NOR2_X1 \SubCellInst_LFInst_5_LFInst_3_U4  ( .A1(PermutationOutput[21]), 
        .A2(\SubCellInst_LFInst_5_LFInst_3_n4 ), .ZN(
        \SubCellInst_LFInst_5_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst_LFInst_5_LFInst_3_U3  ( .A1(PermutationOutput[23]), 
        .A2(PermutationOutput[22]), .ZN(\SubCellInst_LFInst_5_LFInst_3_n4 ) );
  NOR2_X1 \SubCellInst_LFInst_6_LFInst_0_U8  ( .A1(
        \SubCellInst_LFInst_6_LFInst_0_n11 ), .A2(
        \SubCellInst_LFInst_6_LFInst_0_n10 ), .ZN(MCOutput2[24]) );
  AND2_X1 \SubCellInst_LFInst_6_LFInst_0_U7  ( .A1(PermutationOutput[27]), 
        .A2(PermutationOutput[26]), .ZN(\SubCellInst_LFInst_6_LFInst_0_n10 )
         );
  NOR2_X1 \SubCellInst_LFInst_6_LFInst_0_U6  ( .A1(PermutationOutput[25]), 
        .A2(\SubCellInst_LFInst_6_LFInst_0_n9 ), .ZN(
        \SubCellInst_LFInst_6_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst_LFInst_6_LFInst_0_U5  ( .A1(
        \SubCellInst_LFInst_6_LFInst_0_n8 ), .A2(
        \SubCellInst_LFInst_6_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_6_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst_LFInst_6_LFInst_0_U4  ( .A1(PermutationOutput[27]), 
        .A2(PermutationOutput[26]), .ZN(\SubCellInst_LFInst_6_LFInst_0_n7 ) );
  INV_X1 \SubCellInst_LFInst_6_LFInst_0_U3  ( .A(PermutationOutput[24]), .ZN(
        \SubCellInst_LFInst_6_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst_LFInst_6_LFInst_1_U6  ( .A1(
        \SubCellInst_LFInst_6_LFInst_1_n6 ), .A2(
        \SubCellInst_LFInst_6_LFInst_1_n5 ), .ZN(MCOutput2[25]) );
  NAND2_X1 \SubCellInst_LFInst_6_LFInst_1_U5  ( .A1(PermutationOutput[26]), 
        .A2(PermutationOutput[24]), .ZN(\SubCellInst_LFInst_6_LFInst_1_n5 ) );
  OR2_X1 \SubCellInst_LFInst_6_LFInst_1_U4  ( .A1(PermutationOutput[27]), .A2(
        \SubCellInst_LFInst_6_LFInst_1_n4 ), .ZN(
        \SubCellInst_LFInst_6_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst_LFInst_6_LFInst_1_U3  ( .A1(PermutationOutput[26]), 
        .A2(PermutationOutput[24]), .ZN(\SubCellInst_LFInst_6_LFInst_1_n4 ) );
  NAND2_X1 \SubCellInst_LFInst_6_LFInst_2_U8  ( .A1(
        \SubCellInst_LFInst_6_LFInst_2_n11 ), .A2(
        \SubCellInst_LFInst_6_LFInst_2_n10 ), .ZN(MCOutput2[26]) );
  OR2_X1 \SubCellInst_LFInst_6_LFInst_2_U7  ( .A1(PermutationOutput[24]), .A2(
        PermutationOutput[27]), .ZN(\SubCellInst_LFInst_6_LFInst_2_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_6_LFInst_2_U6  ( .A1(PermutationOutput[25]), 
        .A2(\SubCellInst_LFInst_6_LFInst_2_n9 ), .ZN(
        \SubCellInst_LFInst_6_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_6_LFInst_2_U5  ( .A1(
        \SubCellInst_LFInst_6_LFInst_2_n8 ), .A2(
        \SubCellInst_LFInst_6_LFInst_2_n7 ), .ZN(
        \SubCellInst_LFInst_6_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst_LFInst_6_LFInst_2_U4  ( .A1(PermutationOutput[24]), 
        .A2(PermutationOutput[27]), .ZN(\SubCellInst_LFInst_6_LFInst_2_n7 ) );
  INV_X1 \SubCellInst_LFInst_6_LFInst_2_U3  ( .A(PermutationOutput[26]), .ZN(
        \SubCellInst_LFInst_6_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst_LFInst_6_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_6_LFInst_3_n6 ), .A2(
        \SubCellInst_LFInst_6_LFInst_3_n5 ), .ZN(MCOutput2[27]) );
  NOR2_X1 \SubCellInst_LFInst_6_LFInst_3_U5  ( .A1(PermutationOutput[27]), 
        .A2(PermutationOutput[24]), .ZN(\SubCellInst_LFInst_6_LFInst_3_n5 ) );
  NOR2_X1 \SubCellInst_LFInst_6_LFInst_3_U4  ( .A1(PermutationOutput[25]), 
        .A2(\SubCellInst_LFInst_6_LFInst_3_n4 ), .ZN(
        \SubCellInst_LFInst_6_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst_LFInst_6_LFInst_3_U3  ( .A1(PermutationOutput[27]), 
        .A2(PermutationOutput[26]), .ZN(\SubCellInst_LFInst_6_LFInst_3_n4 ) );
  NOR2_X1 \SubCellInst_LFInst_7_LFInst_0_U8  ( .A1(
        \SubCellInst_LFInst_7_LFInst_0_n11 ), .A2(
        \SubCellInst_LFInst_7_LFInst_0_n10 ), .ZN(MCOutput2[28]) );
  AND2_X1 \SubCellInst_LFInst_7_LFInst_0_U7  ( .A1(PermutationOutput[31]), 
        .A2(PermutationOutput[30]), .ZN(\SubCellInst_LFInst_7_LFInst_0_n10 )
         );
  NOR2_X1 \SubCellInst_LFInst_7_LFInst_0_U6  ( .A1(PermutationOutput[29]), 
        .A2(\SubCellInst_LFInst_7_LFInst_0_n9 ), .ZN(
        \SubCellInst_LFInst_7_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst_LFInst_7_LFInst_0_U5  ( .A1(
        \SubCellInst_LFInst_7_LFInst_0_n8 ), .A2(
        \SubCellInst_LFInst_7_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_7_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst_LFInst_7_LFInst_0_U4  ( .A1(PermutationOutput[31]), 
        .A2(PermutationOutput[30]), .ZN(\SubCellInst_LFInst_7_LFInst_0_n7 ) );
  INV_X1 \SubCellInst_LFInst_7_LFInst_0_U3  ( .A(PermutationOutput[28]), .ZN(
        \SubCellInst_LFInst_7_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst_LFInst_7_LFInst_1_U6  ( .A1(
        \SubCellInst_LFInst_7_LFInst_1_n6 ), .A2(
        \SubCellInst_LFInst_7_LFInst_1_n5 ), .ZN(MCOutput2[29]) );
  NAND2_X1 \SubCellInst_LFInst_7_LFInst_1_U5  ( .A1(PermutationOutput[30]), 
        .A2(PermutationOutput[28]), .ZN(\SubCellInst_LFInst_7_LFInst_1_n5 ) );
  OR2_X1 \SubCellInst_LFInst_7_LFInst_1_U4  ( .A1(PermutationOutput[31]), .A2(
        \SubCellInst_LFInst_7_LFInst_1_n4 ), .ZN(
        \SubCellInst_LFInst_7_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst_LFInst_7_LFInst_1_U3  ( .A1(PermutationOutput[30]), 
        .A2(PermutationOutput[28]), .ZN(\SubCellInst_LFInst_7_LFInst_1_n4 ) );
  NAND2_X1 \SubCellInst_LFInst_7_LFInst_2_U8  ( .A1(
        \SubCellInst_LFInst_7_LFInst_2_n11 ), .A2(
        \SubCellInst_LFInst_7_LFInst_2_n10 ), .ZN(MCOutput2[30]) );
  OR2_X1 \SubCellInst_LFInst_7_LFInst_2_U7  ( .A1(PermutationOutput[28]), .A2(
        PermutationOutput[31]), .ZN(\SubCellInst_LFInst_7_LFInst_2_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_7_LFInst_2_U6  ( .A1(PermutationOutput[29]), 
        .A2(\SubCellInst_LFInst_7_LFInst_2_n9 ), .ZN(
        \SubCellInst_LFInst_7_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_7_LFInst_2_U5  ( .A1(
        \SubCellInst_LFInst_7_LFInst_2_n8 ), .A2(
        \SubCellInst_LFInst_7_LFInst_2_n7 ), .ZN(
        \SubCellInst_LFInst_7_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst_LFInst_7_LFInst_2_U4  ( .A1(PermutationOutput[28]), 
        .A2(PermutationOutput[31]), .ZN(\SubCellInst_LFInst_7_LFInst_2_n7 ) );
  INV_X1 \SubCellInst_LFInst_7_LFInst_2_U3  ( .A(PermutationOutput[30]), .ZN(
        \SubCellInst_LFInst_7_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst_LFInst_7_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_7_LFInst_3_n6 ), .A2(
        \SubCellInst_LFInst_7_LFInst_3_n5 ), .ZN(MCOutput2[31]) );
  NOR2_X1 \SubCellInst_LFInst_7_LFInst_3_U5  ( .A1(PermutationOutput[31]), 
        .A2(PermutationOutput[28]), .ZN(\SubCellInst_LFInst_7_LFInst_3_n5 ) );
  NOR2_X1 \SubCellInst_LFInst_7_LFInst_3_U4  ( .A1(PermutationOutput[29]), 
        .A2(\SubCellInst_LFInst_7_LFInst_3_n4 ), .ZN(
        \SubCellInst_LFInst_7_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst_LFInst_7_LFInst_3_U3  ( .A1(PermutationOutput[31]), 
        .A2(PermutationOutput[30]), .ZN(\SubCellInst_LFInst_7_LFInst_3_n4 ) );
  NOR2_X1 \SubCellInst_LFInst_8_LFInst_0_U8  ( .A1(
        \SubCellInst_LFInst_8_LFInst_0_n11 ), .A2(
        \SubCellInst_LFInst_8_LFInst_0_n10 ), .ZN(Feedback[32]) );
  AND2_X1 \SubCellInst_LFInst_8_LFInst_0_U7  ( .A1(PermutationOutput[35]), 
        .A2(PermutationOutput[34]), .ZN(\SubCellInst_LFInst_8_LFInst_0_n10 )
         );
  NOR2_X1 \SubCellInst_LFInst_8_LFInst_0_U6  ( .A1(PermutationOutput[33]), 
        .A2(\SubCellInst_LFInst_8_LFInst_0_n9 ), .ZN(
        \SubCellInst_LFInst_8_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst_LFInst_8_LFInst_0_U5  ( .A1(
        \SubCellInst_LFInst_8_LFInst_0_n8 ), .A2(
        \SubCellInst_LFInst_8_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_8_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst_LFInst_8_LFInst_0_U4  ( .A1(PermutationOutput[35]), 
        .A2(PermutationOutput[34]), .ZN(\SubCellInst_LFInst_8_LFInst_0_n7 ) );
  INV_X1 \SubCellInst_LFInst_8_LFInst_0_U3  ( .A(PermutationOutput[32]), .ZN(
        \SubCellInst_LFInst_8_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst_LFInst_8_LFInst_1_U6  ( .A1(
        \SubCellInst_LFInst_8_LFInst_1_n6 ), .A2(
        \SubCellInst_LFInst_8_LFInst_1_n5 ), .ZN(Feedback[33]) );
  NAND2_X1 \SubCellInst_LFInst_8_LFInst_1_U5  ( .A1(PermutationOutput[34]), 
        .A2(PermutationOutput[32]), .ZN(\SubCellInst_LFInst_8_LFInst_1_n5 ) );
  OR2_X1 \SubCellInst_LFInst_8_LFInst_1_U4  ( .A1(PermutationOutput[35]), .A2(
        \SubCellInst_LFInst_8_LFInst_1_n4 ), .ZN(
        \SubCellInst_LFInst_8_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst_LFInst_8_LFInst_1_U3  ( .A1(PermutationOutput[34]), 
        .A2(PermutationOutput[32]), .ZN(\SubCellInst_LFInst_8_LFInst_1_n4 ) );
  NAND2_X1 \SubCellInst_LFInst_8_LFInst_2_U8  ( .A1(
        \SubCellInst_LFInst_8_LFInst_2_n11 ), .A2(
        \SubCellInst_LFInst_8_LFInst_2_n10 ), .ZN(Feedback[34]) );
  OR2_X1 \SubCellInst_LFInst_8_LFInst_2_U7  ( .A1(PermutationOutput[32]), .A2(
        PermutationOutput[35]), .ZN(\SubCellInst_LFInst_8_LFInst_2_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_8_LFInst_2_U6  ( .A1(PermutationOutput[33]), 
        .A2(\SubCellInst_LFInst_8_LFInst_2_n9 ), .ZN(
        \SubCellInst_LFInst_8_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_8_LFInst_2_U5  ( .A1(
        \SubCellInst_LFInst_8_LFInst_2_n8 ), .A2(
        \SubCellInst_LFInst_8_LFInst_2_n7 ), .ZN(
        \SubCellInst_LFInst_8_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst_LFInst_8_LFInst_2_U4  ( .A1(PermutationOutput[32]), 
        .A2(PermutationOutput[35]), .ZN(\SubCellInst_LFInst_8_LFInst_2_n7 ) );
  INV_X1 \SubCellInst_LFInst_8_LFInst_2_U3  ( .A(PermutationOutput[34]), .ZN(
        \SubCellInst_LFInst_8_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst_LFInst_8_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_8_LFInst_3_n6 ), .A2(
        \SubCellInst_LFInst_8_LFInst_3_n5 ), .ZN(Feedback[35]) );
  NOR2_X1 \SubCellInst_LFInst_8_LFInst_3_U5  ( .A1(PermutationOutput[35]), 
        .A2(PermutationOutput[32]), .ZN(\SubCellInst_LFInst_8_LFInst_3_n5 ) );
  NOR2_X1 \SubCellInst_LFInst_8_LFInst_3_U4  ( .A1(PermutationOutput[33]), 
        .A2(\SubCellInst_LFInst_8_LFInst_3_n4 ), .ZN(
        \SubCellInst_LFInst_8_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst_LFInst_8_LFInst_3_U3  ( .A1(PermutationOutput[35]), 
        .A2(PermutationOutput[34]), .ZN(\SubCellInst_LFInst_8_LFInst_3_n4 ) );
  NOR2_X1 \SubCellInst_LFInst_9_LFInst_0_U8  ( .A1(
        \SubCellInst_LFInst_9_LFInst_0_n11 ), .A2(
        \SubCellInst_LFInst_9_LFInst_0_n10 ), .ZN(Feedback[36]) );
  AND2_X1 \SubCellInst_LFInst_9_LFInst_0_U7  ( .A1(PermutationOutput[39]), 
        .A2(PermutationOutput[38]), .ZN(\SubCellInst_LFInst_9_LFInst_0_n10 )
         );
  NOR2_X1 \SubCellInst_LFInst_9_LFInst_0_U6  ( .A1(PermutationOutput[37]), 
        .A2(\SubCellInst_LFInst_9_LFInst_0_n9 ), .ZN(
        \SubCellInst_LFInst_9_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst_LFInst_9_LFInst_0_U5  ( .A1(
        \SubCellInst_LFInst_9_LFInst_0_n8 ), .A2(
        \SubCellInst_LFInst_9_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_9_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst_LFInst_9_LFInst_0_U4  ( .A1(PermutationOutput[39]), 
        .A2(PermutationOutput[38]), .ZN(\SubCellInst_LFInst_9_LFInst_0_n7 ) );
  INV_X1 \SubCellInst_LFInst_9_LFInst_0_U3  ( .A(PermutationOutput[36]), .ZN(
        \SubCellInst_LFInst_9_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst_LFInst_9_LFInst_1_U6  ( .A1(
        \SubCellInst_LFInst_9_LFInst_1_n6 ), .A2(
        \SubCellInst_LFInst_9_LFInst_1_n5 ), .ZN(Feedback[37]) );
  NAND2_X1 \SubCellInst_LFInst_9_LFInst_1_U5  ( .A1(PermutationOutput[38]), 
        .A2(PermutationOutput[36]), .ZN(\SubCellInst_LFInst_9_LFInst_1_n5 ) );
  OR2_X1 \SubCellInst_LFInst_9_LFInst_1_U4  ( .A1(PermutationOutput[39]), .A2(
        \SubCellInst_LFInst_9_LFInst_1_n4 ), .ZN(
        \SubCellInst_LFInst_9_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst_LFInst_9_LFInst_1_U3  ( .A1(PermutationOutput[38]), 
        .A2(PermutationOutput[36]), .ZN(\SubCellInst_LFInst_9_LFInst_1_n4 ) );
  NAND2_X1 \SubCellInst_LFInst_9_LFInst_2_U8  ( .A1(
        \SubCellInst_LFInst_9_LFInst_2_n11 ), .A2(
        \SubCellInst_LFInst_9_LFInst_2_n10 ), .ZN(Feedback[38]) );
  OR2_X1 \SubCellInst_LFInst_9_LFInst_2_U7  ( .A1(PermutationOutput[36]), .A2(
        PermutationOutput[39]), .ZN(\SubCellInst_LFInst_9_LFInst_2_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_9_LFInst_2_U6  ( .A1(PermutationOutput[37]), 
        .A2(\SubCellInst_LFInst_9_LFInst_2_n9 ), .ZN(
        \SubCellInst_LFInst_9_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_9_LFInst_2_U5  ( .A1(
        \SubCellInst_LFInst_9_LFInst_2_n8 ), .A2(
        \SubCellInst_LFInst_9_LFInst_2_n7 ), .ZN(
        \SubCellInst_LFInst_9_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst_LFInst_9_LFInst_2_U4  ( .A1(PermutationOutput[36]), 
        .A2(PermutationOutput[39]), .ZN(\SubCellInst_LFInst_9_LFInst_2_n7 ) );
  INV_X1 \SubCellInst_LFInst_9_LFInst_2_U3  ( .A(PermutationOutput[38]), .ZN(
        \SubCellInst_LFInst_9_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst_LFInst_9_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_9_LFInst_3_n6 ), .A2(
        \SubCellInst_LFInst_9_LFInst_3_n5 ), .ZN(Feedback[39]) );
  NOR2_X1 \SubCellInst_LFInst_9_LFInst_3_U5  ( .A1(PermutationOutput[39]), 
        .A2(PermutationOutput[36]), .ZN(\SubCellInst_LFInst_9_LFInst_3_n5 ) );
  NOR2_X1 \SubCellInst_LFInst_9_LFInst_3_U4  ( .A1(PermutationOutput[37]), 
        .A2(\SubCellInst_LFInst_9_LFInst_3_n4 ), .ZN(
        \SubCellInst_LFInst_9_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst_LFInst_9_LFInst_3_U3  ( .A1(PermutationOutput[39]), 
        .A2(PermutationOutput[38]), .ZN(\SubCellInst_LFInst_9_LFInst_3_n4 ) );
  NOR2_X1 \SubCellInst_LFInst_10_LFInst_0_U8  ( .A1(
        \SubCellInst_LFInst_10_LFInst_0_n11 ), .A2(
        \SubCellInst_LFInst_10_LFInst_0_n10 ), .ZN(Feedback[40]) );
  AND2_X1 \SubCellInst_LFInst_10_LFInst_0_U7  ( .A1(PermutationOutput[43]), 
        .A2(PermutationOutput[42]), .ZN(\SubCellInst_LFInst_10_LFInst_0_n10 )
         );
  NOR2_X1 \SubCellInst_LFInst_10_LFInst_0_U6  ( .A1(PermutationOutput[41]), 
        .A2(\SubCellInst_LFInst_10_LFInst_0_n9 ), .ZN(
        \SubCellInst_LFInst_10_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst_LFInst_10_LFInst_0_U5  ( .A1(
        \SubCellInst_LFInst_10_LFInst_0_n8 ), .A2(
        \SubCellInst_LFInst_10_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_10_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst_LFInst_10_LFInst_0_U4  ( .A1(PermutationOutput[43]), 
        .A2(PermutationOutput[42]), .ZN(\SubCellInst_LFInst_10_LFInst_0_n7 )
         );
  INV_X1 \SubCellInst_LFInst_10_LFInst_0_U3  ( .A(PermutationOutput[40]), .ZN(
        \SubCellInst_LFInst_10_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst_LFInst_10_LFInst_1_U6  ( .A1(
        \SubCellInst_LFInst_10_LFInst_1_n6 ), .A2(
        \SubCellInst_LFInst_10_LFInst_1_n5 ), .ZN(Feedback[41]) );
  NAND2_X1 \SubCellInst_LFInst_10_LFInst_1_U5  ( .A1(PermutationOutput[42]), 
        .A2(PermutationOutput[40]), .ZN(\SubCellInst_LFInst_10_LFInst_1_n5 )
         );
  OR2_X1 \SubCellInst_LFInst_10_LFInst_1_U4  ( .A1(PermutationOutput[43]), 
        .A2(\SubCellInst_LFInst_10_LFInst_1_n4 ), .ZN(
        \SubCellInst_LFInst_10_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst_LFInst_10_LFInst_1_U3  ( .A1(PermutationOutput[42]), 
        .A2(PermutationOutput[40]), .ZN(\SubCellInst_LFInst_10_LFInst_1_n4 )
         );
  NAND2_X1 \SubCellInst_LFInst_10_LFInst_2_U8  ( .A1(
        \SubCellInst_LFInst_10_LFInst_2_n11 ), .A2(
        \SubCellInst_LFInst_10_LFInst_2_n10 ), .ZN(Feedback[42]) );
  OR2_X1 \SubCellInst_LFInst_10_LFInst_2_U7  ( .A1(PermutationOutput[40]), 
        .A2(PermutationOutput[43]), .ZN(\SubCellInst_LFInst_10_LFInst_2_n10 )
         );
  NAND2_X1 \SubCellInst_LFInst_10_LFInst_2_U6  ( .A1(PermutationOutput[41]), 
        .A2(\SubCellInst_LFInst_10_LFInst_2_n9 ), .ZN(
        \SubCellInst_LFInst_10_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_10_LFInst_2_U5  ( .A1(
        \SubCellInst_LFInst_10_LFInst_2_n8 ), .A2(
        \SubCellInst_LFInst_10_LFInst_2_n7 ), .ZN(
        \SubCellInst_LFInst_10_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst_LFInst_10_LFInst_2_U4  ( .A1(PermutationOutput[40]), 
        .A2(PermutationOutput[43]), .ZN(\SubCellInst_LFInst_10_LFInst_2_n7 )
         );
  INV_X1 \SubCellInst_LFInst_10_LFInst_2_U3  ( .A(PermutationOutput[42]), .ZN(
        \SubCellInst_LFInst_10_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst_LFInst_10_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_10_LFInst_3_n6 ), .A2(
        \SubCellInst_LFInst_10_LFInst_3_n5 ), .ZN(Feedback[43]) );
  NOR2_X1 \SubCellInst_LFInst_10_LFInst_3_U5  ( .A1(PermutationOutput[43]), 
        .A2(PermutationOutput[40]), .ZN(\SubCellInst_LFInst_10_LFInst_3_n5 )
         );
  NOR2_X1 \SubCellInst_LFInst_10_LFInst_3_U4  ( .A1(PermutationOutput[41]), 
        .A2(\SubCellInst_LFInst_10_LFInst_3_n4 ), .ZN(
        \SubCellInst_LFInst_10_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst_LFInst_10_LFInst_3_U3  ( .A1(PermutationOutput[43]), 
        .A2(PermutationOutput[42]), .ZN(\SubCellInst_LFInst_10_LFInst_3_n4 )
         );
  NOR2_X1 \SubCellInst_LFInst_11_LFInst_0_U8  ( .A1(
        \SubCellInst_LFInst_11_LFInst_0_n11 ), .A2(
        \SubCellInst_LFInst_11_LFInst_0_n10 ), .ZN(Feedback[44]) );
  AND2_X1 \SubCellInst_LFInst_11_LFInst_0_U7  ( .A1(PermutationOutput[47]), 
        .A2(PermutationOutput[46]), .ZN(\SubCellInst_LFInst_11_LFInst_0_n10 )
         );
  NOR2_X1 \SubCellInst_LFInst_11_LFInst_0_U6  ( .A1(PermutationOutput[45]), 
        .A2(\SubCellInst_LFInst_11_LFInst_0_n9 ), .ZN(
        \SubCellInst_LFInst_11_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst_LFInst_11_LFInst_0_U5  ( .A1(
        \SubCellInst_LFInst_11_LFInst_0_n8 ), .A2(
        \SubCellInst_LFInst_11_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_11_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst_LFInst_11_LFInst_0_U4  ( .A1(PermutationOutput[47]), 
        .A2(PermutationOutput[46]), .ZN(\SubCellInst_LFInst_11_LFInst_0_n7 )
         );
  INV_X1 \SubCellInst_LFInst_11_LFInst_0_U3  ( .A(PermutationOutput[44]), .ZN(
        \SubCellInst_LFInst_11_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst_LFInst_11_LFInst_1_U6  ( .A1(
        \SubCellInst_LFInst_11_LFInst_1_n6 ), .A2(
        \SubCellInst_LFInst_11_LFInst_1_n5 ), .ZN(Feedback[45]) );
  NAND2_X1 \SubCellInst_LFInst_11_LFInst_1_U5  ( .A1(PermutationOutput[46]), 
        .A2(PermutationOutput[44]), .ZN(\SubCellInst_LFInst_11_LFInst_1_n5 )
         );
  OR2_X1 \SubCellInst_LFInst_11_LFInst_1_U4  ( .A1(PermutationOutput[47]), 
        .A2(\SubCellInst_LFInst_11_LFInst_1_n4 ), .ZN(
        \SubCellInst_LFInst_11_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst_LFInst_11_LFInst_1_U3  ( .A1(PermutationOutput[46]), 
        .A2(PermutationOutput[44]), .ZN(\SubCellInst_LFInst_11_LFInst_1_n4 )
         );
  NAND2_X1 \SubCellInst_LFInst_11_LFInst_2_U8  ( .A1(
        \SubCellInst_LFInst_11_LFInst_2_n11 ), .A2(
        \SubCellInst_LFInst_11_LFInst_2_n10 ), .ZN(Feedback[46]) );
  OR2_X1 \SubCellInst_LFInst_11_LFInst_2_U7  ( .A1(PermutationOutput[44]), 
        .A2(PermutationOutput[47]), .ZN(\SubCellInst_LFInst_11_LFInst_2_n10 )
         );
  NAND2_X1 \SubCellInst_LFInst_11_LFInst_2_U6  ( .A1(PermutationOutput[45]), 
        .A2(\SubCellInst_LFInst_11_LFInst_2_n9 ), .ZN(
        \SubCellInst_LFInst_11_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_11_LFInst_2_U5  ( .A1(
        \SubCellInst_LFInst_11_LFInst_2_n8 ), .A2(
        \SubCellInst_LFInst_11_LFInst_2_n7 ), .ZN(
        \SubCellInst_LFInst_11_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst_LFInst_11_LFInst_2_U4  ( .A1(PermutationOutput[44]), 
        .A2(PermutationOutput[47]), .ZN(\SubCellInst_LFInst_11_LFInst_2_n7 )
         );
  INV_X1 \SubCellInst_LFInst_11_LFInst_2_U3  ( .A(PermutationOutput[46]), .ZN(
        \SubCellInst_LFInst_11_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst_LFInst_11_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_11_LFInst_3_n6 ), .A2(
        \SubCellInst_LFInst_11_LFInst_3_n5 ), .ZN(Feedback[47]) );
  NOR2_X1 \SubCellInst_LFInst_11_LFInst_3_U5  ( .A1(PermutationOutput[47]), 
        .A2(PermutationOutput[44]), .ZN(\SubCellInst_LFInst_11_LFInst_3_n5 )
         );
  NOR2_X1 \SubCellInst_LFInst_11_LFInst_3_U4  ( .A1(PermutationOutput[45]), 
        .A2(\SubCellInst_LFInst_11_LFInst_3_n4 ), .ZN(
        \SubCellInst_LFInst_11_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst_LFInst_11_LFInst_3_U3  ( .A1(PermutationOutput[47]), 
        .A2(PermutationOutput[46]), .ZN(\SubCellInst_LFInst_11_LFInst_3_n4 )
         );
  NOR2_X1 \SubCellInst_LFInst_12_LFInst_0_U8  ( .A1(
        \SubCellInst_LFInst_12_LFInst_0_n11 ), .A2(
        \SubCellInst_LFInst_12_LFInst_0_n10 ), .ZN(Feedback[48]) );
  AND2_X1 \SubCellInst_LFInst_12_LFInst_0_U7  ( .A1(PermutationOutput[51]), 
        .A2(PermutationOutput[50]), .ZN(\SubCellInst_LFInst_12_LFInst_0_n10 )
         );
  NOR2_X1 \SubCellInst_LFInst_12_LFInst_0_U6  ( .A1(PermutationOutput[49]), 
        .A2(\SubCellInst_LFInst_12_LFInst_0_n9 ), .ZN(
        \SubCellInst_LFInst_12_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst_LFInst_12_LFInst_0_U5  ( .A1(
        \SubCellInst_LFInst_12_LFInst_0_n8 ), .A2(
        \SubCellInst_LFInst_12_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_12_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst_LFInst_12_LFInst_0_U4  ( .A1(PermutationOutput[51]), 
        .A2(PermutationOutput[50]), .ZN(\SubCellInst_LFInst_12_LFInst_0_n7 )
         );
  INV_X1 \SubCellInst_LFInst_12_LFInst_0_U3  ( .A(PermutationOutput[48]), .ZN(
        \SubCellInst_LFInst_12_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst_LFInst_12_LFInst_1_U6  ( .A1(
        \SubCellInst_LFInst_12_LFInst_1_n6 ), .A2(
        \SubCellInst_LFInst_12_LFInst_1_n5 ), .ZN(Feedback[49]) );
  NAND2_X1 \SubCellInst_LFInst_12_LFInst_1_U5  ( .A1(PermutationOutput[50]), 
        .A2(PermutationOutput[48]), .ZN(\SubCellInst_LFInst_12_LFInst_1_n5 )
         );
  OR2_X1 \SubCellInst_LFInst_12_LFInst_1_U4  ( .A1(PermutationOutput[51]), 
        .A2(\SubCellInst_LFInst_12_LFInst_1_n4 ), .ZN(
        \SubCellInst_LFInst_12_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst_LFInst_12_LFInst_1_U3  ( .A1(PermutationOutput[50]), 
        .A2(PermutationOutput[48]), .ZN(\SubCellInst_LFInst_12_LFInst_1_n4 )
         );
  NAND2_X1 \SubCellInst_LFInst_12_LFInst_2_U8  ( .A1(
        \SubCellInst_LFInst_12_LFInst_2_n11 ), .A2(
        \SubCellInst_LFInst_12_LFInst_2_n10 ), .ZN(Feedback[50]) );
  OR2_X1 \SubCellInst_LFInst_12_LFInst_2_U7  ( .A1(PermutationOutput[48]), 
        .A2(PermutationOutput[51]), .ZN(\SubCellInst_LFInst_12_LFInst_2_n10 )
         );
  NAND2_X1 \SubCellInst_LFInst_12_LFInst_2_U6  ( .A1(PermutationOutput[49]), 
        .A2(\SubCellInst_LFInst_12_LFInst_2_n9 ), .ZN(
        \SubCellInst_LFInst_12_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_12_LFInst_2_U5  ( .A1(
        \SubCellInst_LFInst_12_LFInst_2_n8 ), .A2(
        \SubCellInst_LFInst_12_LFInst_2_n7 ), .ZN(
        \SubCellInst_LFInst_12_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst_LFInst_12_LFInst_2_U4  ( .A1(PermutationOutput[48]), 
        .A2(PermutationOutput[51]), .ZN(\SubCellInst_LFInst_12_LFInst_2_n7 )
         );
  INV_X1 \SubCellInst_LFInst_12_LFInst_2_U3  ( .A(PermutationOutput[50]), .ZN(
        \SubCellInst_LFInst_12_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst_LFInst_12_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_12_LFInst_3_n6 ), .A2(
        \SubCellInst_LFInst_12_LFInst_3_n5 ), .ZN(Feedback[51]) );
  NOR2_X1 \SubCellInst_LFInst_12_LFInst_3_U5  ( .A1(PermutationOutput[51]), 
        .A2(PermutationOutput[48]), .ZN(\SubCellInst_LFInst_12_LFInst_3_n5 )
         );
  NOR2_X1 \SubCellInst_LFInst_12_LFInst_3_U4  ( .A1(PermutationOutput[49]), 
        .A2(\SubCellInst_LFInst_12_LFInst_3_n4 ), .ZN(
        \SubCellInst_LFInst_12_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst_LFInst_12_LFInst_3_U3  ( .A1(PermutationOutput[51]), 
        .A2(PermutationOutput[50]), .ZN(\SubCellInst_LFInst_12_LFInst_3_n4 )
         );
  NOR2_X1 \SubCellInst_LFInst_13_LFInst_0_U8  ( .A1(
        \SubCellInst_LFInst_13_LFInst_0_n11 ), .A2(
        \SubCellInst_LFInst_13_LFInst_0_n10 ), .ZN(Feedback[52]) );
  AND2_X1 \SubCellInst_LFInst_13_LFInst_0_U7  ( .A1(PermutationOutput[55]), 
        .A2(PermutationOutput[54]), .ZN(\SubCellInst_LFInst_13_LFInst_0_n10 )
         );
  NOR2_X1 \SubCellInst_LFInst_13_LFInst_0_U6  ( .A1(PermutationOutput[53]), 
        .A2(\SubCellInst_LFInst_13_LFInst_0_n9 ), .ZN(
        \SubCellInst_LFInst_13_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst_LFInst_13_LFInst_0_U5  ( .A1(
        \SubCellInst_LFInst_13_LFInst_0_n8 ), .A2(
        \SubCellInst_LFInst_13_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_13_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst_LFInst_13_LFInst_0_U4  ( .A1(PermutationOutput[55]), 
        .A2(PermutationOutput[54]), .ZN(\SubCellInst_LFInst_13_LFInst_0_n7 )
         );
  INV_X1 \SubCellInst_LFInst_13_LFInst_0_U3  ( .A(PermutationOutput[52]), .ZN(
        \SubCellInst_LFInst_13_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst_LFInst_13_LFInst_1_U6  ( .A1(
        \SubCellInst_LFInst_13_LFInst_1_n6 ), .A2(
        \SubCellInst_LFInst_13_LFInst_1_n5 ), .ZN(Feedback[53]) );
  NAND2_X1 \SubCellInst_LFInst_13_LFInst_1_U5  ( .A1(PermutationOutput[54]), 
        .A2(PermutationOutput[52]), .ZN(\SubCellInst_LFInst_13_LFInst_1_n5 )
         );
  OR2_X1 \SubCellInst_LFInst_13_LFInst_1_U4  ( .A1(PermutationOutput[55]), 
        .A2(\SubCellInst_LFInst_13_LFInst_1_n4 ), .ZN(
        \SubCellInst_LFInst_13_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst_LFInst_13_LFInst_1_U3  ( .A1(PermutationOutput[54]), 
        .A2(PermutationOutput[52]), .ZN(\SubCellInst_LFInst_13_LFInst_1_n4 )
         );
  NAND2_X1 \SubCellInst_LFInst_13_LFInst_2_U8  ( .A1(
        \SubCellInst_LFInst_13_LFInst_2_n11 ), .A2(
        \SubCellInst_LFInst_13_LFInst_2_n10 ), .ZN(Feedback[54]) );
  OR2_X1 \SubCellInst_LFInst_13_LFInst_2_U7  ( .A1(PermutationOutput[52]), 
        .A2(PermutationOutput[55]), .ZN(\SubCellInst_LFInst_13_LFInst_2_n10 )
         );
  NAND2_X1 \SubCellInst_LFInst_13_LFInst_2_U6  ( .A1(PermutationOutput[53]), 
        .A2(\SubCellInst_LFInst_13_LFInst_2_n9 ), .ZN(
        \SubCellInst_LFInst_13_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_13_LFInst_2_U5  ( .A1(
        \SubCellInst_LFInst_13_LFInst_2_n8 ), .A2(
        \SubCellInst_LFInst_13_LFInst_2_n7 ), .ZN(
        \SubCellInst_LFInst_13_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst_LFInst_13_LFInst_2_U4  ( .A1(PermutationOutput[52]), 
        .A2(PermutationOutput[55]), .ZN(\SubCellInst_LFInst_13_LFInst_2_n7 )
         );
  INV_X1 \SubCellInst_LFInst_13_LFInst_2_U3  ( .A(PermutationOutput[54]), .ZN(
        \SubCellInst_LFInst_13_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst_LFInst_13_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_13_LFInst_3_n6 ), .A2(
        \SubCellInst_LFInst_13_LFInst_3_n5 ), .ZN(Feedback[55]) );
  NOR2_X1 \SubCellInst_LFInst_13_LFInst_3_U5  ( .A1(PermutationOutput[55]), 
        .A2(PermutationOutput[52]), .ZN(\SubCellInst_LFInst_13_LFInst_3_n5 )
         );
  NOR2_X1 \SubCellInst_LFInst_13_LFInst_3_U4  ( .A1(PermutationOutput[53]), 
        .A2(\SubCellInst_LFInst_13_LFInst_3_n4 ), .ZN(
        \SubCellInst_LFInst_13_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst_LFInst_13_LFInst_3_U3  ( .A1(PermutationOutput[55]), 
        .A2(PermutationOutput[54]), .ZN(\SubCellInst_LFInst_13_LFInst_3_n4 )
         );
  NOR2_X1 \SubCellInst_LFInst_14_LFInst_0_U8  ( .A1(
        \SubCellInst_LFInst_14_LFInst_0_n11 ), .A2(
        \SubCellInst_LFInst_14_LFInst_0_n10 ), .ZN(Feedback[56]) );
  AND2_X1 \SubCellInst_LFInst_14_LFInst_0_U7  ( .A1(PermutationOutput[59]), 
        .A2(PermutationOutput[58]), .ZN(\SubCellInst_LFInst_14_LFInst_0_n10 )
         );
  NOR2_X1 \SubCellInst_LFInst_14_LFInst_0_U6  ( .A1(PermutationOutput[57]), 
        .A2(\SubCellInst_LFInst_14_LFInst_0_n9 ), .ZN(
        \SubCellInst_LFInst_14_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst_LFInst_14_LFInst_0_U5  ( .A1(
        \SubCellInst_LFInst_14_LFInst_0_n8 ), .A2(
        \SubCellInst_LFInst_14_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_14_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst_LFInst_14_LFInst_0_U4  ( .A1(PermutationOutput[59]), 
        .A2(PermutationOutput[58]), .ZN(\SubCellInst_LFInst_14_LFInst_0_n7 )
         );
  INV_X1 \SubCellInst_LFInst_14_LFInst_0_U3  ( .A(PermutationOutput[56]), .ZN(
        \SubCellInst_LFInst_14_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst_LFInst_14_LFInst_1_U6  ( .A1(
        \SubCellInst_LFInst_14_LFInst_1_n6 ), .A2(
        \SubCellInst_LFInst_14_LFInst_1_n5 ), .ZN(Feedback[57]) );
  NAND2_X1 \SubCellInst_LFInst_14_LFInst_1_U5  ( .A1(PermutationOutput[58]), 
        .A2(PermutationOutput[56]), .ZN(\SubCellInst_LFInst_14_LFInst_1_n5 )
         );
  OR2_X1 \SubCellInst_LFInst_14_LFInst_1_U4  ( .A1(PermutationOutput[59]), 
        .A2(\SubCellInst_LFInst_14_LFInst_1_n4 ), .ZN(
        \SubCellInst_LFInst_14_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst_LFInst_14_LFInst_1_U3  ( .A1(PermutationOutput[58]), 
        .A2(PermutationOutput[56]), .ZN(\SubCellInst_LFInst_14_LFInst_1_n4 )
         );
  NAND2_X1 \SubCellInst_LFInst_14_LFInst_2_U8  ( .A1(
        \SubCellInst_LFInst_14_LFInst_2_n11 ), .A2(
        \SubCellInst_LFInst_14_LFInst_2_n10 ), .ZN(Feedback[58]) );
  OR2_X1 \SubCellInst_LFInst_14_LFInst_2_U7  ( .A1(PermutationOutput[56]), 
        .A2(PermutationOutput[59]), .ZN(\SubCellInst_LFInst_14_LFInst_2_n10 )
         );
  NAND2_X1 \SubCellInst_LFInst_14_LFInst_2_U6  ( .A1(PermutationOutput[57]), 
        .A2(\SubCellInst_LFInst_14_LFInst_2_n9 ), .ZN(
        \SubCellInst_LFInst_14_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_14_LFInst_2_U5  ( .A1(
        \SubCellInst_LFInst_14_LFInst_2_n8 ), .A2(
        \SubCellInst_LFInst_14_LFInst_2_n7 ), .ZN(
        \SubCellInst_LFInst_14_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst_LFInst_14_LFInst_2_U4  ( .A1(PermutationOutput[56]), 
        .A2(PermutationOutput[59]), .ZN(\SubCellInst_LFInst_14_LFInst_2_n7 )
         );
  INV_X1 \SubCellInst_LFInst_14_LFInst_2_U3  ( .A(PermutationOutput[58]), .ZN(
        \SubCellInst_LFInst_14_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst_LFInst_14_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_14_LFInst_3_n6 ), .A2(
        \SubCellInst_LFInst_14_LFInst_3_n5 ), .ZN(Feedback[59]) );
  NOR2_X1 \SubCellInst_LFInst_14_LFInst_3_U5  ( .A1(PermutationOutput[59]), 
        .A2(PermutationOutput[56]), .ZN(\SubCellInst_LFInst_14_LFInst_3_n5 )
         );
  NOR2_X1 \SubCellInst_LFInst_14_LFInst_3_U4  ( .A1(PermutationOutput[57]), 
        .A2(\SubCellInst_LFInst_14_LFInst_3_n4 ), .ZN(
        \SubCellInst_LFInst_14_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst_LFInst_14_LFInst_3_U3  ( .A1(PermutationOutput[59]), 
        .A2(PermutationOutput[58]), .ZN(\SubCellInst_LFInst_14_LFInst_3_n4 )
         );
  NOR2_X1 \SubCellInst_LFInst_15_LFInst_0_U8  ( .A1(
        \SubCellInst_LFInst_15_LFInst_0_n11 ), .A2(
        \SubCellInst_LFInst_15_LFInst_0_n10 ), .ZN(Feedback[60]) );
  AND2_X1 \SubCellInst_LFInst_15_LFInst_0_U7  ( .A1(PermutationOutput[63]), 
        .A2(PermutationOutput[62]), .ZN(\SubCellInst_LFInst_15_LFInst_0_n10 )
         );
  NOR2_X1 \SubCellInst_LFInst_15_LFInst_0_U6  ( .A1(PermutationOutput[61]), 
        .A2(\SubCellInst_LFInst_15_LFInst_0_n9 ), .ZN(
        \SubCellInst_LFInst_15_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst_LFInst_15_LFInst_0_U5  ( .A1(
        \SubCellInst_LFInst_15_LFInst_0_n8 ), .A2(
        \SubCellInst_LFInst_15_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_15_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst_LFInst_15_LFInst_0_U4  ( .A1(PermutationOutput[63]), 
        .A2(PermutationOutput[62]), .ZN(\SubCellInst_LFInst_15_LFInst_0_n7 )
         );
  INV_X1 \SubCellInst_LFInst_15_LFInst_0_U3  ( .A(PermutationOutput[60]), .ZN(
        \SubCellInst_LFInst_15_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst_LFInst_15_LFInst_1_U6  ( .A1(
        \SubCellInst_LFInst_15_LFInst_1_n6 ), .A2(
        \SubCellInst_LFInst_15_LFInst_1_n5 ), .ZN(Feedback[61]) );
  NAND2_X1 \SubCellInst_LFInst_15_LFInst_1_U5  ( .A1(PermutationOutput[62]), 
        .A2(PermutationOutput[60]), .ZN(\SubCellInst_LFInst_15_LFInst_1_n5 )
         );
  OR2_X1 \SubCellInst_LFInst_15_LFInst_1_U4  ( .A1(PermutationOutput[63]), 
        .A2(\SubCellInst_LFInst_15_LFInst_1_n4 ), .ZN(
        \SubCellInst_LFInst_15_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst_LFInst_15_LFInst_1_U3  ( .A1(PermutationOutput[62]), 
        .A2(PermutationOutput[60]), .ZN(\SubCellInst_LFInst_15_LFInst_1_n4 )
         );
  NAND2_X1 \SubCellInst_LFInst_15_LFInst_2_U8  ( .A1(
        \SubCellInst_LFInst_15_LFInst_2_n11 ), .A2(
        \SubCellInst_LFInst_15_LFInst_2_n10 ), .ZN(Feedback[62]) );
  OR2_X1 \SubCellInst_LFInst_15_LFInst_2_U7  ( .A1(PermutationOutput[60]), 
        .A2(PermutationOutput[63]), .ZN(\SubCellInst_LFInst_15_LFInst_2_n10 )
         );
  NAND2_X1 \SubCellInst_LFInst_15_LFInst_2_U6  ( .A1(PermutationOutput[61]), 
        .A2(\SubCellInst_LFInst_15_LFInst_2_n9 ), .ZN(
        \SubCellInst_LFInst_15_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_15_LFInst_2_U5  ( .A1(
        \SubCellInst_LFInst_15_LFInst_2_n8 ), .A2(
        \SubCellInst_LFInst_15_LFInst_2_n7 ), .ZN(
        \SubCellInst_LFInst_15_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst_LFInst_15_LFInst_2_U4  ( .A1(PermutationOutput[60]), 
        .A2(PermutationOutput[63]), .ZN(\SubCellInst_LFInst_15_LFInst_2_n7 )
         );
  INV_X1 \SubCellInst_LFInst_15_LFInst_2_U3  ( .A(PermutationOutput[62]), .ZN(
        \SubCellInst_LFInst_15_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst_LFInst_15_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_15_LFInst_3_n6 ), .A2(
        \SubCellInst_LFInst_15_LFInst_3_n5 ), .ZN(Feedback[63]) );
  NOR2_X1 \SubCellInst_LFInst_15_LFInst_3_U5  ( .A1(PermutationOutput[63]), 
        .A2(PermutationOutput[60]), .ZN(\SubCellInst_LFInst_15_LFInst_3_n5 )
         );
  NOR2_X1 \SubCellInst_LFInst_15_LFInst_3_U4  ( .A1(PermutationOutput[61]), 
        .A2(\SubCellInst_LFInst_15_LFInst_3_n4 ), .ZN(
        \SubCellInst_LFInst_15_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst_LFInst_15_LFInst_3_U3  ( .A1(PermutationOutput[63]), 
        .A2(PermutationOutput[62]), .ZN(\SubCellInst_LFInst_15_LFInst_3_n4 )
         );
  XNOR2_X1 \MCInst2_XOR_r0_Inst_0_U2  ( .A(\MCInst2_XOR_r0_Inst_0_n3 ), .B(
        MCOutput2[0]), .ZN(MCOutput2[48]) );
  XNOR2_X1 \MCInst2_XOR_r0_Inst_0_U1  ( .A(Feedback[48]), .B(MCOutput2[16]), 
        .ZN(\MCInst2_XOR_r0_Inst_0_n3 ) );
  XOR2_X1 \MCInst2_XOR_r1_Inst_0_U1  ( .A(Feedback[32]), .B(MCOutput2[0]), .Z(
        MCOutput2[32]) );
  XNOR2_X1 \MCInst2_XOR_r0_Inst_1_U2  ( .A(\MCInst2_XOR_r0_Inst_1_n3 ), .B(
        MCOutput2[1]), .ZN(MCOutput2[49]) );
  XNOR2_X1 \MCInst2_XOR_r0_Inst_1_U1  ( .A(Feedback[49]), .B(MCOutput2[17]), 
        .ZN(\MCInst2_XOR_r0_Inst_1_n3 ) );
  XOR2_X1 \MCInst2_XOR_r1_Inst_1_U1  ( .A(Feedback[33]), .B(MCOutput2[1]), .Z(
        MCOutput2[33]) );
  XNOR2_X1 \MCInst2_XOR_r0_Inst_2_U2  ( .A(\MCInst2_XOR_r0_Inst_2_n3 ), .B(
        MCOutput2[2]), .ZN(MCOutput2[50]) );
  XNOR2_X1 \MCInst2_XOR_r0_Inst_2_U1  ( .A(Feedback[50]), .B(MCOutput2[18]), 
        .ZN(\MCInst2_XOR_r0_Inst_2_n3 ) );
  XOR2_X1 \MCInst2_XOR_r1_Inst_2_U1  ( .A(Feedback[34]), .B(MCOutput2[2]), .Z(
        MCOutput2[34]) );
  XNOR2_X1 \MCInst2_XOR_r0_Inst_3_U2  ( .A(\MCInst2_XOR_r0_Inst_3_n3 ), .B(
        MCOutput2[3]), .ZN(MCOutput2[51]) );
  XNOR2_X1 \MCInst2_XOR_r0_Inst_3_U1  ( .A(Feedback[51]), .B(MCOutput2[19]), 
        .ZN(\MCInst2_XOR_r0_Inst_3_n3 ) );
  XOR2_X1 \MCInst2_XOR_r1_Inst_3_U1  ( .A(Feedback[35]), .B(MCOutput2[3]), .Z(
        MCOutput2[35]) );
  XNOR2_X1 \MCInst2_XOR_r0_Inst_4_U2  ( .A(\MCInst2_XOR_r0_Inst_4_n3 ), .B(
        MCOutput2[4]), .ZN(MCOutput2[52]) );
  XNOR2_X1 \MCInst2_XOR_r0_Inst_4_U1  ( .A(Feedback[52]), .B(MCOutput2[20]), 
        .ZN(\MCInst2_XOR_r0_Inst_4_n3 ) );
  XOR2_X1 \MCInst2_XOR_r1_Inst_4_U1  ( .A(Feedback[36]), .B(MCOutput2[4]), .Z(
        MCOutput2[36]) );
  XNOR2_X1 \MCInst2_XOR_r0_Inst_5_U2  ( .A(\MCInst2_XOR_r0_Inst_5_n3 ), .B(
        MCOutput2[5]), .ZN(MCOutput2[53]) );
  XNOR2_X1 \MCInst2_XOR_r0_Inst_5_U1  ( .A(Feedback[53]), .B(MCOutput2[21]), 
        .ZN(\MCInst2_XOR_r0_Inst_5_n3 ) );
  XOR2_X1 \MCInst2_XOR_r1_Inst_5_U1  ( .A(Feedback[37]), .B(MCOutput2[5]), .Z(
        MCOutput2[37]) );
  XNOR2_X1 \MCInst2_XOR_r0_Inst_6_U2  ( .A(\MCInst2_XOR_r0_Inst_6_n3 ), .B(
        MCOutput2[6]), .ZN(MCOutput2[54]) );
  XNOR2_X1 \MCInst2_XOR_r0_Inst_6_U1  ( .A(Feedback[54]), .B(MCOutput2[22]), 
        .ZN(\MCInst2_XOR_r0_Inst_6_n3 ) );
  XOR2_X1 \MCInst2_XOR_r1_Inst_6_U1  ( .A(Feedback[38]), .B(MCOutput2[6]), .Z(
        MCOutput2[38]) );
  XNOR2_X1 \MCInst2_XOR_r0_Inst_7_U2  ( .A(\MCInst2_XOR_r0_Inst_7_n3 ), .B(
        MCOutput2[7]), .ZN(MCOutput2[55]) );
  XNOR2_X1 \MCInst2_XOR_r0_Inst_7_U1  ( .A(Feedback[55]), .B(MCOutput2[23]), 
        .ZN(\MCInst2_XOR_r0_Inst_7_n3 ) );
  XOR2_X1 \MCInst2_XOR_r1_Inst_7_U1  ( .A(Feedback[39]), .B(MCOutput2[7]), .Z(
        MCOutput2[39]) );
  XNOR2_X1 \MCInst2_XOR_r0_Inst_8_U2  ( .A(\MCInst2_XOR_r0_Inst_8_n3 ), .B(
        MCOutput2[8]), .ZN(MCOutput2[56]) );
  XNOR2_X1 \MCInst2_XOR_r0_Inst_8_U1  ( .A(Feedback[56]), .B(MCOutput2[24]), 
        .ZN(\MCInst2_XOR_r0_Inst_8_n3 ) );
  XOR2_X1 \MCInst2_XOR_r1_Inst_8_U1  ( .A(Feedback[40]), .B(MCOutput2[8]), .Z(
        MCOutput2[40]) );
  XNOR2_X1 \MCInst2_XOR_r0_Inst_9_U2  ( .A(\MCInst2_XOR_r0_Inst_9_n3 ), .B(
        MCOutput2[9]), .ZN(MCOutput2[57]) );
  XNOR2_X1 \MCInst2_XOR_r0_Inst_9_U1  ( .A(Feedback[57]), .B(MCOutput2[25]), 
        .ZN(\MCInst2_XOR_r0_Inst_9_n3 ) );
  XOR2_X1 \MCInst2_XOR_r1_Inst_9_U1  ( .A(Feedback[41]), .B(MCOutput2[9]), .Z(
        MCOutput2[41]) );
  XNOR2_X1 \MCInst2_XOR_r0_Inst_10_U2  ( .A(\MCInst2_XOR_r0_Inst_10_n3 ), .B(
        MCOutput2[10]), .ZN(MCOutput2[58]) );
  XNOR2_X1 \MCInst2_XOR_r0_Inst_10_U1  ( .A(Feedback[58]), .B(MCOutput2[26]), 
        .ZN(\MCInst2_XOR_r0_Inst_10_n3 ) );
  XOR2_X1 \MCInst2_XOR_r1_Inst_10_U1  ( .A(Feedback[42]), .B(MCOutput2[10]), 
        .Z(MCOutput2[42]) );
  XNOR2_X1 \MCInst2_XOR_r0_Inst_11_U2  ( .A(\MCInst2_XOR_r0_Inst_11_n3 ), .B(
        MCOutput2[11]), .ZN(MCOutput2[59]) );
  XNOR2_X1 \MCInst2_XOR_r0_Inst_11_U1  ( .A(Feedback[59]), .B(MCOutput2[27]), 
        .ZN(\MCInst2_XOR_r0_Inst_11_n3 ) );
  XOR2_X1 \MCInst2_XOR_r1_Inst_11_U1  ( .A(Feedback[43]), .B(MCOutput2[11]), 
        .Z(MCOutput2[43]) );
  XNOR2_X1 \MCInst2_XOR_r0_Inst_12_U2  ( .A(\MCInst2_XOR_r0_Inst_12_n3 ), .B(
        MCOutput2[12]), .ZN(MCOutput2[60]) );
  XNOR2_X1 \MCInst2_XOR_r0_Inst_12_U1  ( .A(Feedback[60]), .B(MCOutput2[28]), 
        .ZN(\MCInst2_XOR_r0_Inst_12_n3 ) );
  XOR2_X1 \MCInst2_XOR_r1_Inst_12_U1  ( .A(Feedback[44]), .B(MCOutput2[12]), 
        .Z(MCOutput2[44]) );
  XNOR2_X1 \MCInst2_XOR_r0_Inst_13_U2  ( .A(\MCInst2_XOR_r0_Inst_13_n3 ), .B(
        MCOutput2[13]), .ZN(MCOutput2[61]) );
  XNOR2_X1 \MCInst2_XOR_r0_Inst_13_U1  ( .A(Feedback[61]), .B(MCOutput2[29]), 
        .ZN(\MCInst2_XOR_r0_Inst_13_n3 ) );
  XOR2_X1 \MCInst2_XOR_r1_Inst_13_U1  ( .A(Feedback[45]), .B(MCOutput2[13]), 
        .Z(MCOutput2[45]) );
  XNOR2_X1 \MCInst2_XOR_r0_Inst_14_U2  ( .A(\MCInst2_XOR_r0_Inst_14_n3 ), .B(
        MCOutput2[14]), .ZN(MCOutput2[62]) );
  XNOR2_X1 \MCInst2_XOR_r0_Inst_14_U1  ( .A(Feedback[62]), .B(MCOutput2[30]), 
        .ZN(\MCInst2_XOR_r0_Inst_14_n3 ) );
  XOR2_X1 \MCInst2_XOR_r1_Inst_14_U1  ( .A(Feedback[46]), .B(MCOutput2[14]), 
        .Z(MCOutput2[46]) );
  XNOR2_X1 \MCInst2_XOR_r0_Inst_15_U2  ( .A(\MCInst2_XOR_r0_Inst_15_n3 ), .B(
        MCOutput2[15]), .ZN(MCOutput2[63]) );
  XNOR2_X1 \MCInst2_XOR_r0_Inst_15_U1  ( .A(Feedback[63]), .B(MCOutput2[31]), 
        .ZN(\MCInst2_XOR_r0_Inst_15_n3 ) );
  XOR2_X1 \MCInst2_XOR_r1_Inst_15_U1  ( .A(Feedback[47]), .B(MCOutput2[15]), 
        .Z(MCOutput2[47]) );
  XOR2_X1 \AddKeyXOR12_XORInst_0_0_U1  ( .A(MCOutput2[48]), .B(Key[112]), .Z(
        AddRoundKeyOutput2[48]) );
  XOR2_X1 \AddKeyXOR12_XORInst_0_1_U1  ( .A(MCOutput2[49]), .B(Key[113]), .Z(
        AddRoundKeyOutput2[49]) );
  XOR2_X1 \AddKeyXOR12_XORInst_0_2_U1  ( .A(MCOutput2[50]), .B(Key[114]), .Z(
        AddRoundKeyOutput2[50]) );
  XOR2_X1 \AddKeyXOR12_XORInst_0_3_U1  ( .A(MCOutput2[51]), .B(Key[115]), .Z(
        AddRoundKeyOutput2[51]) );
  XOR2_X1 \AddKeyXOR12_XORInst_1_0_U1  ( .A(MCOutput2[52]), .B(Key[116]), .Z(
        AddRoundKeyOutput2[52]) );
  XOR2_X1 \AddKeyXOR12_XORInst_1_1_U1  ( .A(MCOutput2[53]), .B(Key[117]), .Z(
        AddRoundKeyOutput2[53]) );
  XOR2_X1 \AddKeyXOR12_XORInst_1_2_U1  ( .A(MCOutput2[54]), .B(Key[118]), .Z(
        AddRoundKeyOutput2[54]) );
  XOR2_X1 \AddKeyXOR12_XORInst_1_3_U1  ( .A(MCOutput2[55]), .B(Key[119]), .Z(
        AddRoundKeyOutput2[55]) );
  XOR2_X1 \AddKeyXOR12_XORInst_2_0_U1  ( .A(MCOutput2[56]), .B(Key[120]), .Z(
        AddRoundKeyOutput2[56]) );
  XOR2_X1 \AddKeyXOR12_XORInst_2_1_U1  ( .A(MCOutput2[57]), .B(Key[121]), .Z(
        AddRoundKeyOutput2[57]) );
  XOR2_X1 \AddKeyXOR12_XORInst_2_2_U1  ( .A(MCOutput2[58]), .B(Key[122]), .Z(
        AddRoundKeyOutput2[58]) );
  XOR2_X1 \AddKeyXOR12_XORInst_2_3_U1  ( .A(MCOutput2[59]), .B(Key[123]), .Z(
        AddRoundKeyOutput2[59]) );
  XOR2_X1 \AddKeyXOR12_XORInst_3_0_U1  ( .A(MCOutput2[60]), .B(Key[124]), .Z(
        AddRoundKeyOutput2[60]) );
  XOR2_X1 \AddKeyXOR12_XORInst_3_1_U1  ( .A(MCOutput2[61]), .B(Key[125]), .Z(
        AddRoundKeyOutput2[61]) );
  XOR2_X1 \AddKeyXOR12_XORInst_3_2_U1  ( .A(MCOutput2[62]), .B(Key[126]), .Z(
        AddRoundKeyOutput2[62]) );
  XOR2_X1 \AddKeyXOR12_XORInst_3_3_U1  ( .A(MCOutput2[63]), .B(Key[127]), .Z(
        AddRoundKeyOutput2[63]) );
  XOR2_X1 \AddKeyConstXOR2_XORInst_0_0_U1  ( .A(Key[104]), .B(MCOutput2[40]), 
        .Z(AddRoundKeyOutput2[40]) );
  XOR2_X1 \AddKeyConstXOR2_XORInst_0_1_U1  ( .A(Key[105]), .B(MCOutput2[41]), 
        .Z(AddRoundKeyOutput2[41]) );
  XOR2_X1 \AddKeyConstXOR2_XORInst_0_2_U1  ( .A(Key[106]), .B(MCOutput2[42]), 
        .Z(AddRoundKeyOutput2[42]) );
  XOR2_X1 \AddKeyConstXOR2_XORInst_0_3_U1  ( .A(Key[107]), .B(MCOutput2[43]), 
        .Z(AddRoundKeyOutput2[43]) );
  XOR2_X1 \AddKeyConstXOR2_XORInst_1_0_U1  ( .A(Key[108]), .B(MCOutput2[44]), 
        .Z(AddRoundKeyOutput2[44]) );
  XOR2_X1 \AddKeyConstXOR2_XORInst_1_1_U1  ( .A(Key[109]), .B(MCOutput2[45]), 
        .Z(AddRoundKeyOutput2[45]) );
  XOR2_X1 \AddKeyConstXOR2_XORInst_1_2_U1  ( .A(Key[110]), .B(MCOutput2[46]), 
        .Z(AddRoundKeyOutput2[46]) );
  XOR2_X1 \AddKeyConstXOR2_XORInst_1_3_U1  ( .A(Key[111]), .B(MCOutput2[47]), 
        .Z(AddRoundKeyOutput2[47]) );
  XOR2_X1 \AddKeyXOR22_XORInst_0_0_U1  ( .A(MCOutput2[0]), .B(Key[64]), .Z(
        AddRoundKeyOutput2[0]) );
  XOR2_X1 \AddKeyXOR22_XORInst_0_1_U1  ( .A(MCOutput2[1]), .B(Key[65]), .Z(
        AddRoundKeyOutput2[1]) );
  XOR2_X1 \AddKeyXOR22_XORInst_0_2_U1  ( .A(MCOutput2[2]), .B(Key[66]), .Z(
        AddRoundKeyOutput2[2]) );
  XOR2_X1 \AddKeyXOR22_XORInst_0_3_U1  ( .A(MCOutput2[3]), .B(Key[67]), .Z(
        AddRoundKeyOutput2[3]) );
  XOR2_X1 \AddKeyXOR22_XORInst_1_0_U1  ( .A(MCOutput2[4]), .B(Key[68]), .Z(
        AddRoundKeyOutput2[4]) );
  XOR2_X1 \AddKeyXOR22_XORInst_1_1_U1  ( .A(MCOutput2[5]), .B(Key[69]), .Z(
        AddRoundKeyOutput2[5]) );
  XOR2_X1 \AddKeyXOR22_XORInst_1_2_U1  ( .A(MCOutput2[6]), .B(Key[70]), .Z(
        AddRoundKeyOutput2[6]) );
  XOR2_X1 \AddKeyXOR22_XORInst_1_3_U1  ( .A(MCOutput2[7]), .B(Key[71]), .Z(
        AddRoundKeyOutput2[7]) );
  XOR2_X1 \AddKeyXOR22_XORInst_2_0_U1  ( .A(MCOutput2[8]), .B(Key[72]), .Z(
        AddRoundKeyOutput2[8]) );
  XOR2_X1 \AddKeyXOR22_XORInst_2_1_U1  ( .A(MCOutput2[9]), .B(Key[73]), .Z(
        AddRoundKeyOutput2[9]) );
  XOR2_X1 \AddKeyXOR22_XORInst_2_2_U1  ( .A(MCOutput2[10]), .B(Key[74]), .Z(
        AddRoundKeyOutput2[10]) );
  XOR2_X1 \AddKeyXOR22_XORInst_2_3_U1  ( .A(MCOutput2[11]), .B(Key[75]), .Z(
        AddRoundKeyOutput2[11]) );
  XOR2_X1 \AddKeyXOR22_XORInst_3_0_U1  ( .A(MCOutput2[12]), .B(Key[76]), .Z(
        AddRoundKeyOutput2[12]) );
  XOR2_X1 \AddKeyXOR22_XORInst_3_1_U1  ( .A(MCOutput2[13]), .B(Key[77]), .Z(
        AddRoundKeyOutput2[13]) );
  XOR2_X1 \AddKeyXOR22_XORInst_3_2_U1  ( .A(MCOutput2[14]), .B(Key[78]), .Z(
        AddRoundKeyOutput2[14]) );
  XOR2_X1 \AddKeyXOR22_XORInst_3_3_U1  ( .A(MCOutput2[15]), .B(Key[79]), .Z(
        AddRoundKeyOutput2[15]) );
  XOR2_X1 \AddKeyXOR22_XORInst_4_0_U1  ( .A(MCOutput2[16]), .B(Key[80]), .Z(
        AddRoundKeyOutput2[16]) );
  XOR2_X1 \AddKeyXOR22_XORInst_4_1_U1  ( .A(MCOutput2[17]), .B(Key[81]), .Z(
        AddRoundKeyOutput2[17]) );
  XOR2_X1 \AddKeyXOR22_XORInst_4_2_U1  ( .A(MCOutput2[18]), .B(Key[82]), .Z(
        AddRoundKeyOutput2[18]) );
  XOR2_X1 \AddKeyXOR22_XORInst_4_3_U1  ( .A(MCOutput2[19]), .B(Key[83]), .Z(
        AddRoundKeyOutput2[19]) );
  XOR2_X1 \AddKeyXOR22_XORInst_5_0_U1  ( .A(MCOutput2[20]), .B(Key[84]), .Z(
        AddRoundKeyOutput2[20]) );
  XOR2_X1 \AddKeyXOR22_XORInst_5_1_U1  ( .A(MCOutput2[21]), .B(Key[85]), .Z(
        AddRoundKeyOutput2[21]) );
  XOR2_X1 \AddKeyXOR22_XORInst_5_2_U1  ( .A(MCOutput2[22]), .B(Key[86]), .Z(
        AddRoundKeyOutput2[22]) );
  XOR2_X1 \AddKeyXOR22_XORInst_5_3_U1  ( .A(MCOutput2[23]), .B(Key[87]), .Z(
        AddRoundKeyOutput2[23]) );
  XOR2_X1 \AddKeyXOR22_XORInst_6_0_U1  ( .A(MCOutput2[24]), .B(Key[88]), .Z(
        AddRoundKeyOutput2[24]) );
  XOR2_X1 \AddKeyXOR22_XORInst_6_1_U1  ( .A(MCOutput2[25]), .B(Key[89]), .Z(
        AddRoundKeyOutput2[25]) );
  XOR2_X1 \AddKeyXOR22_XORInst_6_2_U1  ( .A(MCOutput2[26]), .B(Key[90]), .Z(
        AddRoundKeyOutput2[26]) );
  XOR2_X1 \AddKeyXOR22_XORInst_6_3_U1  ( .A(MCOutput2[27]), .B(Key[91]), .Z(
        AddRoundKeyOutput2[27]) );
  XOR2_X1 \AddKeyXOR22_XORInst_7_0_U1  ( .A(MCOutput2[28]), .B(Key[92]), .Z(
        AddRoundKeyOutput2[28]) );
  XOR2_X1 \AddKeyXOR22_XORInst_7_1_U1  ( .A(MCOutput2[29]), .B(Key[93]), .Z(
        AddRoundKeyOutput2[29]) );
  XOR2_X1 \AddKeyXOR22_XORInst_7_2_U1  ( .A(MCOutput2[30]), .B(Key[94]), .Z(
        AddRoundKeyOutput2[30]) );
  XOR2_X1 \AddKeyXOR22_XORInst_7_3_U1  ( .A(MCOutput2[31]), .B(Key[95]), .Z(
        AddRoundKeyOutput2[31]) );
  XOR2_X1 \AddKeyXOR22_XORInst_8_0_U1  ( .A(MCOutput2[32]), .B(Key[96]), .Z(
        AddRoundKeyOutput2[32]) );
  XOR2_X1 \AddKeyXOR22_XORInst_8_1_U1  ( .A(MCOutput2[33]), .B(Key[97]), .Z(
        AddRoundKeyOutput2[33]) );
  XOR2_X1 \AddKeyXOR22_XORInst_8_2_U1  ( .A(MCOutput2[34]), .B(Key[98]), .Z(
        AddRoundKeyOutput2[34]) );
  XOR2_X1 \AddKeyXOR22_XORInst_8_3_U1  ( .A(MCOutput2[35]), .B(Key[99]), .Z(
        AddRoundKeyOutput2[35]) );
  XOR2_X1 \AddKeyXOR22_XORInst_9_0_U1  ( .A(MCOutput2[36]), .B(Key[100]), .Z(
        AddRoundKeyOutput2[36]) );
  XOR2_X1 \AddKeyXOR22_XORInst_9_1_U1  ( .A(MCOutput2[37]), .B(Key[101]), .Z(
        AddRoundKeyOutput2[37]) );
  XOR2_X1 \AddKeyXOR22_XORInst_9_2_U1  ( .A(MCOutput2[38]), .B(Key[102]), .Z(
        AddRoundKeyOutput2[38]) );
  XOR2_X1 \AddKeyXOR22_XORInst_9_3_U1  ( .A(MCOutput2[39]), .B(Key[103]), .Z(
        AddRoundKeyOutput2[39]) );
  DFF_X1 \StateReg2_s_current_state_reg[0]  ( .D(AddRoundKeyOutput2[0]), .CK(
        clk), .Q(PermutationOutput2[60]) );
  DFF_X1 \StateReg2_s_current_state_reg[1]  ( .D(AddRoundKeyOutput2[1]), .CK(
        clk), .Q(PermutationOutput2[61]) );
  DFF_X1 \StateReg2_s_current_state_reg[2]  ( .D(AddRoundKeyOutput2[2]), .CK(
        clk), .Q(PermutationOutput2[62]) );
  DFF_X1 \StateReg2_s_current_state_reg[3]  ( .D(AddRoundKeyOutput2[3]), .CK(
        clk), .Q(PermutationOutput2[63]) );
  DFF_X1 \StateReg2_s_current_state_reg[4]  ( .D(AddRoundKeyOutput2[4]), .CK(
        clk), .Q(PermutationOutput2[48]) );
  DFF_X1 \StateReg2_s_current_state_reg[5]  ( .D(AddRoundKeyOutput2[5]), .CK(
        clk), .Q(PermutationOutput2[49]) );
  DFF_X1 \StateReg2_s_current_state_reg[6]  ( .D(AddRoundKeyOutput2[6]), .CK(
        clk), .Q(PermutationOutput2[50]) );
  DFF_X1 \StateReg2_s_current_state_reg[7]  ( .D(AddRoundKeyOutput2[7]), .CK(
        clk), .Q(PermutationOutput2[51]) );
  DFF_X1 \StateReg2_s_current_state_reg[8]  ( .D(AddRoundKeyOutput2[8]), .CK(
        clk), .Q(PermutationOutput2[52]) );
  DFF_X1 \StateReg2_s_current_state_reg[9]  ( .D(AddRoundKeyOutput2[9]), .CK(
        clk), .Q(PermutationOutput2[53]) );
  DFF_X1 \StateReg2_s_current_state_reg[10]  ( .D(AddRoundKeyOutput2[10]), 
        .CK(clk), .Q(PermutationOutput2[54]) );
  DFF_X1 \StateReg2_s_current_state_reg[11]  ( .D(AddRoundKeyOutput2[11]), 
        .CK(clk), .Q(PermutationOutput2[55]) );
  DFF_X1 \StateReg2_s_current_state_reg[12]  ( .D(AddRoundKeyOutput2[12]), 
        .CK(clk), .Q(PermutationOutput2[56]) );
  DFF_X1 \StateReg2_s_current_state_reg[13]  ( .D(AddRoundKeyOutput2[13]), 
        .CK(clk), .Q(PermutationOutput2[57]) );
  DFF_X1 \StateReg2_s_current_state_reg[14]  ( .D(AddRoundKeyOutput2[14]), 
        .CK(clk), .Q(PermutationOutput2[58]) );
  DFF_X1 \StateReg2_s_current_state_reg[15]  ( .D(AddRoundKeyOutput2[15]), 
        .CK(clk), .Q(PermutationOutput2[59]) );
  DFF_X1 \StateReg2_s_current_state_reg[16]  ( .D(AddRoundKeyOutput2[16]), 
        .CK(clk), .Q(PermutationOutput2[32]) );
  DFF_X1 \StateReg2_s_current_state_reg[17]  ( .D(AddRoundKeyOutput2[17]), 
        .CK(clk), .Q(PermutationOutput2[33]) );
  DFF_X1 \StateReg2_s_current_state_reg[18]  ( .D(AddRoundKeyOutput2[18]), 
        .CK(clk), .Q(PermutationOutput2[34]) );
  DFF_X1 \StateReg2_s_current_state_reg[19]  ( .D(AddRoundKeyOutput2[19]), 
        .CK(clk), .Q(PermutationOutput2[35]) );
  DFF_X1 \StateReg2_s_current_state_reg[20]  ( .D(AddRoundKeyOutput2[20]), 
        .CK(clk), .Q(PermutationOutput2[44]) );
  DFF_X1 \StateReg2_s_current_state_reg[21]  ( .D(AddRoundKeyOutput2[21]), 
        .CK(clk), .Q(PermutationOutput2[45]) );
  DFF_X1 \StateReg2_s_current_state_reg[22]  ( .D(AddRoundKeyOutput2[22]), 
        .CK(clk), .Q(PermutationOutput2[46]) );
  DFF_X1 \StateReg2_s_current_state_reg[23]  ( .D(AddRoundKeyOutput2[23]), 
        .CK(clk), .Q(PermutationOutput2[47]) );
  DFF_X1 \StateReg2_s_current_state_reg[24]  ( .D(AddRoundKeyOutput2[24]), 
        .CK(clk), .Q(PermutationOutput2[40]) );
  DFF_X1 \StateReg2_s_current_state_reg[25]  ( .D(AddRoundKeyOutput2[25]), 
        .CK(clk), .Q(PermutationOutput2[41]) );
  DFF_X1 \StateReg2_s_current_state_reg[26]  ( .D(AddRoundKeyOutput2[26]), 
        .CK(clk), .Q(PermutationOutput2[42]) );
  DFF_X1 \StateReg2_s_current_state_reg[27]  ( .D(AddRoundKeyOutput2[27]), 
        .CK(clk), .Q(PermutationOutput2[43]) );
  DFF_X1 \StateReg2_s_current_state_reg[28]  ( .D(AddRoundKeyOutput2[28]), 
        .CK(clk), .Q(PermutationOutput2[36]) );
  DFF_X1 \StateReg2_s_current_state_reg[29]  ( .D(AddRoundKeyOutput2[29]), 
        .CK(clk), .Q(PermutationOutput2[37]) );
  DFF_X1 \StateReg2_s_current_state_reg[30]  ( .D(AddRoundKeyOutput2[30]), 
        .CK(clk), .Q(PermutationOutput2[38]) );
  DFF_X1 \StateReg2_s_current_state_reg[31]  ( .D(AddRoundKeyOutput2[31]), 
        .CK(clk), .Q(PermutationOutput2[39]) );
  DFF_X1 \StateReg2_s_current_state_reg[32]  ( .D(AddRoundKeyOutput2[32]), 
        .CK(clk), .Q(PermutationOutput2[16]) );
  DFF_X1 \StateReg2_s_current_state_reg[33]  ( .D(AddRoundKeyOutput2[33]), 
        .CK(clk), .Q(PermutationOutput2[17]) );
  DFF_X1 \StateReg2_s_current_state_reg[34]  ( .D(AddRoundKeyOutput2[34]), 
        .CK(clk), .Q(PermutationOutput2[18]) );
  DFF_X1 \StateReg2_s_current_state_reg[35]  ( .D(AddRoundKeyOutput2[35]), 
        .CK(clk), .Q(PermutationOutput2[19]) );
  DFF_X1 \StateReg2_s_current_state_reg[36]  ( .D(AddRoundKeyOutput2[36]), 
        .CK(clk), .Q(PermutationOutput2[28]) );
  DFF_X1 \StateReg2_s_current_state_reg[37]  ( .D(AddRoundKeyOutput2[37]), 
        .CK(clk), .Q(PermutationOutput2[29]) );
  DFF_X1 \StateReg2_s_current_state_reg[38]  ( .D(AddRoundKeyOutput2[38]), 
        .CK(clk), .Q(PermutationOutput2[30]) );
  DFF_X1 \StateReg2_s_current_state_reg[39]  ( .D(AddRoundKeyOutput2[39]), 
        .CK(clk), .Q(PermutationOutput2[31]) );
  DFF_X1 \StateReg2_s_current_state_reg[40]  ( .D(AddRoundKeyOutput2[40]), 
        .CK(clk), .Q(PermutationOutput2[24]) );
  DFF_X1 \StateReg2_s_current_state_reg[41]  ( .D(AddRoundKeyOutput2[41]), 
        .CK(clk), .Q(PermutationOutput2[25]) );
  DFF_X1 \StateReg2_s_current_state_reg[42]  ( .D(AddRoundKeyOutput2[42]), 
        .CK(clk), .Q(PermutationOutput2[26]) );
  DFF_X1 \StateReg2_s_current_state_reg[43]  ( .D(AddRoundKeyOutput2[43]), 
        .CK(clk), .Q(PermutationOutput2[27]) );
  DFF_X1 \StateReg2_s_current_state_reg[44]  ( .D(AddRoundKeyOutput2[44]), 
        .CK(clk), .Q(PermutationOutput2[20]) );
  DFF_X1 \StateReg2_s_current_state_reg[45]  ( .D(AddRoundKeyOutput2[45]), 
        .CK(clk), .Q(PermutationOutput2[21]) );
  DFF_X1 \StateReg2_s_current_state_reg[46]  ( .D(AddRoundKeyOutput2[46]), 
        .CK(clk), .Q(PermutationOutput2[22]) );
  DFF_X1 \StateReg2_s_current_state_reg[47]  ( .D(AddRoundKeyOutput2[47]), 
        .CK(clk), .Q(PermutationOutput2[23]) );
  DFF_X1 \StateReg2_s_current_state_reg[48]  ( .D(AddRoundKeyOutput2[48]), 
        .CK(clk), .Q(PermutationOutput2[4]) );
  DFF_X1 \StateReg2_s_current_state_reg[49]  ( .D(AddRoundKeyOutput2[49]), 
        .CK(clk), .Q(PermutationOutput2[5]) );
  DFF_X1 \StateReg2_s_current_state_reg[50]  ( .D(AddRoundKeyOutput2[50]), 
        .CK(clk), .Q(PermutationOutput2[6]) );
  DFF_X1 \StateReg2_s_current_state_reg[51]  ( .D(AddRoundKeyOutput2[51]), 
        .CK(clk), .Q(PermutationOutput2[7]) );
  DFF_X1 \StateReg2_s_current_state_reg[52]  ( .D(AddRoundKeyOutput2[52]), 
        .CK(clk), .Q(PermutationOutput2[8]) );
  DFF_X1 \StateReg2_s_current_state_reg[53]  ( .D(AddRoundKeyOutput2[53]), 
        .CK(clk), .Q(PermutationOutput2[9]) );
  DFF_X1 \StateReg2_s_current_state_reg[54]  ( .D(AddRoundKeyOutput2[54]), 
        .CK(clk), .Q(PermutationOutput2[10]) );
  DFF_X1 \StateReg2_s_current_state_reg[55]  ( .D(AddRoundKeyOutput2[55]), 
        .CK(clk), .Q(PermutationOutput2[11]) );
  DFF_X1 \StateReg2_s_current_state_reg[56]  ( .D(AddRoundKeyOutput2[56]), 
        .CK(clk), .Q(PermutationOutput2[12]) );
  DFF_X1 \StateReg2_s_current_state_reg[57]  ( .D(AddRoundKeyOutput2[57]), 
        .CK(clk), .Q(PermutationOutput2[13]) );
  DFF_X1 \StateReg2_s_current_state_reg[58]  ( .D(AddRoundKeyOutput2[58]), 
        .CK(clk), .Q(PermutationOutput2[14]) );
  DFF_X1 \StateReg2_s_current_state_reg[59]  ( .D(AddRoundKeyOutput2[59]), 
        .CK(clk), .Q(PermutationOutput2[15]) );
  DFF_X1 \StateReg2_s_current_state_reg[60]  ( .D(AddRoundKeyOutput2[60]), 
        .CK(clk), .Q(PermutationOutput2[0]) );
  DFF_X1 \StateReg2_s_current_state_reg[61]  ( .D(AddRoundKeyOutput2[61]), 
        .CK(clk), .Q(PermutationOutput2[1]) );
  DFF_X1 \StateReg2_s_current_state_reg[62]  ( .D(AddRoundKeyOutput2[62]), 
        .CK(clk), .Q(PermutationOutput2[2]) );
  DFF_X1 \StateReg2_s_current_state_reg[63]  ( .D(AddRoundKeyOutput2[63]), 
        .CK(clk), .Q(PermutationOutput2[3]) );
  NOR2_X1 \SubCellInst2_LFInst_0_LFInst_0_U8  ( .A1(
        \SubCellInst2_LFInst_0_LFInst_0_n11 ), .A2(
        \SubCellInst2_LFInst_0_LFInst_0_n10 ), .ZN(MCOutput3[0]) );
  AND2_X1 \SubCellInst2_LFInst_0_LFInst_0_U7  ( .A1(PermutationOutput2[3]), 
        .A2(PermutationOutput2[2]), .ZN(\SubCellInst2_LFInst_0_LFInst_0_n10 )
         );
  NOR2_X1 \SubCellInst2_LFInst_0_LFInst_0_U6  ( .A1(PermutationOutput2[1]), 
        .A2(\SubCellInst2_LFInst_0_LFInst_0_n9 ), .ZN(
        \SubCellInst2_LFInst_0_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst2_LFInst_0_LFInst_0_U5  ( .A1(
        \SubCellInst2_LFInst_0_LFInst_0_n8 ), .A2(
        \SubCellInst2_LFInst_0_LFInst_0_n7 ), .ZN(
        \SubCellInst2_LFInst_0_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst2_LFInst_0_LFInst_0_U4  ( .A1(PermutationOutput2[3]), 
        .A2(PermutationOutput2[2]), .ZN(\SubCellInst2_LFInst_0_LFInst_0_n7 )
         );
  INV_X1 \SubCellInst2_LFInst_0_LFInst_0_U3  ( .A(PermutationOutput2[0]), .ZN(
        \SubCellInst2_LFInst_0_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst2_LFInst_0_LFInst_1_U6  ( .A1(
        \SubCellInst2_LFInst_0_LFInst_1_n6 ), .A2(
        \SubCellInst2_LFInst_0_LFInst_1_n5 ), .ZN(MCOutput3[1]) );
  NAND2_X1 \SubCellInst2_LFInst_0_LFInst_1_U5  ( .A1(PermutationOutput2[2]), 
        .A2(PermutationOutput2[0]), .ZN(\SubCellInst2_LFInst_0_LFInst_1_n5 )
         );
  OR2_X1 \SubCellInst2_LFInst_0_LFInst_1_U4  ( .A1(PermutationOutput2[3]), 
        .A2(\SubCellInst2_LFInst_0_LFInst_1_n4 ), .ZN(
        \SubCellInst2_LFInst_0_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst2_LFInst_0_LFInst_1_U3  ( .A1(PermutationOutput2[2]), 
        .A2(PermutationOutput2[0]), .ZN(\SubCellInst2_LFInst_0_LFInst_1_n4 )
         );
  NAND2_X1 \SubCellInst2_LFInst_0_LFInst_2_U8  ( .A1(
        \SubCellInst2_LFInst_0_LFInst_2_n11 ), .A2(
        \SubCellInst2_LFInst_0_LFInst_2_n10 ), .ZN(MCOutput3[2]) );
  OR2_X1 \SubCellInst2_LFInst_0_LFInst_2_U7  ( .A1(PermutationOutput2[0]), 
        .A2(PermutationOutput2[3]), .ZN(\SubCellInst2_LFInst_0_LFInst_2_n10 )
         );
  NAND2_X1 \SubCellInst2_LFInst_0_LFInst_2_U6  ( .A1(PermutationOutput2[1]), 
        .A2(\SubCellInst2_LFInst_0_LFInst_2_n9 ), .ZN(
        \SubCellInst2_LFInst_0_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst2_LFInst_0_LFInst_2_U5  ( .A1(
        \SubCellInst2_LFInst_0_LFInst_2_n8 ), .A2(
        \SubCellInst2_LFInst_0_LFInst_2_n7 ), .ZN(
        \SubCellInst2_LFInst_0_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst2_LFInst_0_LFInst_2_U4  ( .A1(PermutationOutput2[0]), 
        .A2(PermutationOutput2[3]), .ZN(\SubCellInst2_LFInst_0_LFInst_2_n7 )
         );
  INV_X1 \SubCellInst2_LFInst_0_LFInst_2_U3  ( .A(PermutationOutput2[2]), .ZN(
        \SubCellInst2_LFInst_0_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst2_LFInst_0_LFInst_3_U6  ( .A1(
        \SubCellInst2_LFInst_0_LFInst_3_n6 ), .A2(
        \SubCellInst2_LFInst_0_LFInst_3_n5 ), .ZN(MCOutput3[3]) );
  NOR2_X1 \SubCellInst2_LFInst_0_LFInst_3_U5  ( .A1(PermutationOutput2[3]), 
        .A2(PermutationOutput2[0]), .ZN(\SubCellInst2_LFInst_0_LFInst_3_n5 )
         );
  NOR2_X1 \SubCellInst2_LFInst_0_LFInst_3_U4  ( .A1(PermutationOutput2[1]), 
        .A2(\SubCellInst2_LFInst_0_LFInst_3_n4 ), .ZN(
        \SubCellInst2_LFInst_0_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst2_LFInst_0_LFInst_3_U3  ( .A1(PermutationOutput2[3]), 
        .A2(PermutationOutput2[2]), .ZN(\SubCellInst2_LFInst_0_LFInst_3_n4 )
         );
  NOR2_X1 \SubCellInst2_LFInst_1_LFInst_0_U8  ( .A1(
        \SubCellInst2_LFInst_1_LFInst_0_n11 ), .A2(
        \SubCellInst2_LFInst_1_LFInst_0_n10 ), .ZN(MCOutput3[4]) );
  AND2_X1 \SubCellInst2_LFInst_1_LFInst_0_U7  ( .A1(PermutationOutput2[7]), 
        .A2(PermutationOutput2[6]), .ZN(\SubCellInst2_LFInst_1_LFInst_0_n10 )
         );
  NOR2_X1 \SubCellInst2_LFInst_1_LFInst_0_U6  ( .A1(PermutationOutput2[5]), 
        .A2(\SubCellInst2_LFInst_1_LFInst_0_n9 ), .ZN(
        \SubCellInst2_LFInst_1_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst2_LFInst_1_LFInst_0_U5  ( .A1(
        \SubCellInst2_LFInst_1_LFInst_0_n8 ), .A2(
        \SubCellInst2_LFInst_1_LFInst_0_n7 ), .ZN(
        \SubCellInst2_LFInst_1_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst2_LFInst_1_LFInst_0_U4  ( .A1(PermutationOutput2[7]), 
        .A2(PermutationOutput2[6]), .ZN(\SubCellInst2_LFInst_1_LFInst_0_n7 )
         );
  INV_X1 \SubCellInst2_LFInst_1_LFInst_0_U3  ( .A(PermutationOutput2[4]), .ZN(
        \SubCellInst2_LFInst_1_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst2_LFInst_1_LFInst_1_U6  ( .A1(
        \SubCellInst2_LFInst_1_LFInst_1_n6 ), .A2(
        \SubCellInst2_LFInst_1_LFInst_1_n5 ), .ZN(MCOutput3[5]) );
  NAND2_X1 \SubCellInst2_LFInst_1_LFInst_1_U5  ( .A1(PermutationOutput2[6]), 
        .A2(PermutationOutput2[4]), .ZN(\SubCellInst2_LFInst_1_LFInst_1_n5 )
         );
  OR2_X1 \SubCellInst2_LFInst_1_LFInst_1_U4  ( .A1(PermutationOutput2[7]), 
        .A2(\SubCellInst2_LFInst_1_LFInst_1_n4 ), .ZN(
        \SubCellInst2_LFInst_1_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst2_LFInst_1_LFInst_1_U3  ( .A1(PermutationOutput2[6]), 
        .A2(PermutationOutput2[4]), .ZN(\SubCellInst2_LFInst_1_LFInst_1_n4 )
         );
  NAND2_X1 \SubCellInst2_LFInst_1_LFInst_2_U8  ( .A1(
        \SubCellInst2_LFInst_1_LFInst_2_n11 ), .A2(
        \SubCellInst2_LFInst_1_LFInst_2_n10 ), .ZN(MCOutput3[6]) );
  OR2_X1 \SubCellInst2_LFInst_1_LFInst_2_U7  ( .A1(PermutationOutput2[4]), 
        .A2(PermutationOutput2[7]), .ZN(\SubCellInst2_LFInst_1_LFInst_2_n10 )
         );
  NAND2_X1 \SubCellInst2_LFInst_1_LFInst_2_U6  ( .A1(PermutationOutput2[5]), 
        .A2(\SubCellInst2_LFInst_1_LFInst_2_n9 ), .ZN(
        \SubCellInst2_LFInst_1_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst2_LFInst_1_LFInst_2_U5  ( .A1(
        \SubCellInst2_LFInst_1_LFInst_2_n8 ), .A2(
        \SubCellInst2_LFInst_1_LFInst_2_n7 ), .ZN(
        \SubCellInst2_LFInst_1_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst2_LFInst_1_LFInst_2_U4  ( .A1(PermutationOutput2[4]), 
        .A2(PermutationOutput2[7]), .ZN(\SubCellInst2_LFInst_1_LFInst_2_n7 )
         );
  INV_X1 \SubCellInst2_LFInst_1_LFInst_2_U3  ( .A(PermutationOutput2[6]), .ZN(
        \SubCellInst2_LFInst_1_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst2_LFInst_1_LFInst_3_U6  ( .A1(
        \SubCellInst2_LFInst_1_LFInst_3_n6 ), .A2(
        \SubCellInst2_LFInst_1_LFInst_3_n5 ), .ZN(MCOutput3[7]) );
  NOR2_X1 \SubCellInst2_LFInst_1_LFInst_3_U5  ( .A1(PermutationOutput2[7]), 
        .A2(PermutationOutput2[4]), .ZN(\SubCellInst2_LFInst_1_LFInst_3_n5 )
         );
  NOR2_X1 \SubCellInst2_LFInst_1_LFInst_3_U4  ( .A1(PermutationOutput2[5]), 
        .A2(\SubCellInst2_LFInst_1_LFInst_3_n4 ), .ZN(
        \SubCellInst2_LFInst_1_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst2_LFInst_1_LFInst_3_U3  ( .A1(PermutationOutput2[7]), 
        .A2(PermutationOutput2[6]), .ZN(\SubCellInst2_LFInst_1_LFInst_3_n4 )
         );
  NOR2_X1 \SubCellInst2_LFInst_2_LFInst_0_U8  ( .A1(
        \SubCellInst2_LFInst_2_LFInst_0_n11 ), .A2(
        \SubCellInst2_LFInst_2_LFInst_0_n10 ), .ZN(MCOutput3[8]) );
  AND2_X1 \SubCellInst2_LFInst_2_LFInst_0_U7  ( .A1(PermutationOutput2[11]), 
        .A2(PermutationOutput2[10]), .ZN(\SubCellInst2_LFInst_2_LFInst_0_n10 )
         );
  NOR2_X1 \SubCellInst2_LFInst_2_LFInst_0_U6  ( .A1(PermutationOutput2[9]), 
        .A2(\SubCellInst2_LFInst_2_LFInst_0_n9 ), .ZN(
        \SubCellInst2_LFInst_2_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst2_LFInst_2_LFInst_0_U5  ( .A1(
        \SubCellInst2_LFInst_2_LFInst_0_n8 ), .A2(
        \SubCellInst2_LFInst_2_LFInst_0_n7 ), .ZN(
        \SubCellInst2_LFInst_2_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst2_LFInst_2_LFInst_0_U4  ( .A1(PermutationOutput2[11]), 
        .A2(PermutationOutput2[10]), .ZN(\SubCellInst2_LFInst_2_LFInst_0_n7 )
         );
  INV_X1 \SubCellInst2_LFInst_2_LFInst_0_U3  ( .A(PermutationOutput2[8]), .ZN(
        \SubCellInst2_LFInst_2_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst2_LFInst_2_LFInst_1_U6  ( .A1(
        \SubCellInst2_LFInst_2_LFInst_1_n6 ), .A2(
        \SubCellInst2_LFInst_2_LFInst_1_n5 ), .ZN(MCOutput3[9]) );
  NAND2_X1 \SubCellInst2_LFInst_2_LFInst_1_U5  ( .A1(PermutationOutput2[10]), 
        .A2(PermutationOutput2[8]), .ZN(\SubCellInst2_LFInst_2_LFInst_1_n5 )
         );
  OR2_X1 \SubCellInst2_LFInst_2_LFInst_1_U4  ( .A1(PermutationOutput2[11]), 
        .A2(\SubCellInst2_LFInst_2_LFInst_1_n4 ), .ZN(
        \SubCellInst2_LFInst_2_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst2_LFInst_2_LFInst_1_U3  ( .A1(PermutationOutput2[10]), 
        .A2(PermutationOutput2[8]), .ZN(\SubCellInst2_LFInst_2_LFInst_1_n4 )
         );
  NAND2_X1 \SubCellInst2_LFInst_2_LFInst_2_U8  ( .A1(
        \SubCellInst2_LFInst_2_LFInst_2_n11 ), .A2(
        \SubCellInst2_LFInst_2_LFInst_2_n10 ), .ZN(MCOutput3[10]) );
  OR2_X1 \SubCellInst2_LFInst_2_LFInst_2_U7  ( .A1(PermutationOutput2[8]), 
        .A2(PermutationOutput2[11]), .ZN(\SubCellInst2_LFInst_2_LFInst_2_n10 )
         );
  NAND2_X1 \SubCellInst2_LFInst_2_LFInst_2_U6  ( .A1(PermutationOutput2[9]), 
        .A2(\SubCellInst2_LFInst_2_LFInst_2_n9 ), .ZN(
        \SubCellInst2_LFInst_2_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst2_LFInst_2_LFInst_2_U5  ( .A1(
        \SubCellInst2_LFInst_2_LFInst_2_n8 ), .A2(
        \SubCellInst2_LFInst_2_LFInst_2_n7 ), .ZN(
        \SubCellInst2_LFInst_2_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst2_LFInst_2_LFInst_2_U4  ( .A1(PermutationOutput2[8]), 
        .A2(PermutationOutput2[11]), .ZN(\SubCellInst2_LFInst_2_LFInst_2_n7 )
         );
  INV_X1 \SubCellInst2_LFInst_2_LFInst_2_U3  ( .A(PermutationOutput2[10]), 
        .ZN(\SubCellInst2_LFInst_2_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst2_LFInst_2_LFInst_3_U6  ( .A1(
        \SubCellInst2_LFInst_2_LFInst_3_n6 ), .A2(
        \SubCellInst2_LFInst_2_LFInst_3_n5 ), .ZN(MCOutput3[11]) );
  NOR2_X1 \SubCellInst2_LFInst_2_LFInst_3_U5  ( .A1(PermutationOutput2[11]), 
        .A2(PermutationOutput2[8]), .ZN(\SubCellInst2_LFInst_2_LFInst_3_n5 )
         );
  NOR2_X1 \SubCellInst2_LFInst_2_LFInst_3_U4  ( .A1(PermutationOutput2[9]), 
        .A2(\SubCellInst2_LFInst_2_LFInst_3_n4 ), .ZN(
        \SubCellInst2_LFInst_2_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst2_LFInst_2_LFInst_3_U3  ( .A1(PermutationOutput2[11]), 
        .A2(PermutationOutput2[10]), .ZN(\SubCellInst2_LFInst_2_LFInst_3_n4 )
         );
  NOR2_X1 \SubCellInst2_LFInst_3_LFInst_0_U8  ( .A1(
        \SubCellInst2_LFInst_3_LFInst_0_n11 ), .A2(
        \SubCellInst2_LFInst_3_LFInst_0_n10 ), .ZN(MCOutput3[12]) );
  AND2_X1 \SubCellInst2_LFInst_3_LFInst_0_U7  ( .A1(PermutationOutput2[15]), 
        .A2(PermutationOutput2[14]), .ZN(\SubCellInst2_LFInst_3_LFInst_0_n10 )
         );
  NOR2_X1 \SubCellInst2_LFInst_3_LFInst_0_U6  ( .A1(PermutationOutput2[13]), 
        .A2(\SubCellInst2_LFInst_3_LFInst_0_n9 ), .ZN(
        \SubCellInst2_LFInst_3_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst2_LFInst_3_LFInst_0_U5  ( .A1(
        \SubCellInst2_LFInst_3_LFInst_0_n8 ), .A2(
        \SubCellInst2_LFInst_3_LFInst_0_n7 ), .ZN(
        \SubCellInst2_LFInst_3_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst2_LFInst_3_LFInst_0_U4  ( .A1(PermutationOutput2[15]), 
        .A2(PermutationOutput2[14]), .ZN(\SubCellInst2_LFInst_3_LFInst_0_n7 )
         );
  INV_X1 \SubCellInst2_LFInst_3_LFInst_0_U3  ( .A(PermutationOutput2[12]), 
        .ZN(\SubCellInst2_LFInst_3_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst2_LFInst_3_LFInst_1_U6  ( .A1(
        \SubCellInst2_LFInst_3_LFInst_1_n6 ), .A2(
        \SubCellInst2_LFInst_3_LFInst_1_n5 ), .ZN(MCOutput3[13]) );
  NAND2_X1 \SubCellInst2_LFInst_3_LFInst_1_U5  ( .A1(PermutationOutput2[14]), 
        .A2(PermutationOutput2[12]), .ZN(\SubCellInst2_LFInst_3_LFInst_1_n5 )
         );
  OR2_X1 \SubCellInst2_LFInst_3_LFInst_1_U4  ( .A1(PermutationOutput2[15]), 
        .A2(\SubCellInst2_LFInst_3_LFInst_1_n4 ), .ZN(
        \SubCellInst2_LFInst_3_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst2_LFInst_3_LFInst_1_U3  ( .A1(PermutationOutput2[14]), 
        .A2(PermutationOutput2[12]), .ZN(\SubCellInst2_LFInst_3_LFInst_1_n4 )
         );
  NAND2_X1 \SubCellInst2_LFInst_3_LFInst_2_U8  ( .A1(
        \SubCellInst2_LFInst_3_LFInst_2_n11 ), .A2(
        \SubCellInst2_LFInst_3_LFInst_2_n10 ), .ZN(MCOutput3[14]) );
  OR2_X1 \SubCellInst2_LFInst_3_LFInst_2_U7  ( .A1(PermutationOutput2[12]), 
        .A2(PermutationOutput2[15]), .ZN(\SubCellInst2_LFInst_3_LFInst_2_n10 )
         );
  NAND2_X1 \SubCellInst2_LFInst_3_LFInst_2_U6  ( .A1(PermutationOutput2[13]), 
        .A2(\SubCellInst2_LFInst_3_LFInst_2_n9 ), .ZN(
        \SubCellInst2_LFInst_3_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst2_LFInst_3_LFInst_2_U5  ( .A1(
        \SubCellInst2_LFInst_3_LFInst_2_n8 ), .A2(
        \SubCellInst2_LFInst_3_LFInst_2_n7 ), .ZN(
        \SubCellInst2_LFInst_3_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst2_LFInst_3_LFInst_2_U4  ( .A1(PermutationOutput2[12]), 
        .A2(PermutationOutput2[15]), .ZN(\SubCellInst2_LFInst_3_LFInst_2_n7 )
         );
  INV_X1 \SubCellInst2_LFInst_3_LFInst_2_U3  ( .A(PermutationOutput2[14]), 
        .ZN(\SubCellInst2_LFInst_3_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst2_LFInst_3_LFInst_3_U6  ( .A1(
        \SubCellInst2_LFInst_3_LFInst_3_n6 ), .A2(
        \SubCellInst2_LFInst_3_LFInst_3_n5 ), .ZN(MCOutput3[15]) );
  NOR2_X1 \SubCellInst2_LFInst_3_LFInst_3_U5  ( .A1(PermutationOutput2[15]), 
        .A2(PermutationOutput2[12]), .ZN(\SubCellInst2_LFInst_3_LFInst_3_n5 )
         );
  NOR2_X1 \SubCellInst2_LFInst_3_LFInst_3_U4  ( .A1(PermutationOutput2[13]), 
        .A2(\SubCellInst2_LFInst_3_LFInst_3_n4 ), .ZN(
        \SubCellInst2_LFInst_3_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst2_LFInst_3_LFInst_3_U3  ( .A1(PermutationOutput2[15]), 
        .A2(PermutationOutput2[14]), .ZN(\SubCellInst2_LFInst_3_LFInst_3_n4 )
         );
  NOR2_X1 \SubCellInst2_LFInst_4_LFInst_0_U8  ( .A1(
        \SubCellInst2_LFInst_4_LFInst_0_n11 ), .A2(
        \SubCellInst2_LFInst_4_LFInst_0_n10 ), .ZN(MCOutput3[16]) );
  AND2_X1 \SubCellInst2_LFInst_4_LFInst_0_U7  ( .A1(PermutationOutput2[19]), 
        .A2(PermutationOutput2[18]), .ZN(\SubCellInst2_LFInst_4_LFInst_0_n10 )
         );
  NOR2_X1 \SubCellInst2_LFInst_4_LFInst_0_U6  ( .A1(PermutationOutput2[17]), 
        .A2(\SubCellInst2_LFInst_4_LFInst_0_n9 ), .ZN(
        \SubCellInst2_LFInst_4_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst2_LFInst_4_LFInst_0_U5  ( .A1(
        \SubCellInst2_LFInst_4_LFInst_0_n8 ), .A2(
        \SubCellInst2_LFInst_4_LFInst_0_n7 ), .ZN(
        \SubCellInst2_LFInst_4_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst2_LFInst_4_LFInst_0_U4  ( .A1(PermutationOutput2[19]), 
        .A2(PermutationOutput2[18]), .ZN(\SubCellInst2_LFInst_4_LFInst_0_n7 )
         );
  INV_X1 \SubCellInst2_LFInst_4_LFInst_0_U3  ( .A(PermutationOutput2[16]), 
        .ZN(\SubCellInst2_LFInst_4_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst2_LFInst_4_LFInst_1_U6  ( .A1(
        \SubCellInst2_LFInst_4_LFInst_1_n6 ), .A2(
        \SubCellInst2_LFInst_4_LFInst_1_n5 ), .ZN(MCOutput3[17]) );
  NAND2_X1 \SubCellInst2_LFInst_4_LFInst_1_U5  ( .A1(PermutationOutput2[18]), 
        .A2(PermutationOutput2[16]), .ZN(\SubCellInst2_LFInst_4_LFInst_1_n5 )
         );
  OR2_X1 \SubCellInst2_LFInst_4_LFInst_1_U4  ( .A1(PermutationOutput2[19]), 
        .A2(\SubCellInst2_LFInst_4_LFInst_1_n4 ), .ZN(
        \SubCellInst2_LFInst_4_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst2_LFInst_4_LFInst_1_U3  ( .A1(PermutationOutput2[18]), 
        .A2(PermutationOutput2[16]), .ZN(\SubCellInst2_LFInst_4_LFInst_1_n4 )
         );
  NAND2_X1 \SubCellInst2_LFInst_4_LFInst_2_U8  ( .A1(
        \SubCellInst2_LFInst_4_LFInst_2_n11 ), .A2(
        \SubCellInst2_LFInst_4_LFInst_2_n10 ), .ZN(MCOutput3[18]) );
  OR2_X1 \SubCellInst2_LFInst_4_LFInst_2_U7  ( .A1(PermutationOutput2[16]), 
        .A2(PermutationOutput2[19]), .ZN(\SubCellInst2_LFInst_4_LFInst_2_n10 )
         );
  NAND2_X1 \SubCellInst2_LFInst_4_LFInst_2_U6  ( .A1(PermutationOutput2[17]), 
        .A2(\SubCellInst2_LFInst_4_LFInst_2_n9 ), .ZN(
        \SubCellInst2_LFInst_4_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst2_LFInst_4_LFInst_2_U5  ( .A1(
        \SubCellInst2_LFInst_4_LFInst_2_n8 ), .A2(
        \SubCellInst2_LFInst_4_LFInst_2_n7 ), .ZN(
        \SubCellInst2_LFInst_4_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst2_LFInst_4_LFInst_2_U4  ( .A1(PermutationOutput2[16]), 
        .A2(PermutationOutput2[19]), .ZN(\SubCellInst2_LFInst_4_LFInst_2_n7 )
         );
  INV_X1 \SubCellInst2_LFInst_4_LFInst_2_U3  ( .A(PermutationOutput2[18]), 
        .ZN(\SubCellInst2_LFInst_4_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst2_LFInst_4_LFInst_3_U6  ( .A1(
        \SubCellInst2_LFInst_4_LFInst_3_n6 ), .A2(
        \SubCellInst2_LFInst_4_LFInst_3_n5 ), .ZN(MCOutput3[19]) );
  NOR2_X1 \SubCellInst2_LFInst_4_LFInst_3_U5  ( .A1(PermutationOutput2[19]), 
        .A2(PermutationOutput2[16]), .ZN(\SubCellInst2_LFInst_4_LFInst_3_n5 )
         );
  NOR2_X1 \SubCellInst2_LFInst_4_LFInst_3_U4  ( .A1(PermutationOutput2[17]), 
        .A2(\SubCellInst2_LFInst_4_LFInst_3_n4 ), .ZN(
        \SubCellInst2_LFInst_4_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst2_LFInst_4_LFInst_3_U3  ( .A1(PermutationOutput2[19]), 
        .A2(PermutationOutput2[18]), .ZN(\SubCellInst2_LFInst_4_LFInst_3_n4 )
         );
  NOR2_X1 \SubCellInst2_LFInst_5_LFInst_0_U8  ( .A1(
        \SubCellInst2_LFInst_5_LFInst_0_n11 ), .A2(
        \SubCellInst2_LFInst_5_LFInst_0_n10 ), .ZN(MCOutput3[20]) );
  AND2_X1 \SubCellInst2_LFInst_5_LFInst_0_U7  ( .A1(PermutationOutput2[23]), 
        .A2(PermutationOutput2[22]), .ZN(\SubCellInst2_LFInst_5_LFInst_0_n10 )
         );
  NOR2_X1 \SubCellInst2_LFInst_5_LFInst_0_U6  ( .A1(PermutationOutput2[21]), 
        .A2(\SubCellInst2_LFInst_5_LFInst_0_n9 ), .ZN(
        \SubCellInst2_LFInst_5_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst2_LFInst_5_LFInst_0_U5  ( .A1(
        \SubCellInst2_LFInst_5_LFInst_0_n8 ), .A2(
        \SubCellInst2_LFInst_5_LFInst_0_n7 ), .ZN(
        \SubCellInst2_LFInst_5_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst2_LFInst_5_LFInst_0_U4  ( .A1(PermutationOutput2[23]), 
        .A2(PermutationOutput2[22]), .ZN(\SubCellInst2_LFInst_5_LFInst_0_n7 )
         );
  INV_X1 \SubCellInst2_LFInst_5_LFInst_0_U3  ( .A(PermutationOutput2[20]), 
        .ZN(\SubCellInst2_LFInst_5_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst2_LFInst_5_LFInst_1_U6  ( .A1(
        \SubCellInst2_LFInst_5_LFInst_1_n6 ), .A2(
        \SubCellInst2_LFInst_5_LFInst_1_n5 ), .ZN(MCOutput3[21]) );
  NAND2_X1 \SubCellInst2_LFInst_5_LFInst_1_U5  ( .A1(PermutationOutput2[22]), 
        .A2(PermutationOutput2[20]), .ZN(\SubCellInst2_LFInst_5_LFInst_1_n5 )
         );
  OR2_X1 \SubCellInst2_LFInst_5_LFInst_1_U4  ( .A1(PermutationOutput2[23]), 
        .A2(\SubCellInst2_LFInst_5_LFInst_1_n4 ), .ZN(
        \SubCellInst2_LFInst_5_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst2_LFInst_5_LFInst_1_U3  ( .A1(PermutationOutput2[22]), 
        .A2(PermutationOutput2[20]), .ZN(\SubCellInst2_LFInst_5_LFInst_1_n4 )
         );
  NAND2_X1 \SubCellInst2_LFInst_5_LFInst_2_U8  ( .A1(
        \SubCellInst2_LFInst_5_LFInst_2_n11 ), .A2(
        \SubCellInst2_LFInst_5_LFInst_2_n10 ), .ZN(MCOutput3[22]) );
  OR2_X1 \SubCellInst2_LFInst_5_LFInst_2_U7  ( .A1(PermutationOutput2[20]), 
        .A2(PermutationOutput2[23]), .ZN(\SubCellInst2_LFInst_5_LFInst_2_n10 )
         );
  NAND2_X1 \SubCellInst2_LFInst_5_LFInst_2_U6  ( .A1(PermutationOutput2[21]), 
        .A2(\SubCellInst2_LFInst_5_LFInst_2_n9 ), .ZN(
        \SubCellInst2_LFInst_5_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst2_LFInst_5_LFInst_2_U5  ( .A1(
        \SubCellInst2_LFInst_5_LFInst_2_n8 ), .A2(
        \SubCellInst2_LFInst_5_LFInst_2_n7 ), .ZN(
        \SubCellInst2_LFInst_5_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst2_LFInst_5_LFInst_2_U4  ( .A1(PermutationOutput2[20]), 
        .A2(PermutationOutput2[23]), .ZN(\SubCellInst2_LFInst_5_LFInst_2_n7 )
         );
  INV_X1 \SubCellInst2_LFInst_5_LFInst_2_U3  ( .A(PermutationOutput2[22]), 
        .ZN(\SubCellInst2_LFInst_5_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst2_LFInst_5_LFInst_3_U6  ( .A1(
        \SubCellInst2_LFInst_5_LFInst_3_n6 ), .A2(
        \SubCellInst2_LFInst_5_LFInst_3_n5 ), .ZN(MCOutput3[23]) );
  NOR2_X1 \SubCellInst2_LFInst_5_LFInst_3_U5  ( .A1(PermutationOutput2[23]), 
        .A2(PermutationOutput2[20]), .ZN(\SubCellInst2_LFInst_5_LFInst_3_n5 )
         );
  NOR2_X1 \SubCellInst2_LFInst_5_LFInst_3_U4  ( .A1(PermutationOutput2[21]), 
        .A2(\SubCellInst2_LFInst_5_LFInst_3_n4 ), .ZN(
        \SubCellInst2_LFInst_5_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst2_LFInst_5_LFInst_3_U3  ( .A1(PermutationOutput2[23]), 
        .A2(PermutationOutput2[22]), .ZN(\SubCellInst2_LFInst_5_LFInst_3_n4 )
         );
  NOR2_X1 \SubCellInst2_LFInst_6_LFInst_0_U8  ( .A1(
        \SubCellInst2_LFInst_6_LFInst_0_n11 ), .A2(
        \SubCellInst2_LFInst_6_LFInst_0_n10 ), .ZN(MCOutput3[24]) );
  AND2_X1 \SubCellInst2_LFInst_6_LFInst_0_U7  ( .A1(PermutationOutput2[27]), 
        .A2(PermutationOutput2[26]), .ZN(\SubCellInst2_LFInst_6_LFInst_0_n10 )
         );
  NOR2_X1 \SubCellInst2_LFInst_6_LFInst_0_U6  ( .A1(PermutationOutput2[25]), 
        .A2(\SubCellInst2_LFInst_6_LFInst_0_n9 ), .ZN(
        \SubCellInst2_LFInst_6_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst2_LFInst_6_LFInst_0_U5  ( .A1(
        \SubCellInst2_LFInst_6_LFInst_0_n8 ), .A2(
        \SubCellInst2_LFInst_6_LFInst_0_n7 ), .ZN(
        \SubCellInst2_LFInst_6_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst2_LFInst_6_LFInst_0_U4  ( .A1(PermutationOutput2[27]), 
        .A2(PermutationOutput2[26]), .ZN(\SubCellInst2_LFInst_6_LFInst_0_n7 )
         );
  INV_X1 \SubCellInst2_LFInst_6_LFInst_0_U3  ( .A(PermutationOutput2[24]), 
        .ZN(\SubCellInst2_LFInst_6_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst2_LFInst_6_LFInst_1_U6  ( .A1(
        \SubCellInst2_LFInst_6_LFInst_1_n6 ), .A2(
        \SubCellInst2_LFInst_6_LFInst_1_n5 ), .ZN(MCOutput3[25]) );
  NAND2_X1 \SubCellInst2_LFInst_6_LFInst_1_U5  ( .A1(PermutationOutput2[26]), 
        .A2(PermutationOutput2[24]), .ZN(\SubCellInst2_LFInst_6_LFInst_1_n5 )
         );
  OR2_X1 \SubCellInst2_LFInst_6_LFInst_1_U4  ( .A1(PermutationOutput2[27]), 
        .A2(\SubCellInst2_LFInst_6_LFInst_1_n4 ), .ZN(
        \SubCellInst2_LFInst_6_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst2_LFInst_6_LFInst_1_U3  ( .A1(PermutationOutput2[26]), 
        .A2(PermutationOutput2[24]), .ZN(\SubCellInst2_LFInst_6_LFInst_1_n4 )
         );
  NAND2_X1 \SubCellInst2_LFInst_6_LFInst_2_U8  ( .A1(
        \SubCellInst2_LFInst_6_LFInst_2_n11 ), .A2(
        \SubCellInst2_LFInst_6_LFInst_2_n10 ), .ZN(MCOutput3[26]) );
  OR2_X1 \SubCellInst2_LFInst_6_LFInst_2_U7  ( .A1(PermutationOutput2[24]), 
        .A2(PermutationOutput2[27]), .ZN(\SubCellInst2_LFInst_6_LFInst_2_n10 )
         );
  NAND2_X1 \SubCellInst2_LFInst_6_LFInst_2_U6  ( .A1(PermutationOutput2[25]), 
        .A2(\SubCellInst2_LFInst_6_LFInst_2_n9 ), .ZN(
        \SubCellInst2_LFInst_6_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst2_LFInst_6_LFInst_2_U5  ( .A1(
        \SubCellInst2_LFInst_6_LFInst_2_n8 ), .A2(
        \SubCellInst2_LFInst_6_LFInst_2_n7 ), .ZN(
        \SubCellInst2_LFInst_6_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst2_LFInst_6_LFInst_2_U4  ( .A1(PermutationOutput2[24]), 
        .A2(PermutationOutput2[27]), .ZN(\SubCellInst2_LFInst_6_LFInst_2_n7 )
         );
  INV_X1 \SubCellInst2_LFInst_6_LFInst_2_U3  ( .A(PermutationOutput2[26]), 
        .ZN(\SubCellInst2_LFInst_6_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst2_LFInst_6_LFInst_3_U6  ( .A1(
        \SubCellInst2_LFInst_6_LFInst_3_n6 ), .A2(
        \SubCellInst2_LFInst_6_LFInst_3_n5 ), .ZN(MCOutput3[27]) );
  NOR2_X1 \SubCellInst2_LFInst_6_LFInst_3_U5  ( .A1(PermutationOutput2[27]), 
        .A2(PermutationOutput2[24]), .ZN(\SubCellInst2_LFInst_6_LFInst_3_n5 )
         );
  NOR2_X1 \SubCellInst2_LFInst_6_LFInst_3_U4  ( .A1(PermutationOutput2[25]), 
        .A2(\SubCellInst2_LFInst_6_LFInst_3_n4 ), .ZN(
        \SubCellInst2_LFInst_6_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst2_LFInst_6_LFInst_3_U3  ( .A1(PermutationOutput2[27]), 
        .A2(PermutationOutput2[26]), .ZN(\SubCellInst2_LFInst_6_LFInst_3_n4 )
         );
  NOR2_X1 \SubCellInst2_LFInst_7_LFInst_0_U8  ( .A1(
        \SubCellInst2_LFInst_7_LFInst_0_n11 ), .A2(
        \SubCellInst2_LFInst_7_LFInst_0_n10 ), .ZN(MCOutput3[28]) );
  AND2_X1 \SubCellInst2_LFInst_7_LFInst_0_U7  ( .A1(PermutationOutput2[31]), 
        .A2(PermutationOutput2[30]), .ZN(\SubCellInst2_LFInst_7_LFInst_0_n10 )
         );
  NOR2_X1 \SubCellInst2_LFInst_7_LFInst_0_U6  ( .A1(PermutationOutput2[29]), 
        .A2(\SubCellInst2_LFInst_7_LFInst_0_n9 ), .ZN(
        \SubCellInst2_LFInst_7_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst2_LFInst_7_LFInst_0_U5  ( .A1(
        \SubCellInst2_LFInst_7_LFInst_0_n8 ), .A2(
        \SubCellInst2_LFInst_7_LFInst_0_n7 ), .ZN(
        \SubCellInst2_LFInst_7_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst2_LFInst_7_LFInst_0_U4  ( .A1(PermutationOutput2[31]), 
        .A2(PermutationOutput2[30]), .ZN(\SubCellInst2_LFInst_7_LFInst_0_n7 )
         );
  INV_X1 \SubCellInst2_LFInst_7_LFInst_0_U3  ( .A(PermutationOutput2[28]), 
        .ZN(\SubCellInst2_LFInst_7_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst2_LFInst_7_LFInst_1_U6  ( .A1(
        \SubCellInst2_LFInst_7_LFInst_1_n6 ), .A2(
        \SubCellInst2_LFInst_7_LFInst_1_n5 ), .ZN(MCOutput3[29]) );
  NAND2_X1 \SubCellInst2_LFInst_7_LFInst_1_U5  ( .A1(PermutationOutput2[30]), 
        .A2(PermutationOutput2[28]), .ZN(\SubCellInst2_LFInst_7_LFInst_1_n5 )
         );
  OR2_X1 \SubCellInst2_LFInst_7_LFInst_1_U4  ( .A1(PermutationOutput2[31]), 
        .A2(\SubCellInst2_LFInst_7_LFInst_1_n4 ), .ZN(
        \SubCellInst2_LFInst_7_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst2_LFInst_7_LFInst_1_U3  ( .A1(PermutationOutput2[30]), 
        .A2(PermutationOutput2[28]), .ZN(\SubCellInst2_LFInst_7_LFInst_1_n4 )
         );
  NAND2_X1 \SubCellInst2_LFInst_7_LFInst_2_U8  ( .A1(
        \SubCellInst2_LFInst_7_LFInst_2_n11 ), .A2(
        \SubCellInst2_LFInst_7_LFInst_2_n10 ), .ZN(MCOutput3[30]) );
  OR2_X1 \SubCellInst2_LFInst_7_LFInst_2_U7  ( .A1(PermutationOutput2[28]), 
        .A2(PermutationOutput2[31]), .ZN(\SubCellInst2_LFInst_7_LFInst_2_n10 )
         );
  NAND2_X1 \SubCellInst2_LFInst_7_LFInst_2_U6  ( .A1(PermutationOutput2[29]), 
        .A2(\SubCellInst2_LFInst_7_LFInst_2_n9 ), .ZN(
        \SubCellInst2_LFInst_7_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst2_LFInst_7_LFInst_2_U5  ( .A1(
        \SubCellInst2_LFInst_7_LFInst_2_n8 ), .A2(
        \SubCellInst2_LFInst_7_LFInst_2_n7 ), .ZN(
        \SubCellInst2_LFInst_7_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst2_LFInst_7_LFInst_2_U4  ( .A1(PermutationOutput2[28]), 
        .A2(PermutationOutput2[31]), .ZN(\SubCellInst2_LFInst_7_LFInst_2_n7 )
         );
  INV_X1 \SubCellInst2_LFInst_7_LFInst_2_U3  ( .A(PermutationOutput2[30]), 
        .ZN(\SubCellInst2_LFInst_7_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst2_LFInst_7_LFInst_3_U6  ( .A1(
        \SubCellInst2_LFInst_7_LFInst_3_n6 ), .A2(
        \SubCellInst2_LFInst_7_LFInst_3_n5 ), .ZN(MCOutput3[31]) );
  NOR2_X1 \SubCellInst2_LFInst_7_LFInst_3_U5  ( .A1(PermutationOutput2[31]), 
        .A2(PermutationOutput2[28]), .ZN(\SubCellInst2_LFInst_7_LFInst_3_n5 )
         );
  NOR2_X1 \SubCellInst2_LFInst_7_LFInst_3_U4  ( .A1(PermutationOutput2[29]), 
        .A2(\SubCellInst2_LFInst_7_LFInst_3_n4 ), .ZN(
        \SubCellInst2_LFInst_7_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst2_LFInst_7_LFInst_3_U3  ( .A1(PermutationOutput2[31]), 
        .A2(PermutationOutput2[30]), .ZN(\SubCellInst2_LFInst_7_LFInst_3_n4 )
         );
  NOR2_X1 \SubCellInst2_LFInst_8_LFInst_0_U8  ( .A1(
        \SubCellInst2_LFInst_8_LFInst_0_n11 ), .A2(
        \SubCellInst2_LFInst_8_LFInst_0_n10 ), .ZN(Feedback2[32]) );
  AND2_X1 \SubCellInst2_LFInst_8_LFInst_0_U7  ( .A1(PermutationOutput2[35]), 
        .A2(PermutationOutput2[34]), .ZN(\SubCellInst2_LFInst_8_LFInst_0_n10 )
         );
  NOR2_X1 \SubCellInst2_LFInst_8_LFInst_0_U6  ( .A1(PermutationOutput2[33]), 
        .A2(\SubCellInst2_LFInst_8_LFInst_0_n9 ), .ZN(
        \SubCellInst2_LFInst_8_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst2_LFInst_8_LFInst_0_U5  ( .A1(
        \SubCellInst2_LFInst_8_LFInst_0_n8 ), .A2(
        \SubCellInst2_LFInst_8_LFInst_0_n7 ), .ZN(
        \SubCellInst2_LFInst_8_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst2_LFInst_8_LFInst_0_U4  ( .A1(PermutationOutput2[35]), 
        .A2(PermutationOutput2[34]), .ZN(\SubCellInst2_LFInst_8_LFInst_0_n7 )
         );
  INV_X1 \SubCellInst2_LFInst_8_LFInst_0_U3  ( .A(PermutationOutput2[32]), 
        .ZN(\SubCellInst2_LFInst_8_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst2_LFInst_8_LFInst_1_U6  ( .A1(
        \SubCellInst2_LFInst_8_LFInst_1_n6 ), .A2(
        \SubCellInst2_LFInst_8_LFInst_1_n5 ), .ZN(Feedback2[33]) );
  NAND2_X1 \SubCellInst2_LFInst_8_LFInst_1_U5  ( .A1(PermutationOutput2[34]), 
        .A2(PermutationOutput2[32]), .ZN(\SubCellInst2_LFInst_8_LFInst_1_n5 )
         );
  OR2_X1 \SubCellInst2_LFInst_8_LFInst_1_U4  ( .A1(PermutationOutput2[35]), 
        .A2(\SubCellInst2_LFInst_8_LFInst_1_n4 ), .ZN(
        \SubCellInst2_LFInst_8_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst2_LFInst_8_LFInst_1_U3  ( .A1(PermutationOutput2[34]), 
        .A2(PermutationOutput2[32]), .ZN(\SubCellInst2_LFInst_8_LFInst_1_n4 )
         );
  NAND2_X1 \SubCellInst2_LFInst_8_LFInst_2_U8  ( .A1(
        \SubCellInst2_LFInst_8_LFInst_2_n11 ), .A2(
        \SubCellInst2_LFInst_8_LFInst_2_n10 ), .ZN(Feedback2[34]) );
  OR2_X1 \SubCellInst2_LFInst_8_LFInst_2_U7  ( .A1(PermutationOutput2[32]), 
        .A2(PermutationOutput2[35]), .ZN(\SubCellInst2_LFInst_8_LFInst_2_n10 )
         );
  NAND2_X1 \SubCellInst2_LFInst_8_LFInst_2_U6  ( .A1(PermutationOutput2[33]), 
        .A2(\SubCellInst2_LFInst_8_LFInst_2_n9 ), .ZN(
        \SubCellInst2_LFInst_8_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst2_LFInst_8_LFInst_2_U5  ( .A1(
        \SubCellInst2_LFInst_8_LFInst_2_n8 ), .A2(
        \SubCellInst2_LFInst_8_LFInst_2_n7 ), .ZN(
        \SubCellInst2_LFInst_8_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst2_LFInst_8_LFInst_2_U4  ( .A1(PermutationOutput2[32]), 
        .A2(PermutationOutput2[35]), .ZN(\SubCellInst2_LFInst_8_LFInst_2_n7 )
         );
  INV_X1 \SubCellInst2_LFInst_8_LFInst_2_U3  ( .A(PermutationOutput2[34]), 
        .ZN(\SubCellInst2_LFInst_8_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst2_LFInst_8_LFInst_3_U6  ( .A1(
        \SubCellInst2_LFInst_8_LFInst_3_n6 ), .A2(
        \SubCellInst2_LFInst_8_LFInst_3_n5 ), .ZN(Feedback2[35]) );
  NOR2_X1 \SubCellInst2_LFInst_8_LFInst_3_U5  ( .A1(PermutationOutput2[35]), 
        .A2(PermutationOutput2[32]), .ZN(\SubCellInst2_LFInst_8_LFInst_3_n5 )
         );
  NOR2_X1 \SubCellInst2_LFInst_8_LFInst_3_U4  ( .A1(PermutationOutput2[33]), 
        .A2(\SubCellInst2_LFInst_8_LFInst_3_n4 ), .ZN(
        \SubCellInst2_LFInst_8_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst2_LFInst_8_LFInst_3_U3  ( .A1(PermutationOutput2[35]), 
        .A2(PermutationOutput2[34]), .ZN(\SubCellInst2_LFInst_8_LFInst_3_n4 )
         );
  NOR2_X1 \SubCellInst2_LFInst_9_LFInst_0_U8  ( .A1(
        \SubCellInst2_LFInst_9_LFInst_0_n11 ), .A2(
        \SubCellInst2_LFInst_9_LFInst_0_n10 ), .ZN(Feedback2[36]) );
  AND2_X1 \SubCellInst2_LFInst_9_LFInst_0_U7  ( .A1(PermutationOutput2[39]), 
        .A2(PermutationOutput2[38]), .ZN(\SubCellInst2_LFInst_9_LFInst_0_n10 )
         );
  NOR2_X1 \SubCellInst2_LFInst_9_LFInst_0_U6  ( .A1(PermutationOutput2[37]), 
        .A2(\SubCellInst2_LFInst_9_LFInst_0_n9 ), .ZN(
        \SubCellInst2_LFInst_9_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst2_LFInst_9_LFInst_0_U5  ( .A1(
        \SubCellInst2_LFInst_9_LFInst_0_n8 ), .A2(
        \SubCellInst2_LFInst_9_LFInst_0_n7 ), .ZN(
        \SubCellInst2_LFInst_9_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst2_LFInst_9_LFInst_0_U4  ( .A1(PermutationOutput2[39]), 
        .A2(PermutationOutput2[38]), .ZN(\SubCellInst2_LFInst_9_LFInst_0_n7 )
         );
  INV_X1 \SubCellInst2_LFInst_9_LFInst_0_U3  ( .A(PermutationOutput2[36]), 
        .ZN(\SubCellInst2_LFInst_9_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst2_LFInst_9_LFInst_1_U6  ( .A1(
        \SubCellInst2_LFInst_9_LFInst_1_n6 ), .A2(
        \SubCellInst2_LFInst_9_LFInst_1_n5 ), .ZN(Feedback2[37]) );
  NAND2_X1 \SubCellInst2_LFInst_9_LFInst_1_U5  ( .A1(PermutationOutput2[38]), 
        .A2(PermutationOutput2[36]), .ZN(\SubCellInst2_LFInst_9_LFInst_1_n5 )
         );
  OR2_X1 \SubCellInst2_LFInst_9_LFInst_1_U4  ( .A1(PermutationOutput2[39]), 
        .A2(\SubCellInst2_LFInst_9_LFInst_1_n4 ), .ZN(
        \SubCellInst2_LFInst_9_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst2_LFInst_9_LFInst_1_U3  ( .A1(PermutationOutput2[38]), 
        .A2(PermutationOutput2[36]), .ZN(\SubCellInst2_LFInst_9_LFInst_1_n4 )
         );
  NAND2_X1 \SubCellInst2_LFInst_9_LFInst_2_U8  ( .A1(
        \SubCellInst2_LFInst_9_LFInst_2_n11 ), .A2(
        \SubCellInst2_LFInst_9_LFInst_2_n10 ), .ZN(Feedback2[38]) );
  OR2_X1 \SubCellInst2_LFInst_9_LFInst_2_U7  ( .A1(PermutationOutput2[36]), 
        .A2(PermutationOutput2[39]), .ZN(\SubCellInst2_LFInst_9_LFInst_2_n10 )
         );
  NAND2_X1 \SubCellInst2_LFInst_9_LFInst_2_U6  ( .A1(PermutationOutput2[37]), 
        .A2(\SubCellInst2_LFInst_9_LFInst_2_n9 ), .ZN(
        \SubCellInst2_LFInst_9_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst2_LFInst_9_LFInst_2_U5  ( .A1(
        \SubCellInst2_LFInst_9_LFInst_2_n8 ), .A2(
        \SubCellInst2_LFInst_9_LFInst_2_n7 ), .ZN(
        \SubCellInst2_LFInst_9_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst2_LFInst_9_LFInst_2_U4  ( .A1(PermutationOutput2[36]), 
        .A2(PermutationOutput2[39]), .ZN(\SubCellInst2_LFInst_9_LFInst_2_n7 )
         );
  INV_X1 \SubCellInst2_LFInst_9_LFInst_2_U3  ( .A(PermutationOutput2[38]), 
        .ZN(\SubCellInst2_LFInst_9_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst2_LFInst_9_LFInst_3_U6  ( .A1(
        \SubCellInst2_LFInst_9_LFInst_3_n6 ), .A2(
        \SubCellInst2_LFInst_9_LFInst_3_n5 ), .ZN(Feedback2[39]) );
  NOR2_X1 \SubCellInst2_LFInst_9_LFInst_3_U5  ( .A1(PermutationOutput2[39]), 
        .A2(PermutationOutput2[36]), .ZN(\SubCellInst2_LFInst_9_LFInst_3_n5 )
         );
  NOR2_X1 \SubCellInst2_LFInst_9_LFInst_3_U4  ( .A1(PermutationOutput2[37]), 
        .A2(\SubCellInst2_LFInst_9_LFInst_3_n4 ), .ZN(
        \SubCellInst2_LFInst_9_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst2_LFInst_9_LFInst_3_U3  ( .A1(PermutationOutput2[39]), 
        .A2(PermutationOutput2[38]), .ZN(\SubCellInst2_LFInst_9_LFInst_3_n4 )
         );
  NOR2_X1 \SubCellInst2_LFInst_10_LFInst_0_U8  ( .A1(
        \SubCellInst2_LFInst_10_LFInst_0_n11 ), .A2(
        \SubCellInst2_LFInst_10_LFInst_0_n10 ), .ZN(Feedback2[40]) );
  AND2_X1 \SubCellInst2_LFInst_10_LFInst_0_U7  ( .A1(PermutationOutput2[43]), 
        .A2(PermutationOutput2[42]), .ZN(\SubCellInst2_LFInst_10_LFInst_0_n10 ) );
  NOR2_X1 \SubCellInst2_LFInst_10_LFInst_0_U6  ( .A1(PermutationOutput2[41]), 
        .A2(\SubCellInst2_LFInst_10_LFInst_0_n9 ), .ZN(
        \SubCellInst2_LFInst_10_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst2_LFInst_10_LFInst_0_U5  ( .A1(
        \SubCellInst2_LFInst_10_LFInst_0_n8 ), .A2(
        \SubCellInst2_LFInst_10_LFInst_0_n7 ), .ZN(
        \SubCellInst2_LFInst_10_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst2_LFInst_10_LFInst_0_U4  ( .A1(PermutationOutput2[43]), 
        .A2(PermutationOutput2[42]), .ZN(\SubCellInst2_LFInst_10_LFInst_0_n7 )
         );
  INV_X1 \SubCellInst2_LFInst_10_LFInst_0_U3  ( .A(PermutationOutput2[40]), 
        .ZN(\SubCellInst2_LFInst_10_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst2_LFInst_10_LFInst_1_U6  ( .A1(
        \SubCellInst2_LFInst_10_LFInst_1_n6 ), .A2(
        \SubCellInst2_LFInst_10_LFInst_1_n5 ), .ZN(Feedback2[41]) );
  NAND2_X1 \SubCellInst2_LFInst_10_LFInst_1_U5  ( .A1(PermutationOutput2[42]), 
        .A2(PermutationOutput2[40]), .ZN(\SubCellInst2_LFInst_10_LFInst_1_n5 )
         );
  OR2_X1 \SubCellInst2_LFInst_10_LFInst_1_U4  ( .A1(PermutationOutput2[43]), 
        .A2(\SubCellInst2_LFInst_10_LFInst_1_n4 ), .ZN(
        \SubCellInst2_LFInst_10_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst2_LFInst_10_LFInst_1_U3  ( .A1(PermutationOutput2[42]), 
        .A2(PermutationOutput2[40]), .ZN(\SubCellInst2_LFInst_10_LFInst_1_n4 )
         );
  NAND2_X1 \SubCellInst2_LFInst_10_LFInst_2_U8  ( .A1(
        \SubCellInst2_LFInst_10_LFInst_2_n11 ), .A2(
        \SubCellInst2_LFInst_10_LFInst_2_n10 ), .ZN(Feedback2[42]) );
  OR2_X1 \SubCellInst2_LFInst_10_LFInst_2_U7  ( .A1(PermutationOutput2[40]), 
        .A2(PermutationOutput2[43]), .ZN(\SubCellInst2_LFInst_10_LFInst_2_n10 ) );
  NAND2_X1 \SubCellInst2_LFInst_10_LFInst_2_U6  ( .A1(PermutationOutput2[41]), 
        .A2(\SubCellInst2_LFInst_10_LFInst_2_n9 ), .ZN(
        \SubCellInst2_LFInst_10_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst2_LFInst_10_LFInst_2_U5  ( .A1(
        \SubCellInst2_LFInst_10_LFInst_2_n8 ), .A2(
        \SubCellInst2_LFInst_10_LFInst_2_n7 ), .ZN(
        \SubCellInst2_LFInst_10_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst2_LFInst_10_LFInst_2_U4  ( .A1(PermutationOutput2[40]), 
        .A2(PermutationOutput2[43]), .ZN(\SubCellInst2_LFInst_10_LFInst_2_n7 )
         );
  INV_X1 \SubCellInst2_LFInst_10_LFInst_2_U3  ( .A(PermutationOutput2[42]), 
        .ZN(\SubCellInst2_LFInst_10_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst2_LFInst_10_LFInst_3_U6  ( .A1(
        \SubCellInst2_LFInst_10_LFInst_3_n6 ), .A2(
        \SubCellInst2_LFInst_10_LFInst_3_n5 ), .ZN(Feedback2[43]) );
  NOR2_X1 \SubCellInst2_LFInst_10_LFInst_3_U5  ( .A1(PermutationOutput2[43]), 
        .A2(PermutationOutput2[40]), .ZN(\SubCellInst2_LFInst_10_LFInst_3_n5 )
         );
  NOR2_X1 \SubCellInst2_LFInst_10_LFInst_3_U4  ( .A1(PermutationOutput2[41]), 
        .A2(\SubCellInst2_LFInst_10_LFInst_3_n4 ), .ZN(
        \SubCellInst2_LFInst_10_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst2_LFInst_10_LFInst_3_U3  ( .A1(PermutationOutput2[43]), 
        .A2(PermutationOutput2[42]), .ZN(\SubCellInst2_LFInst_10_LFInst_3_n4 )
         );
  NOR2_X1 \SubCellInst2_LFInst_11_LFInst_0_U8  ( .A1(
        \SubCellInst2_LFInst_11_LFInst_0_n11 ), .A2(
        \SubCellInst2_LFInst_11_LFInst_0_n10 ), .ZN(Feedback2[44]) );
  AND2_X1 \SubCellInst2_LFInst_11_LFInst_0_U7  ( .A1(PermutationOutput2[47]), 
        .A2(PermutationOutput2[46]), .ZN(\SubCellInst2_LFInst_11_LFInst_0_n10 ) );
  NOR2_X1 \SubCellInst2_LFInst_11_LFInst_0_U6  ( .A1(PermutationOutput2[45]), 
        .A2(\SubCellInst2_LFInst_11_LFInst_0_n9 ), .ZN(
        \SubCellInst2_LFInst_11_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst2_LFInst_11_LFInst_0_U5  ( .A1(
        \SubCellInst2_LFInst_11_LFInst_0_n8 ), .A2(
        \SubCellInst2_LFInst_11_LFInst_0_n7 ), .ZN(
        \SubCellInst2_LFInst_11_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst2_LFInst_11_LFInst_0_U4  ( .A1(PermutationOutput2[47]), 
        .A2(PermutationOutput2[46]), .ZN(\SubCellInst2_LFInst_11_LFInst_0_n7 )
         );
  INV_X1 \SubCellInst2_LFInst_11_LFInst_0_U3  ( .A(PermutationOutput2[44]), 
        .ZN(\SubCellInst2_LFInst_11_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst2_LFInst_11_LFInst_1_U6  ( .A1(
        \SubCellInst2_LFInst_11_LFInst_1_n6 ), .A2(
        \SubCellInst2_LFInst_11_LFInst_1_n5 ), .ZN(Feedback2[45]) );
  NAND2_X1 \SubCellInst2_LFInst_11_LFInst_1_U5  ( .A1(PermutationOutput2[46]), 
        .A2(PermutationOutput2[44]), .ZN(\SubCellInst2_LFInst_11_LFInst_1_n5 )
         );
  OR2_X1 \SubCellInst2_LFInst_11_LFInst_1_U4  ( .A1(PermutationOutput2[47]), 
        .A2(\SubCellInst2_LFInst_11_LFInst_1_n4 ), .ZN(
        \SubCellInst2_LFInst_11_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst2_LFInst_11_LFInst_1_U3  ( .A1(PermutationOutput2[46]), 
        .A2(PermutationOutput2[44]), .ZN(\SubCellInst2_LFInst_11_LFInst_1_n4 )
         );
  NAND2_X1 \SubCellInst2_LFInst_11_LFInst_2_U8  ( .A1(
        \SubCellInst2_LFInst_11_LFInst_2_n11 ), .A2(
        \SubCellInst2_LFInst_11_LFInst_2_n10 ), .ZN(Feedback2[46]) );
  OR2_X1 \SubCellInst2_LFInst_11_LFInst_2_U7  ( .A1(PermutationOutput2[44]), 
        .A2(PermutationOutput2[47]), .ZN(\SubCellInst2_LFInst_11_LFInst_2_n10 ) );
  NAND2_X1 \SubCellInst2_LFInst_11_LFInst_2_U6  ( .A1(PermutationOutput2[45]), 
        .A2(\SubCellInst2_LFInst_11_LFInst_2_n9 ), .ZN(
        \SubCellInst2_LFInst_11_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst2_LFInst_11_LFInst_2_U5  ( .A1(
        \SubCellInst2_LFInst_11_LFInst_2_n8 ), .A2(
        \SubCellInst2_LFInst_11_LFInst_2_n7 ), .ZN(
        \SubCellInst2_LFInst_11_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst2_LFInst_11_LFInst_2_U4  ( .A1(PermutationOutput2[44]), 
        .A2(PermutationOutput2[47]), .ZN(\SubCellInst2_LFInst_11_LFInst_2_n7 )
         );
  INV_X1 \SubCellInst2_LFInst_11_LFInst_2_U3  ( .A(PermutationOutput2[46]), 
        .ZN(\SubCellInst2_LFInst_11_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst2_LFInst_11_LFInst_3_U6  ( .A1(
        \SubCellInst2_LFInst_11_LFInst_3_n6 ), .A2(
        \SubCellInst2_LFInst_11_LFInst_3_n5 ), .ZN(Feedback2[47]) );
  NOR2_X1 \SubCellInst2_LFInst_11_LFInst_3_U5  ( .A1(PermutationOutput2[47]), 
        .A2(PermutationOutput2[44]), .ZN(\SubCellInst2_LFInst_11_LFInst_3_n5 )
         );
  NOR2_X1 \SubCellInst2_LFInst_11_LFInst_3_U4  ( .A1(PermutationOutput2[45]), 
        .A2(\SubCellInst2_LFInst_11_LFInst_3_n4 ), .ZN(
        \SubCellInst2_LFInst_11_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst2_LFInst_11_LFInst_3_U3  ( .A1(PermutationOutput2[47]), 
        .A2(PermutationOutput2[46]), .ZN(\SubCellInst2_LFInst_11_LFInst_3_n4 )
         );
  NOR2_X1 \SubCellInst2_LFInst_12_LFInst_0_U8  ( .A1(
        \SubCellInst2_LFInst_12_LFInst_0_n11 ), .A2(
        \SubCellInst2_LFInst_12_LFInst_0_n10 ), .ZN(Feedback2[48]) );
  AND2_X1 \SubCellInst2_LFInst_12_LFInst_0_U7  ( .A1(PermutationOutput2[51]), 
        .A2(PermutationOutput2[50]), .ZN(\SubCellInst2_LFInst_12_LFInst_0_n10 ) );
  NOR2_X1 \SubCellInst2_LFInst_12_LFInst_0_U6  ( .A1(PermutationOutput2[49]), 
        .A2(\SubCellInst2_LFInst_12_LFInst_0_n9 ), .ZN(
        \SubCellInst2_LFInst_12_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst2_LFInst_12_LFInst_0_U5  ( .A1(
        \SubCellInst2_LFInst_12_LFInst_0_n8 ), .A2(
        \SubCellInst2_LFInst_12_LFInst_0_n7 ), .ZN(
        \SubCellInst2_LFInst_12_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst2_LFInst_12_LFInst_0_U4  ( .A1(PermutationOutput2[51]), 
        .A2(PermutationOutput2[50]), .ZN(\SubCellInst2_LFInst_12_LFInst_0_n7 )
         );
  INV_X1 \SubCellInst2_LFInst_12_LFInst_0_U3  ( .A(PermutationOutput2[48]), 
        .ZN(\SubCellInst2_LFInst_12_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst2_LFInst_12_LFInst_1_U6  ( .A1(
        \SubCellInst2_LFInst_12_LFInst_1_n6 ), .A2(
        \SubCellInst2_LFInst_12_LFInst_1_n5 ), .ZN(Feedback2[49]) );
  NAND2_X1 \SubCellInst2_LFInst_12_LFInst_1_U5  ( .A1(PermutationOutput2[50]), 
        .A2(PermutationOutput2[48]), .ZN(\SubCellInst2_LFInst_12_LFInst_1_n5 )
         );
  OR2_X1 \SubCellInst2_LFInst_12_LFInst_1_U4  ( .A1(PermutationOutput2[51]), 
        .A2(\SubCellInst2_LFInst_12_LFInst_1_n4 ), .ZN(
        \SubCellInst2_LFInst_12_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst2_LFInst_12_LFInst_1_U3  ( .A1(PermutationOutput2[50]), 
        .A2(PermutationOutput2[48]), .ZN(\SubCellInst2_LFInst_12_LFInst_1_n4 )
         );
  NAND2_X1 \SubCellInst2_LFInst_12_LFInst_2_U8  ( .A1(
        \SubCellInst2_LFInst_12_LFInst_2_n11 ), .A2(
        \SubCellInst2_LFInst_12_LFInst_2_n10 ), .ZN(Feedback2[50]) );
  OR2_X1 \SubCellInst2_LFInst_12_LFInst_2_U7  ( .A1(PermutationOutput2[48]), 
        .A2(PermutationOutput2[51]), .ZN(\SubCellInst2_LFInst_12_LFInst_2_n10 ) );
  NAND2_X1 \SubCellInst2_LFInst_12_LFInst_2_U6  ( .A1(PermutationOutput2[49]), 
        .A2(\SubCellInst2_LFInst_12_LFInst_2_n9 ), .ZN(
        \SubCellInst2_LFInst_12_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst2_LFInst_12_LFInst_2_U5  ( .A1(
        \SubCellInst2_LFInst_12_LFInst_2_n8 ), .A2(
        \SubCellInst2_LFInst_12_LFInst_2_n7 ), .ZN(
        \SubCellInst2_LFInst_12_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst2_LFInst_12_LFInst_2_U4  ( .A1(PermutationOutput2[48]), 
        .A2(PermutationOutput2[51]), .ZN(\SubCellInst2_LFInst_12_LFInst_2_n7 )
         );
  INV_X1 \SubCellInst2_LFInst_12_LFInst_2_U3  ( .A(PermutationOutput2[50]), 
        .ZN(\SubCellInst2_LFInst_12_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst2_LFInst_12_LFInst_3_U6  ( .A1(
        \SubCellInst2_LFInst_12_LFInst_3_n6 ), .A2(
        \SubCellInst2_LFInst_12_LFInst_3_n5 ), .ZN(Feedback2[51]) );
  NOR2_X1 \SubCellInst2_LFInst_12_LFInst_3_U5  ( .A1(PermutationOutput2[51]), 
        .A2(PermutationOutput2[48]), .ZN(\SubCellInst2_LFInst_12_LFInst_3_n5 )
         );
  NOR2_X1 \SubCellInst2_LFInst_12_LFInst_3_U4  ( .A1(PermutationOutput2[49]), 
        .A2(\SubCellInst2_LFInst_12_LFInst_3_n4 ), .ZN(
        \SubCellInst2_LFInst_12_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst2_LFInst_12_LFInst_3_U3  ( .A1(PermutationOutput2[51]), 
        .A2(PermutationOutput2[50]), .ZN(\SubCellInst2_LFInst_12_LFInst_3_n4 )
         );
  NOR2_X1 \SubCellInst2_LFInst_13_LFInst_0_U8  ( .A1(
        \SubCellInst2_LFInst_13_LFInst_0_n11 ), .A2(
        \SubCellInst2_LFInst_13_LFInst_0_n10 ), .ZN(Feedback2[52]) );
  AND2_X1 \SubCellInst2_LFInst_13_LFInst_0_U7  ( .A1(PermutationOutput2[55]), 
        .A2(PermutationOutput2[54]), .ZN(\SubCellInst2_LFInst_13_LFInst_0_n10 ) );
  NOR2_X1 \SubCellInst2_LFInst_13_LFInst_0_U6  ( .A1(PermutationOutput2[53]), 
        .A2(\SubCellInst2_LFInst_13_LFInst_0_n9 ), .ZN(
        \SubCellInst2_LFInst_13_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst2_LFInst_13_LFInst_0_U5  ( .A1(
        \SubCellInst2_LFInst_13_LFInst_0_n8 ), .A2(
        \SubCellInst2_LFInst_13_LFInst_0_n7 ), .ZN(
        \SubCellInst2_LFInst_13_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst2_LFInst_13_LFInst_0_U4  ( .A1(PermutationOutput2[55]), 
        .A2(PermutationOutput2[54]), .ZN(\SubCellInst2_LFInst_13_LFInst_0_n7 )
         );
  INV_X1 \SubCellInst2_LFInst_13_LFInst_0_U3  ( .A(PermutationOutput2[52]), 
        .ZN(\SubCellInst2_LFInst_13_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst2_LFInst_13_LFInst_1_U6  ( .A1(
        \SubCellInst2_LFInst_13_LFInst_1_n6 ), .A2(
        \SubCellInst2_LFInst_13_LFInst_1_n5 ), .ZN(Feedback2[53]) );
  NAND2_X1 \SubCellInst2_LFInst_13_LFInst_1_U5  ( .A1(PermutationOutput2[54]), 
        .A2(PermutationOutput2[52]), .ZN(\SubCellInst2_LFInst_13_LFInst_1_n5 )
         );
  OR2_X1 \SubCellInst2_LFInst_13_LFInst_1_U4  ( .A1(PermutationOutput2[55]), 
        .A2(\SubCellInst2_LFInst_13_LFInst_1_n4 ), .ZN(
        \SubCellInst2_LFInst_13_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst2_LFInst_13_LFInst_1_U3  ( .A1(PermutationOutput2[54]), 
        .A2(PermutationOutput2[52]), .ZN(\SubCellInst2_LFInst_13_LFInst_1_n4 )
         );
  NAND2_X1 \SubCellInst2_LFInst_13_LFInst_2_U8  ( .A1(
        \SubCellInst2_LFInst_13_LFInst_2_n11 ), .A2(
        \SubCellInst2_LFInst_13_LFInst_2_n10 ), .ZN(Feedback2[54]) );
  OR2_X1 \SubCellInst2_LFInst_13_LFInst_2_U7  ( .A1(PermutationOutput2[52]), 
        .A2(PermutationOutput2[55]), .ZN(\SubCellInst2_LFInst_13_LFInst_2_n10 ) );
  NAND2_X1 \SubCellInst2_LFInst_13_LFInst_2_U6  ( .A1(PermutationOutput2[53]), 
        .A2(\SubCellInst2_LFInst_13_LFInst_2_n9 ), .ZN(
        \SubCellInst2_LFInst_13_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst2_LFInst_13_LFInst_2_U5  ( .A1(
        \SubCellInst2_LFInst_13_LFInst_2_n8 ), .A2(
        \SubCellInst2_LFInst_13_LFInst_2_n7 ), .ZN(
        \SubCellInst2_LFInst_13_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst2_LFInst_13_LFInst_2_U4  ( .A1(PermutationOutput2[52]), 
        .A2(PermutationOutput2[55]), .ZN(\SubCellInst2_LFInst_13_LFInst_2_n7 )
         );
  INV_X1 \SubCellInst2_LFInst_13_LFInst_2_U3  ( .A(PermutationOutput2[54]), 
        .ZN(\SubCellInst2_LFInst_13_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst2_LFInst_13_LFInst_3_U6  ( .A1(
        \SubCellInst2_LFInst_13_LFInst_3_n6 ), .A2(
        \SubCellInst2_LFInst_13_LFInst_3_n5 ), .ZN(Feedback2[55]) );
  NOR2_X1 \SubCellInst2_LFInst_13_LFInst_3_U5  ( .A1(PermutationOutput2[55]), 
        .A2(PermutationOutput2[52]), .ZN(\SubCellInst2_LFInst_13_LFInst_3_n5 )
         );
  NOR2_X1 \SubCellInst2_LFInst_13_LFInst_3_U4  ( .A1(PermutationOutput2[53]), 
        .A2(\SubCellInst2_LFInst_13_LFInst_3_n4 ), .ZN(
        \SubCellInst2_LFInst_13_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst2_LFInst_13_LFInst_3_U3  ( .A1(PermutationOutput2[55]), 
        .A2(PermutationOutput2[54]), .ZN(\SubCellInst2_LFInst_13_LFInst_3_n4 )
         );
  NOR2_X1 \SubCellInst2_LFInst_14_LFInst_0_U8  ( .A1(
        \SubCellInst2_LFInst_14_LFInst_0_n11 ), .A2(
        \SubCellInst2_LFInst_14_LFInst_0_n10 ), .ZN(Feedback2[56]) );
  AND2_X1 \SubCellInst2_LFInst_14_LFInst_0_U7  ( .A1(PermutationOutput2[59]), 
        .A2(PermutationOutput2[58]), .ZN(\SubCellInst2_LFInst_14_LFInst_0_n10 ) );
  NOR2_X1 \SubCellInst2_LFInst_14_LFInst_0_U6  ( .A1(PermutationOutput2[57]), 
        .A2(\SubCellInst2_LFInst_14_LFInst_0_n9 ), .ZN(
        \SubCellInst2_LFInst_14_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst2_LFInst_14_LFInst_0_U5  ( .A1(
        \SubCellInst2_LFInst_14_LFInst_0_n8 ), .A2(
        \SubCellInst2_LFInst_14_LFInst_0_n7 ), .ZN(
        \SubCellInst2_LFInst_14_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst2_LFInst_14_LFInst_0_U4  ( .A1(PermutationOutput2[59]), 
        .A2(PermutationOutput2[58]), .ZN(\SubCellInst2_LFInst_14_LFInst_0_n7 )
         );
  INV_X1 \SubCellInst2_LFInst_14_LFInst_0_U3  ( .A(PermutationOutput2[56]), 
        .ZN(\SubCellInst2_LFInst_14_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst2_LFInst_14_LFInst_1_U6  ( .A1(
        \SubCellInst2_LFInst_14_LFInst_1_n6 ), .A2(
        \SubCellInst2_LFInst_14_LFInst_1_n5 ), .ZN(Feedback2[57]) );
  NAND2_X1 \SubCellInst2_LFInst_14_LFInst_1_U5  ( .A1(PermutationOutput2[58]), 
        .A2(PermutationOutput2[56]), .ZN(\SubCellInst2_LFInst_14_LFInst_1_n5 )
         );
  OR2_X1 \SubCellInst2_LFInst_14_LFInst_1_U4  ( .A1(PermutationOutput2[59]), 
        .A2(\SubCellInst2_LFInst_14_LFInst_1_n4 ), .ZN(
        \SubCellInst2_LFInst_14_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst2_LFInst_14_LFInst_1_U3  ( .A1(PermutationOutput2[58]), 
        .A2(PermutationOutput2[56]), .ZN(\SubCellInst2_LFInst_14_LFInst_1_n4 )
         );
  NAND2_X1 \SubCellInst2_LFInst_14_LFInst_2_U8  ( .A1(
        \SubCellInst2_LFInst_14_LFInst_2_n11 ), .A2(
        \SubCellInst2_LFInst_14_LFInst_2_n10 ), .ZN(Feedback2[58]) );
  OR2_X1 \SubCellInst2_LFInst_14_LFInst_2_U7  ( .A1(PermutationOutput2[56]), 
        .A2(PermutationOutput2[59]), .ZN(\SubCellInst2_LFInst_14_LFInst_2_n10 ) );
  NAND2_X1 \SubCellInst2_LFInst_14_LFInst_2_U6  ( .A1(PermutationOutput2[57]), 
        .A2(\SubCellInst2_LFInst_14_LFInst_2_n9 ), .ZN(
        \SubCellInst2_LFInst_14_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst2_LFInst_14_LFInst_2_U5  ( .A1(
        \SubCellInst2_LFInst_14_LFInst_2_n8 ), .A2(
        \SubCellInst2_LFInst_14_LFInst_2_n7 ), .ZN(
        \SubCellInst2_LFInst_14_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst2_LFInst_14_LFInst_2_U4  ( .A1(PermutationOutput2[56]), 
        .A2(PermutationOutput2[59]), .ZN(\SubCellInst2_LFInst_14_LFInst_2_n7 )
         );
  INV_X1 \SubCellInst2_LFInst_14_LFInst_2_U3  ( .A(PermutationOutput2[58]), 
        .ZN(\SubCellInst2_LFInst_14_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst2_LFInst_14_LFInst_3_U6  ( .A1(
        \SubCellInst2_LFInst_14_LFInst_3_n6 ), .A2(
        \SubCellInst2_LFInst_14_LFInst_3_n5 ), .ZN(Feedback2[59]) );
  NOR2_X1 \SubCellInst2_LFInst_14_LFInst_3_U5  ( .A1(PermutationOutput2[59]), 
        .A2(PermutationOutput2[56]), .ZN(\SubCellInst2_LFInst_14_LFInst_3_n5 )
         );
  NOR2_X1 \SubCellInst2_LFInst_14_LFInst_3_U4  ( .A1(PermutationOutput2[57]), 
        .A2(\SubCellInst2_LFInst_14_LFInst_3_n4 ), .ZN(
        \SubCellInst2_LFInst_14_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst2_LFInst_14_LFInst_3_U3  ( .A1(PermutationOutput2[59]), 
        .A2(PermutationOutput2[58]), .ZN(\SubCellInst2_LFInst_14_LFInst_3_n4 )
         );
  NOR2_X1 \SubCellInst2_LFInst_15_LFInst_0_U8  ( .A1(
        \SubCellInst2_LFInst_15_LFInst_0_n11 ), .A2(
        \SubCellInst2_LFInst_15_LFInst_0_n10 ), .ZN(Feedback2[60]) );
  AND2_X1 \SubCellInst2_LFInst_15_LFInst_0_U7  ( .A1(PermutationOutput2[63]), 
        .A2(PermutationOutput2[62]), .ZN(\SubCellInst2_LFInst_15_LFInst_0_n10 ) );
  NOR2_X1 \SubCellInst2_LFInst_15_LFInst_0_U6  ( .A1(PermutationOutput2[61]), 
        .A2(\SubCellInst2_LFInst_15_LFInst_0_n9 ), .ZN(
        \SubCellInst2_LFInst_15_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst2_LFInst_15_LFInst_0_U5  ( .A1(
        \SubCellInst2_LFInst_15_LFInst_0_n8 ), .A2(
        \SubCellInst2_LFInst_15_LFInst_0_n7 ), .ZN(
        \SubCellInst2_LFInst_15_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst2_LFInst_15_LFInst_0_U4  ( .A1(PermutationOutput2[63]), 
        .A2(PermutationOutput2[62]), .ZN(\SubCellInst2_LFInst_15_LFInst_0_n7 )
         );
  INV_X1 \SubCellInst2_LFInst_15_LFInst_0_U3  ( .A(PermutationOutput2[60]), 
        .ZN(\SubCellInst2_LFInst_15_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst2_LFInst_15_LFInst_1_U6  ( .A1(
        \SubCellInst2_LFInst_15_LFInst_1_n6 ), .A2(
        \SubCellInst2_LFInst_15_LFInst_1_n5 ), .ZN(Feedback2[61]) );
  NAND2_X1 \SubCellInst2_LFInst_15_LFInst_1_U5  ( .A1(PermutationOutput2[62]), 
        .A2(PermutationOutput2[60]), .ZN(\SubCellInst2_LFInst_15_LFInst_1_n5 )
         );
  OR2_X1 \SubCellInst2_LFInst_15_LFInst_1_U4  ( .A1(PermutationOutput2[63]), 
        .A2(\SubCellInst2_LFInst_15_LFInst_1_n4 ), .ZN(
        \SubCellInst2_LFInst_15_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst2_LFInst_15_LFInst_1_U3  ( .A1(PermutationOutput2[62]), 
        .A2(PermutationOutput2[60]), .ZN(\SubCellInst2_LFInst_15_LFInst_1_n4 )
         );
  NAND2_X1 \SubCellInst2_LFInst_15_LFInst_2_U8  ( .A1(
        \SubCellInst2_LFInst_15_LFInst_2_n11 ), .A2(
        \SubCellInst2_LFInst_15_LFInst_2_n10 ), .ZN(Feedback2[62]) );
  OR2_X1 \SubCellInst2_LFInst_15_LFInst_2_U7  ( .A1(PermutationOutput2[60]), 
        .A2(PermutationOutput2[63]), .ZN(\SubCellInst2_LFInst_15_LFInst_2_n10 ) );
  NAND2_X1 \SubCellInst2_LFInst_15_LFInst_2_U6  ( .A1(PermutationOutput2[61]), 
        .A2(\SubCellInst2_LFInst_15_LFInst_2_n9 ), .ZN(
        \SubCellInst2_LFInst_15_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst2_LFInst_15_LFInst_2_U5  ( .A1(
        \SubCellInst2_LFInst_15_LFInst_2_n8 ), .A2(
        \SubCellInst2_LFInst_15_LFInst_2_n7 ), .ZN(
        \SubCellInst2_LFInst_15_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst2_LFInst_15_LFInst_2_U4  ( .A1(PermutationOutput2[60]), 
        .A2(PermutationOutput2[63]), .ZN(\SubCellInst2_LFInst_15_LFInst_2_n7 )
         );
  INV_X1 \SubCellInst2_LFInst_15_LFInst_2_U3  ( .A(PermutationOutput2[62]), 
        .ZN(\SubCellInst2_LFInst_15_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst2_LFInst_15_LFInst_3_U6  ( .A1(
        \SubCellInst2_LFInst_15_LFInst_3_n6 ), .A2(
        \SubCellInst2_LFInst_15_LFInst_3_n5 ), .ZN(Feedback2[63]) );
  NOR2_X1 \SubCellInst2_LFInst_15_LFInst_3_U5  ( .A1(PermutationOutput2[63]), 
        .A2(PermutationOutput2[60]), .ZN(\SubCellInst2_LFInst_15_LFInst_3_n5 )
         );
  NOR2_X1 \SubCellInst2_LFInst_15_LFInst_3_U4  ( .A1(PermutationOutput2[61]), 
        .A2(\SubCellInst2_LFInst_15_LFInst_3_n4 ), .ZN(
        \SubCellInst2_LFInst_15_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst2_LFInst_15_LFInst_3_U3  ( .A1(PermutationOutput2[63]), 
        .A2(PermutationOutput2[62]), .ZN(\SubCellInst2_LFInst_15_LFInst_3_n4 )
         );
  XNOR2_X1 \MCInst3_XOR_r0_Inst_0_U2  ( .A(\MCInst3_XOR_r0_Inst_0_n3 ), .B(
        MCOutput3[0]), .ZN(MCOutput3[48]) );
  XNOR2_X1 \MCInst3_XOR_r0_Inst_0_U1  ( .A(Feedback2[48]), .B(MCOutput3[16]), 
        .ZN(\MCInst3_XOR_r0_Inst_0_n3 ) );
  XOR2_X1 \MCInst3_XOR_r1_Inst_0_U1  ( .A(Feedback2[32]), .B(MCOutput3[0]), 
        .Z(MCOutput3[32]) );
  XNOR2_X1 \MCInst3_XOR_r0_Inst_1_U2  ( .A(\MCInst3_XOR_r0_Inst_1_n3 ), .B(
        MCOutput3[1]), .ZN(MCOutput3[49]) );
  XNOR2_X1 \MCInst3_XOR_r0_Inst_1_U1  ( .A(Feedback2[49]), .B(MCOutput3[17]), 
        .ZN(\MCInst3_XOR_r0_Inst_1_n3 ) );
  XOR2_X1 \MCInst3_XOR_r1_Inst_1_U1  ( .A(Feedback2[33]), .B(MCOutput3[1]), 
        .Z(MCOutput3[33]) );
  XNOR2_X1 \MCInst3_XOR_r0_Inst_2_U2  ( .A(\MCInst3_XOR_r0_Inst_2_n3 ), .B(
        MCOutput3[2]), .ZN(MCOutput3[50]) );
  XNOR2_X1 \MCInst3_XOR_r0_Inst_2_U1  ( .A(Feedback2[50]), .B(MCOutput3[18]), 
        .ZN(\MCInst3_XOR_r0_Inst_2_n3 ) );
  XOR2_X1 \MCInst3_XOR_r1_Inst_2_U1  ( .A(Feedback2[34]), .B(MCOutput3[2]), 
        .Z(MCOutput3[34]) );
  XNOR2_X1 \MCInst3_XOR_r0_Inst_3_U2  ( .A(\MCInst3_XOR_r0_Inst_3_n3 ), .B(
        MCOutput3[3]), .ZN(MCOutput3[51]) );
  XNOR2_X1 \MCInst3_XOR_r0_Inst_3_U1  ( .A(Feedback2[51]), .B(MCOutput3[19]), 
        .ZN(\MCInst3_XOR_r0_Inst_3_n3 ) );
  XOR2_X1 \MCInst3_XOR_r1_Inst_3_U1  ( .A(Feedback2[35]), .B(MCOutput3[3]), 
        .Z(MCOutput3[35]) );
  XNOR2_X1 \MCInst3_XOR_r0_Inst_4_U2  ( .A(\MCInst3_XOR_r0_Inst_4_n3 ), .B(
        MCOutput3[4]), .ZN(MCOutput3[52]) );
  XNOR2_X1 \MCInst3_XOR_r0_Inst_4_U1  ( .A(Feedback2[52]), .B(MCOutput3[20]), 
        .ZN(\MCInst3_XOR_r0_Inst_4_n3 ) );
  XOR2_X1 \MCInst3_XOR_r1_Inst_4_U1  ( .A(Feedback2[36]), .B(MCOutput3[4]), 
        .Z(MCOutput3[36]) );
  XNOR2_X1 \MCInst3_XOR_r0_Inst_5_U2  ( .A(\MCInst3_XOR_r0_Inst_5_n3 ), .B(
        MCOutput3[5]), .ZN(MCOutput3[53]) );
  XNOR2_X1 \MCInst3_XOR_r0_Inst_5_U1  ( .A(Feedback2[53]), .B(MCOutput3[21]), 
        .ZN(\MCInst3_XOR_r0_Inst_5_n3 ) );
  XOR2_X1 \MCInst3_XOR_r1_Inst_5_U1  ( .A(Feedback2[37]), .B(MCOutput3[5]), 
        .Z(MCOutput3[37]) );
  XNOR2_X1 \MCInst3_XOR_r0_Inst_6_U2  ( .A(\MCInst3_XOR_r0_Inst_6_n3 ), .B(
        MCOutput3[6]), .ZN(MCOutput3[54]) );
  XNOR2_X1 \MCInst3_XOR_r0_Inst_6_U1  ( .A(Feedback2[54]), .B(MCOutput3[22]), 
        .ZN(\MCInst3_XOR_r0_Inst_6_n3 ) );
  XOR2_X1 \MCInst3_XOR_r1_Inst_6_U1  ( .A(Feedback2[38]), .B(MCOutput3[6]), 
        .Z(MCOutput3[38]) );
  XNOR2_X1 \MCInst3_XOR_r0_Inst_7_U2  ( .A(\MCInst3_XOR_r0_Inst_7_n3 ), .B(
        MCOutput3[7]), .ZN(MCOutput3[55]) );
  XNOR2_X1 \MCInst3_XOR_r0_Inst_7_U1  ( .A(Feedback2[55]), .B(MCOutput3[23]), 
        .ZN(\MCInst3_XOR_r0_Inst_7_n3 ) );
  XOR2_X1 \MCInst3_XOR_r1_Inst_7_U1  ( .A(Feedback2[39]), .B(MCOutput3[7]), 
        .Z(MCOutput3[39]) );
  XNOR2_X1 \MCInst3_XOR_r0_Inst_8_U2  ( .A(\MCInst3_XOR_r0_Inst_8_n3 ), .B(
        MCOutput3[8]), .ZN(MCOutput3[56]) );
  XNOR2_X1 \MCInst3_XOR_r0_Inst_8_U1  ( .A(Feedback2[56]), .B(MCOutput3[24]), 
        .ZN(\MCInst3_XOR_r0_Inst_8_n3 ) );
  XOR2_X1 \MCInst3_XOR_r1_Inst_8_U1  ( .A(Feedback2[40]), .B(MCOutput3[8]), 
        .Z(MCOutput3[40]) );
  XNOR2_X1 \MCInst3_XOR_r0_Inst_9_U2  ( .A(\MCInst3_XOR_r0_Inst_9_n3 ), .B(
        MCOutput3[9]), .ZN(MCOutput3[57]) );
  XNOR2_X1 \MCInst3_XOR_r0_Inst_9_U1  ( .A(Feedback2[57]), .B(MCOutput3[25]), 
        .ZN(\MCInst3_XOR_r0_Inst_9_n3 ) );
  XOR2_X1 \MCInst3_XOR_r1_Inst_9_U1  ( .A(Feedback2[41]), .B(MCOutput3[9]), 
        .Z(MCOutput3[41]) );
  XNOR2_X1 \MCInst3_XOR_r0_Inst_10_U2  ( .A(\MCInst3_XOR_r0_Inst_10_n3 ), .B(
        MCOutput3[10]), .ZN(MCOutput3[58]) );
  XNOR2_X1 \MCInst3_XOR_r0_Inst_10_U1  ( .A(Feedback2[58]), .B(MCOutput3[26]), 
        .ZN(\MCInst3_XOR_r0_Inst_10_n3 ) );
  XOR2_X1 \MCInst3_XOR_r1_Inst_10_U1  ( .A(Feedback2[42]), .B(MCOutput3[10]), 
        .Z(MCOutput3[42]) );
  XNOR2_X1 \MCInst3_XOR_r0_Inst_11_U2  ( .A(\MCInst3_XOR_r0_Inst_11_n3 ), .B(
        MCOutput3[11]), .ZN(MCOutput3[59]) );
  XNOR2_X1 \MCInst3_XOR_r0_Inst_11_U1  ( .A(Feedback2[59]), .B(MCOutput3[27]), 
        .ZN(\MCInst3_XOR_r0_Inst_11_n3 ) );
  XOR2_X1 \MCInst3_XOR_r1_Inst_11_U1  ( .A(Feedback2[43]), .B(MCOutput3[11]), 
        .Z(MCOutput3[43]) );
  XNOR2_X1 \MCInst3_XOR_r0_Inst_12_U2  ( .A(\MCInst3_XOR_r0_Inst_12_n3 ), .B(
        MCOutput3[12]), .ZN(MCOutput3[60]) );
  XNOR2_X1 \MCInst3_XOR_r0_Inst_12_U1  ( .A(Feedback2[60]), .B(MCOutput3[28]), 
        .ZN(\MCInst3_XOR_r0_Inst_12_n3 ) );
  XOR2_X1 \MCInst3_XOR_r1_Inst_12_U1  ( .A(Feedback2[44]), .B(MCOutput3[12]), 
        .Z(MCOutput3[44]) );
  XNOR2_X1 \MCInst3_XOR_r0_Inst_13_U2  ( .A(\MCInst3_XOR_r0_Inst_13_n3 ), .B(
        MCOutput3[13]), .ZN(MCOutput3[61]) );
  XNOR2_X1 \MCInst3_XOR_r0_Inst_13_U1  ( .A(Feedback2[61]), .B(MCOutput3[29]), 
        .ZN(\MCInst3_XOR_r0_Inst_13_n3 ) );
  XOR2_X1 \MCInst3_XOR_r1_Inst_13_U1  ( .A(Feedback2[45]), .B(MCOutput3[13]), 
        .Z(MCOutput3[45]) );
  XNOR2_X1 \MCInst3_XOR_r0_Inst_14_U2  ( .A(\MCInst3_XOR_r0_Inst_14_n3 ), .B(
        MCOutput3[14]), .ZN(MCOutput3[62]) );
  XNOR2_X1 \MCInst3_XOR_r0_Inst_14_U1  ( .A(Feedback2[62]), .B(MCOutput3[30]), 
        .ZN(\MCInst3_XOR_r0_Inst_14_n3 ) );
  XOR2_X1 \MCInst3_XOR_r1_Inst_14_U1  ( .A(Feedback2[46]), .B(MCOutput3[14]), 
        .Z(MCOutput3[46]) );
  XNOR2_X1 \MCInst3_XOR_r0_Inst_15_U2  ( .A(\MCInst3_XOR_r0_Inst_15_n3 ), .B(
        MCOutput3[15]), .ZN(MCOutput3[63]) );
  XNOR2_X1 \MCInst3_XOR_r0_Inst_15_U1  ( .A(Feedback2[63]), .B(MCOutput3[31]), 
        .ZN(\MCInst3_XOR_r0_Inst_15_n3 ) );
  XOR2_X1 \MCInst3_XOR_r1_Inst_15_U1  ( .A(Feedback2[47]), .B(MCOutput3[15]), 
        .Z(MCOutput3[47]) );
  XOR2_X1 \AddKeyXOR13_XORInst_0_0_U1  ( .A(MCOutput3[48]), .B(Key[48]), .Z(
        AddRoundKeyOutput3[48]) );
  XOR2_X1 \AddKeyXOR13_XORInst_0_1_U1  ( .A(MCOutput3[49]), .B(Key[49]), .Z(
        AddRoundKeyOutput3[49]) );
  XOR2_X1 \AddKeyXOR13_XORInst_0_2_U1  ( .A(MCOutput3[50]), .B(Key[50]), .Z(
        AddRoundKeyOutput3[50]) );
  XOR2_X1 \AddKeyXOR13_XORInst_0_3_U1  ( .A(MCOutput3[51]), .B(Key[51]), .Z(
        AddRoundKeyOutput3[51]) );
  XOR2_X1 \AddKeyXOR13_XORInst_1_0_U1  ( .A(MCOutput3[52]), .B(Key[52]), .Z(
        AddRoundKeyOutput3[52]) );
  XOR2_X1 \AddKeyXOR13_XORInst_1_1_U1  ( .A(MCOutput3[53]), .B(Key[53]), .Z(
        AddRoundKeyOutput3[53]) );
  XOR2_X1 \AddKeyXOR13_XORInst_1_2_U1  ( .A(MCOutput3[54]), .B(Key[54]), .Z(
        AddRoundKeyOutput3[54]) );
  XOR2_X1 \AddKeyXOR13_XORInst_1_3_U1  ( .A(MCOutput3[55]), .B(Key[55]), .Z(
        AddRoundKeyOutput3[55]) );
  XOR2_X1 \AddKeyXOR13_XORInst_2_0_U1  ( .A(MCOutput3[56]), .B(Key[56]), .Z(
        AddRoundKeyOutput3[56]) );
  XOR2_X1 \AddKeyXOR13_XORInst_2_1_U1  ( .A(MCOutput3[57]), .B(Key[57]), .Z(
        AddRoundKeyOutput3[57]) );
  XOR2_X1 \AddKeyXOR13_XORInst_2_2_U1  ( .A(MCOutput3[58]), .B(Key[58]), .Z(
        AddRoundKeyOutput3[58]) );
  XOR2_X1 \AddKeyXOR13_XORInst_2_3_U1  ( .A(MCOutput3[59]), .B(Key[59]), .Z(
        AddRoundKeyOutput3[59]) );
  XOR2_X1 \AddKeyXOR13_XORInst_3_0_U1  ( .A(MCOutput3[60]), .B(Key[60]), .Z(
        AddRoundKeyOutput3[60]) );
  XOR2_X1 \AddKeyXOR13_XORInst_3_1_U1  ( .A(MCOutput3[61]), .B(Key[61]), .Z(
        AddRoundKeyOutput3[61]) );
  XOR2_X1 \AddKeyXOR13_XORInst_3_2_U1  ( .A(MCOutput3[62]), .B(Key[62]), .Z(
        AddRoundKeyOutput3[62]) );
  XOR2_X1 \AddKeyXOR13_XORInst_3_3_U1  ( .A(MCOutput3[63]), .B(Key[63]), .Z(
        AddRoundKeyOutput3[63]) );
  XOR2_X1 \AddKeyConstXOR3_XORInst_0_0_U1  ( .A(Key[40]), .B(MCOutput3[40]), 
        .Z(AddRoundKeyOutput3[40]) );
  XOR2_X1 \AddKeyConstXOR3_XORInst_0_1_U1  ( .A(Key[41]), .B(MCOutput3[41]), 
        .Z(AddRoundKeyOutput3[41]) );
  XOR2_X1 \AddKeyConstXOR3_XORInst_0_2_U1  ( .A(Key[42]), .B(MCOutput3[42]), 
        .Z(AddRoundKeyOutput3[42]) );
  XOR2_X1 \AddKeyConstXOR3_XORInst_0_3_U1  ( .A(Key[43]), .B(MCOutput3[43]), 
        .Z(AddRoundKeyOutput3[43]) );
  XOR2_X1 \AddKeyConstXOR3_XORInst_1_0_U1  ( .A(Key[44]), .B(MCOutput3[44]), 
        .Z(AddRoundKeyOutput3[44]) );
  XOR2_X1 \AddKeyConstXOR3_XORInst_1_1_U1  ( .A(Key[45]), .B(MCOutput3[45]), 
        .Z(AddRoundKeyOutput3[45]) );
  XOR2_X1 \AddKeyConstXOR3_XORInst_1_2_U1  ( .A(Key[46]), .B(MCOutput3[46]), 
        .Z(AddRoundKeyOutput3[46]) );
  XOR2_X1 \AddKeyConstXOR3_XORInst_1_3_U1  ( .A(Key[47]), .B(MCOutput3[47]), 
        .Z(AddRoundKeyOutput3[47]) );
  XOR2_X1 \AddKeyXOR23_XORInst_0_0_U1  ( .A(MCOutput3[0]), .B(Key[0]), .Z(
        AddRoundKeyOutput3[0]) );
  XOR2_X1 \AddKeyXOR23_XORInst_0_1_U1  ( .A(MCOutput3[1]), .B(Key[1]), .Z(
        AddRoundKeyOutput3[1]) );
  XOR2_X1 \AddKeyXOR23_XORInst_0_2_U1  ( .A(MCOutput3[2]), .B(Key[2]), .Z(
        AddRoundKeyOutput3[2]) );
  XOR2_X1 \AddKeyXOR23_XORInst_0_3_U1  ( .A(MCOutput3[3]), .B(Key[3]), .Z(
        AddRoundKeyOutput3[3]) );
  XOR2_X1 \AddKeyXOR23_XORInst_1_0_U1  ( .A(MCOutput3[4]), .B(Key[4]), .Z(
        AddRoundKeyOutput3[4]) );
  XOR2_X1 \AddKeyXOR23_XORInst_1_1_U1  ( .A(MCOutput3[5]), .B(Key[5]), .Z(
        AddRoundKeyOutput3[5]) );
  XOR2_X1 \AddKeyXOR23_XORInst_1_2_U1  ( .A(MCOutput3[6]), .B(Key[6]), .Z(
        AddRoundKeyOutput3[6]) );
  XOR2_X1 \AddKeyXOR23_XORInst_1_3_U1  ( .A(MCOutput3[7]), .B(Key[7]), .Z(
        AddRoundKeyOutput3[7]) );
  XOR2_X1 \AddKeyXOR23_XORInst_2_0_U1  ( .A(MCOutput3[8]), .B(Key[8]), .Z(
        AddRoundKeyOutput3[8]) );
  XOR2_X1 \AddKeyXOR23_XORInst_2_1_U1  ( .A(MCOutput3[9]), .B(Key[9]), .Z(
        AddRoundKeyOutput3[9]) );
  XOR2_X1 \AddKeyXOR23_XORInst_2_2_U1  ( .A(MCOutput3[10]), .B(Key[10]), .Z(
        AddRoundKeyOutput3[10]) );
  XOR2_X1 \AddKeyXOR23_XORInst_2_3_U1  ( .A(MCOutput3[11]), .B(Key[11]), .Z(
        AddRoundKeyOutput3[11]) );
  XOR2_X1 \AddKeyXOR23_XORInst_3_0_U1  ( .A(MCOutput3[12]), .B(Key[12]), .Z(
        AddRoundKeyOutput3[12]) );
  XOR2_X1 \AddKeyXOR23_XORInst_3_1_U1  ( .A(MCOutput3[13]), .B(Key[13]), .Z(
        AddRoundKeyOutput3[13]) );
  XOR2_X1 \AddKeyXOR23_XORInst_3_2_U1  ( .A(MCOutput3[14]), .B(Key[14]), .Z(
        AddRoundKeyOutput3[14]) );
  XOR2_X1 \AddKeyXOR23_XORInst_3_3_U1  ( .A(MCOutput3[15]), .B(Key[15]), .Z(
        AddRoundKeyOutput3[15]) );
  XOR2_X1 \AddKeyXOR23_XORInst_4_0_U1  ( .A(MCOutput3[16]), .B(Key[16]), .Z(
        AddRoundKeyOutput3[16]) );
  XOR2_X1 \AddKeyXOR23_XORInst_4_1_U1  ( .A(MCOutput3[17]), .B(Key[17]), .Z(
        AddRoundKeyOutput3[17]) );
  XOR2_X1 \AddKeyXOR23_XORInst_4_2_U1  ( .A(MCOutput3[18]), .B(Key[18]), .Z(
        AddRoundKeyOutput3[18]) );
  XOR2_X1 \AddKeyXOR23_XORInst_4_3_U1  ( .A(MCOutput3[19]), .B(Key[19]), .Z(
        AddRoundKeyOutput3[19]) );
  XOR2_X1 \AddKeyXOR23_XORInst_5_0_U1  ( .A(MCOutput3[20]), .B(Key[20]), .Z(
        AddRoundKeyOutput3[20]) );
  XOR2_X1 \AddKeyXOR23_XORInst_5_1_U1  ( .A(MCOutput3[21]), .B(Key[21]), .Z(
        AddRoundKeyOutput3[21]) );
  XOR2_X1 \AddKeyXOR23_XORInst_5_2_U1  ( .A(MCOutput3[22]), .B(Key[22]), .Z(
        AddRoundKeyOutput3[22]) );
  XOR2_X1 \AddKeyXOR23_XORInst_5_3_U1  ( .A(MCOutput3[23]), .B(Key[23]), .Z(
        AddRoundKeyOutput3[23]) );
  XOR2_X1 \AddKeyXOR23_XORInst_6_0_U1  ( .A(MCOutput3[24]), .B(Key[24]), .Z(
        AddRoundKeyOutput3[24]) );
  XOR2_X1 \AddKeyXOR23_XORInst_6_1_U1  ( .A(MCOutput3[25]), .B(Key[25]), .Z(
        AddRoundKeyOutput3[25]) );
  XOR2_X1 \AddKeyXOR23_XORInst_6_2_U1  ( .A(MCOutput3[26]), .B(Key[26]), .Z(
        AddRoundKeyOutput3[26]) );
  XOR2_X1 \AddKeyXOR23_XORInst_6_3_U1  ( .A(MCOutput3[27]), .B(Key[27]), .Z(
        AddRoundKeyOutput3[27]) );
  XOR2_X1 \AddKeyXOR23_XORInst_7_0_U1  ( .A(MCOutput3[28]), .B(Key[28]), .Z(
        AddRoundKeyOutput3[28]) );
  XOR2_X1 \AddKeyXOR23_XORInst_7_1_U1  ( .A(MCOutput3[29]), .B(Key[29]), .Z(
        AddRoundKeyOutput3[29]) );
  XOR2_X1 \AddKeyXOR23_XORInst_7_2_U1  ( .A(MCOutput3[30]), .B(Key[30]), .Z(
        AddRoundKeyOutput3[30]) );
  XOR2_X1 \AddKeyXOR23_XORInst_7_3_U1  ( .A(MCOutput3[31]), .B(Key[31]), .Z(
        AddRoundKeyOutput3[31]) );
  XOR2_X1 \AddKeyXOR23_XORInst_8_0_U1  ( .A(MCOutput3[32]), .B(Key[32]), .Z(
        AddRoundKeyOutput3[32]) );
  XOR2_X1 \AddKeyXOR23_XORInst_8_1_U1  ( .A(MCOutput3[33]), .B(Key[33]), .Z(
        AddRoundKeyOutput3[33]) );
  XOR2_X1 \AddKeyXOR23_XORInst_8_2_U1  ( .A(MCOutput3[34]), .B(Key[34]), .Z(
        AddRoundKeyOutput3[34]) );
  XOR2_X1 \AddKeyXOR23_XORInst_8_3_U1  ( .A(MCOutput3[35]), .B(Key[35]), .Z(
        AddRoundKeyOutput3[35]) );
  XOR2_X1 \AddKeyXOR23_XORInst_9_0_U1  ( .A(MCOutput3[36]), .B(Key[36]), .Z(
        AddRoundKeyOutput3[36]) );
  XOR2_X1 \AddKeyXOR23_XORInst_9_1_U1  ( .A(MCOutput3[37]), .B(Key[37]), .Z(
        AddRoundKeyOutput3[37]) );
  XOR2_X1 \AddKeyXOR23_XORInst_9_2_U1  ( .A(MCOutput3[38]), .B(Key[38]), .Z(
        AddRoundKeyOutput3[38]) );
  XOR2_X1 \AddKeyXOR23_XORInst_9_3_U1  ( .A(MCOutput3[39]), .B(Key[39]), .Z(
        AddRoundKeyOutput3[39]) );
  DFF_X1 \StateReg3_s_current_state_reg[0]  ( .D(AddRoundKeyOutput3[0]), .CK(
        clk), .Q(PermutationOutput3[60]) );
  DFF_X1 \StateReg3_s_current_state_reg[1]  ( .D(AddRoundKeyOutput3[1]), .CK(
        clk), .Q(PermutationOutput3[61]) );
  DFF_X1 \StateReg3_s_current_state_reg[2]  ( .D(AddRoundKeyOutput3[2]), .CK(
        clk), .Q(PermutationOutput3[62]) );
  DFF_X1 \StateReg3_s_current_state_reg[3]  ( .D(AddRoundKeyOutput3[3]), .CK(
        clk), .Q(PermutationOutput3[63]) );
  DFF_X1 \StateReg3_s_current_state_reg[4]  ( .D(AddRoundKeyOutput3[4]), .CK(
        clk), .Q(PermutationOutput3[48]) );
  DFF_X1 \StateReg3_s_current_state_reg[5]  ( .D(AddRoundKeyOutput3[5]), .CK(
        clk), .Q(PermutationOutput3[49]) );
  DFF_X1 \StateReg3_s_current_state_reg[6]  ( .D(AddRoundKeyOutput3[6]), .CK(
        clk), .Q(PermutationOutput3[50]) );
  DFF_X1 \StateReg3_s_current_state_reg[7]  ( .D(AddRoundKeyOutput3[7]), .CK(
        clk), .Q(PermutationOutput3[51]) );
  DFF_X1 \StateReg3_s_current_state_reg[8]  ( .D(AddRoundKeyOutput3[8]), .CK(
        clk), .Q(PermutationOutput3[52]) );
  DFF_X1 \StateReg3_s_current_state_reg[9]  ( .D(AddRoundKeyOutput3[9]), .CK(
        clk), .Q(PermutationOutput3[53]) );
  DFF_X1 \StateReg3_s_current_state_reg[10]  ( .D(AddRoundKeyOutput3[10]), 
        .CK(clk), .Q(PermutationOutput3[54]) );
  DFF_X1 \StateReg3_s_current_state_reg[11]  ( .D(AddRoundKeyOutput3[11]), 
        .CK(clk), .Q(PermutationOutput3[55]) );
  DFF_X1 \StateReg3_s_current_state_reg[12]  ( .D(AddRoundKeyOutput3[12]), 
        .CK(clk), .Q(PermutationOutput3[56]) );
  DFF_X1 \StateReg3_s_current_state_reg[13]  ( .D(AddRoundKeyOutput3[13]), 
        .CK(clk), .Q(PermutationOutput3[57]) );
  DFF_X1 \StateReg3_s_current_state_reg[14]  ( .D(AddRoundKeyOutput3[14]), 
        .CK(clk), .Q(PermutationOutput3[58]) );
  DFF_X1 \StateReg3_s_current_state_reg[15]  ( .D(AddRoundKeyOutput3[15]), 
        .CK(clk), .Q(PermutationOutput3[59]) );
  DFF_X1 \StateReg3_s_current_state_reg[16]  ( .D(AddRoundKeyOutput3[16]), 
        .CK(clk), .Q(PermutationOutput3[32]) );
  DFF_X1 \StateReg3_s_current_state_reg[17]  ( .D(AddRoundKeyOutput3[17]), 
        .CK(clk), .Q(PermutationOutput3[33]) );
  DFF_X1 \StateReg3_s_current_state_reg[18]  ( .D(AddRoundKeyOutput3[18]), 
        .CK(clk), .Q(PermutationOutput3[34]) );
  DFF_X1 \StateReg3_s_current_state_reg[19]  ( .D(AddRoundKeyOutput3[19]), 
        .CK(clk), .Q(PermutationOutput3[35]) );
  DFF_X1 \StateReg3_s_current_state_reg[20]  ( .D(AddRoundKeyOutput3[20]), 
        .CK(clk), .Q(PermutationOutput3[44]) );
  DFF_X1 \StateReg3_s_current_state_reg[21]  ( .D(AddRoundKeyOutput3[21]), 
        .CK(clk), .Q(PermutationOutput3[45]) );
  DFF_X1 \StateReg3_s_current_state_reg[22]  ( .D(AddRoundKeyOutput3[22]), 
        .CK(clk), .Q(PermutationOutput3[46]) );
  DFF_X1 \StateReg3_s_current_state_reg[23]  ( .D(AddRoundKeyOutput3[23]), 
        .CK(clk), .Q(PermutationOutput3[47]) );
  DFF_X1 \StateReg3_s_current_state_reg[24]  ( .D(AddRoundKeyOutput3[24]), 
        .CK(clk), .Q(PermutationOutput3[40]) );
  DFF_X1 \StateReg3_s_current_state_reg[25]  ( .D(AddRoundKeyOutput3[25]), 
        .CK(clk), .Q(PermutationOutput3[41]) );
  DFF_X1 \StateReg3_s_current_state_reg[26]  ( .D(AddRoundKeyOutput3[26]), 
        .CK(clk), .Q(PermutationOutput3[42]) );
  DFF_X1 \StateReg3_s_current_state_reg[27]  ( .D(AddRoundKeyOutput3[27]), 
        .CK(clk), .Q(PermutationOutput3[43]) );
  DFF_X1 \StateReg3_s_current_state_reg[28]  ( .D(AddRoundKeyOutput3[28]), 
        .CK(clk), .Q(PermutationOutput3[36]) );
  DFF_X1 \StateReg3_s_current_state_reg[29]  ( .D(AddRoundKeyOutput3[29]), 
        .CK(clk), .Q(PermutationOutput3[37]) );
  DFF_X1 \StateReg3_s_current_state_reg[30]  ( .D(AddRoundKeyOutput3[30]), 
        .CK(clk), .Q(PermutationOutput3[38]) );
  DFF_X1 \StateReg3_s_current_state_reg[31]  ( .D(AddRoundKeyOutput3[31]), 
        .CK(clk), .Q(PermutationOutput3[39]) );
  DFF_X1 \StateReg3_s_current_state_reg[32]  ( .D(AddRoundKeyOutput3[32]), 
        .CK(clk), .Q(PermutationOutput3[16]) );
  DFF_X1 \StateReg3_s_current_state_reg[33]  ( .D(AddRoundKeyOutput3[33]), 
        .CK(clk), .Q(PermutationOutput3[17]) );
  DFF_X1 \StateReg3_s_current_state_reg[34]  ( .D(AddRoundKeyOutput3[34]), 
        .CK(clk), .Q(PermutationOutput3[18]) );
  DFF_X1 \StateReg3_s_current_state_reg[35]  ( .D(AddRoundKeyOutput3[35]), 
        .CK(clk), .Q(PermutationOutput3[19]) );
  DFF_X1 \StateReg3_s_current_state_reg[36]  ( .D(AddRoundKeyOutput3[36]), 
        .CK(clk), .Q(PermutationOutput3[28]) );
  DFF_X1 \StateReg3_s_current_state_reg[37]  ( .D(AddRoundKeyOutput3[37]), 
        .CK(clk), .Q(PermutationOutput3[29]) );
  DFF_X1 \StateReg3_s_current_state_reg[38]  ( .D(AddRoundKeyOutput3[38]), 
        .CK(clk), .Q(PermutationOutput3[30]) );
  DFF_X1 \StateReg3_s_current_state_reg[39]  ( .D(AddRoundKeyOutput3[39]), 
        .CK(clk), .Q(PermutationOutput3[31]) );
  DFF_X1 \StateReg3_s_current_state_reg[40]  ( .D(AddRoundKeyOutput3[40]), 
        .CK(clk), .Q(PermutationOutput3[24]) );
  DFF_X1 \StateReg3_s_current_state_reg[41]  ( .D(AddRoundKeyOutput3[41]), 
        .CK(clk), .Q(PermutationOutput3[25]) );
  DFF_X1 \StateReg3_s_current_state_reg[42]  ( .D(AddRoundKeyOutput3[42]), 
        .CK(clk), .Q(PermutationOutput3[26]) );
  DFF_X1 \StateReg3_s_current_state_reg[43]  ( .D(AddRoundKeyOutput3[43]), 
        .CK(clk), .Q(PermutationOutput3[27]) );
  DFF_X1 \StateReg3_s_current_state_reg[44]  ( .D(AddRoundKeyOutput3[44]), 
        .CK(clk), .Q(PermutationOutput3[20]) );
  DFF_X1 \StateReg3_s_current_state_reg[45]  ( .D(AddRoundKeyOutput3[45]), 
        .CK(clk), .Q(PermutationOutput3[21]) );
  DFF_X1 \StateReg3_s_current_state_reg[46]  ( .D(AddRoundKeyOutput3[46]), 
        .CK(clk), .Q(PermutationOutput3[22]) );
  DFF_X1 \StateReg3_s_current_state_reg[47]  ( .D(AddRoundKeyOutput3[47]), 
        .CK(clk), .Q(PermutationOutput3[23]) );
  DFF_X1 \StateReg3_s_current_state_reg[48]  ( .D(AddRoundKeyOutput3[48]), 
        .CK(clk), .Q(PermutationOutput3[4]) );
  DFF_X1 \StateReg3_s_current_state_reg[49]  ( .D(AddRoundKeyOutput3[49]), 
        .CK(clk), .Q(PermutationOutput3[5]) );
  DFF_X1 \StateReg3_s_current_state_reg[50]  ( .D(AddRoundKeyOutput3[50]), 
        .CK(clk), .Q(PermutationOutput3[6]) );
  DFF_X1 \StateReg3_s_current_state_reg[51]  ( .D(AddRoundKeyOutput3[51]), 
        .CK(clk), .Q(PermutationOutput3[7]) );
  DFF_X1 \StateReg3_s_current_state_reg[52]  ( .D(AddRoundKeyOutput3[52]), 
        .CK(clk), .Q(PermutationOutput3[8]) );
  DFF_X1 \StateReg3_s_current_state_reg[53]  ( .D(AddRoundKeyOutput3[53]), 
        .CK(clk), .Q(PermutationOutput3[9]) );
  DFF_X1 \StateReg3_s_current_state_reg[54]  ( .D(AddRoundKeyOutput3[54]), 
        .CK(clk), .Q(PermutationOutput3[10]) );
  DFF_X1 \StateReg3_s_current_state_reg[55]  ( .D(AddRoundKeyOutput3[55]), 
        .CK(clk), .Q(PermutationOutput3[11]) );
  DFF_X1 \StateReg3_s_current_state_reg[56]  ( .D(AddRoundKeyOutput3[56]), 
        .CK(clk), .Q(PermutationOutput3[12]) );
  DFF_X1 \StateReg3_s_current_state_reg[57]  ( .D(AddRoundKeyOutput3[57]), 
        .CK(clk), .Q(PermutationOutput3[13]) );
  DFF_X1 \StateReg3_s_current_state_reg[58]  ( .D(AddRoundKeyOutput3[58]), 
        .CK(clk), .Q(PermutationOutput3[14]) );
  DFF_X1 \StateReg3_s_current_state_reg[59]  ( .D(AddRoundKeyOutput3[59]), 
        .CK(clk), .Q(PermutationOutput3[15]) );
  DFF_X1 \StateReg3_s_current_state_reg[60]  ( .D(AddRoundKeyOutput3[60]), 
        .CK(clk), .Q(PermutationOutput3[0]) );
  DFF_X1 \StateReg3_s_current_state_reg[61]  ( .D(AddRoundKeyOutput3[61]), 
        .CK(clk), .Q(PermutationOutput3[1]) );
  DFF_X1 \StateReg3_s_current_state_reg[62]  ( .D(AddRoundKeyOutput3[62]), 
        .CK(clk), .Q(PermutationOutput3[2]) );
  DFF_X1 \StateReg3_s_current_state_reg[63]  ( .D(AddRoundKeyOutput3[63]), 
        .CK(clk), .Q(PermutationOutput3[3]) );
  NOR2_X1 \SubCellInst3_LFInst_0_LFInst_0_U8  ( .A1(
        \SubCellInst3_LFInst_0_LFInst_0_n11 ), .A2(
        \SubCellInst3_LFInst_0_LFInst_0_n10 ), .ZN(Output[0]) );
  AND2_X1 \SubCellInst3_LFInst_0_LFInst_0_U7  ( .A1(PermutationOutput3[3]), 
        .A2(PermutationOutput3[2]), .ZN(\SubCellInst3_LFInst_0_LFInst_0_n10 )
         );
  NOR2_X1 \SubCellInst3_LFInst_0_LFInst_0_U6  ( .A1(PermutationOutput3[1]), 
        .A2(\SubCellInst3_LFInst_0_LFInst_0_n9 ), .ZN(
        \SubCellInst3_LFInst_0_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst3_LFInst_0_LFInst_0_U5  ( .A1(
        \SubCellInst3_LFInst_0_LFInst_0_n8 ), .A2(
        \SubCellInst3_LFInst_0_LFInst_0_n7 ), .ZN(
        \SubCellInst3_LFInst_0_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst3_LFInst_0_LFInst_0_U4  ( .A1(PermutationOutput3[3]), 
        .A2(PermutationOutput3[2]), .ZN(\SubCellInst3_LFInst_0_LFInst_0_n7 )
         );
  INV_X1 \SubCellInst3_LFInst_0_LFInst_0_U3  ( .A(PermutationOutput3[0]), .ZN(
        \SubCellInst3_LFInst_0_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst3_LFInst_0_LFInst_1_U6  ( .A1(
        \SubCellInst3_LFInst_0_LFInst_1_n6 ), .A2(
        \SubCellInst3_LFInst_0_LFInst_1_n5 ), .ZN(Output[1]) );
  NAND2_X1 \SubCellInst3_LFInst_0_LFInst_1_U5  ( .A1(PermutationOutput3[2]), 
        .A2(PermutationOutput3[0]), .ZN(\SubCellInst3_LFInst_0_LFInst_1_n5 )
         );
  OR2_X1 \SubCellInst3_LFInst_0_LFInst_1_U4  ( .A1(PermutationOutput3[3]), 
        .A2(\SubCellInst3_LFInst_0_LFInst_1_n4 ), .ZN(
        \SubCellInst3_LFInst_0_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst3_LFInst_0_LFInst_1_U3  ( .A1(PermutationOutput3[2]), 
        .A2(PermutationOutput3[0]), .ZN(\SubCellInst3_LFInst_0_LFInst_1_n4 )
         );
  NAND2_X1 \SubCellInst3_LFInst_0_LFInst_2_U8  ( .A1(
        \SubCellInst3_LFInst_0_LFInst_2_n11 ), .A2(
        \SubCellInst3_LFInst_0_LFInst_2_n10 ), .ZN(Output[2]) );
  OR2_X1 \SubCellInst3_LFInst_0_LFInst_2_U7  ( .A1(PermutationOutput3[0]), 
        .A2(PermutationOutput3[3]), .ZN(\SubCellInst3_LFInst_0_LFInst_2_n10 )
         );
  NAND2_X1 \SubCellInst3_LFInst_0_LFInst_2_U6  ( .A1(PermutationOutput3[1]), 
        .A2(\SubCellInst3_LFInst_0_LFInst_2_n9 ), .ZN(
        \SubCellInst3_LFInst_0_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst3_LFInst_0_LFInst_2_U5  ( .A1(
        \SubCellInst3_LFInst_0_LFInst_2_n8 ), .A2(
        \SubCellInst3_LFInst_0_LFInst_2_n7 ), .ZN(
        \SubCellInst3_LFInst_0_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst3_LFInst_0_LFInst_2_U4  ( .A1(PermutationOutput3[0]), 
        .A2(PermutationOutput3[3]), .ZN(\SubCellInst3_LFInst_0_LFInst_2_n7 )
         );
  INV_X1 \SubCellInst3_LFInst_0_LFInst_2_U3  ( .A(PermutationOutput3[2]), .ZN(
        \SubCellInst3_LFInst_0_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst3_LFInst_0_LFInst_3_U6  ( .A1(
        \SubCellInst3_LFInst_0_LFInst_3_n6 ), .A2(
        \SubCellInst3_LFInst_0_LFInst_3_n5 ), .ZN(Output[3]) );
  NOR2_X1 \SubCellInst3_LFInst_0_LFInst_3_U5  ( .A1(PermutationOutput3[3]), 
        .A2(PermutationOutput3[0]), .ZN(\SubCellInst3_LFInst_0_LFInst_3_n5 )
         );
  NOR2_X1 \SubCellInst3_LFInst_0_LFInst_3_U4  ( .A1(PermutationOutput3[1]), 
        .A2(\SubCellInst3_LFInst_0_LFInst_3_n4 ), .ZN(
        \SubCellInst3_LFInst_0_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst3_LFInst_0_LFInst_3_U3  ( .A1(PermutationOutput3[3]), 
        .A2(PermutationOutput3[2]), .ZN(\SubCellInst3_LFInst_0_LFInst_3_n4 )
         );
  NOR2_X1 \SubCellInst3_LFInst_1_LFInst_0_U8  ( .A1(
        \SubCellInst3_LFInst_1_LFInst_0_n11 ), .A2(
        \SubCellInst3_LFInst_1_LFInst_0_n10 ), .ZN(Output[4]) );
  AND2_X1 \SubCellInst3_LFInst_1_LFInst_0_U7  ( .A1(PermutationOutput3[7]), 
        .A2(PermutationOutput3[6]), .ZN(\SubCellInst3_LFInst_1_LFInst_0_n10 )
         );
  NOR2_X1 \SubCellInst3_LFInst_1_LFInst_0_U6  ( .A1(PermutationOutput3[5]), 
        .A2(\SubCellInst3_LFInst_1_LFInst_0_n9 ), .ZN(
        \SubCellInst3_LFInst_1_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst3_LFInst_1_LFInst_0_U5  ( .A1(
        \SubCellInst3_LFInst_1_LFInst_0_n8 ), .A2(
        \SubCellInst3_LFInst_1_LFInst_0_n7 ), .ZN(
        \SubCellInst3_LFInst_1_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst3_LFInst_1_LFInst_0_U4  ( .A1(PermutationOutput3[7]), 
        .A2(PermutationOutput3[6]), .ZN(\SubCellInst3_LFInst_1_LFInst_0_n7 )
         );
  INV_X1 \SubCellInst3_LFInst_1_LFInst_0_U3  ( .A(PermutationOutput3[4]), .ZN(
        \SubCellInst3_LFInst_1_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst3_LFInst_1_LFInst_1_U6  ( .A1(
        \SubCellInst3_LFInst_1_LFInst_1_n6 ), .A2(
        \SubCellInst3_LFInst_1_LFInst_1_n5 ), .ZN(Output[5]) );
  NAND2_X1 \SubCellInst3_LFInst_1_LFInst_1_U5  ( .A1(PermutationOutput3[6]), 
        .A2(PermutationOutput3[4]), .ZN(\SubCellInst3_LFInst_1_LFInst_1_n5 )
         );
  OR2_X1 \SubCellInst3_LFInst_1_LFInst_1_U4  ( .A1(PermutationOutput3[7]), 
        .A2(\SubCellInst3_LFInst_1_LFInst_1_n4 ), .ZN(
        \SubCellInst3_LFInst_1_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst3_LFInst_1_LFInst_1_U3  ( .A1(PermutationOutput3[6]), 
        .A2(PermutationOutput3[4]), .ZN(\SubCellInst3_LFInst_1_LFInst_1_n4 )
         );
  NAND2_X1 \SubCellInst3_LFInst_1_LFInst_2_U8  ( .A1(
        \SubCellInst3_LFInst_1_LFInst_2_n11 ), .A2(
        \SubCellInst3_LFInst_1_LFInst_2_n10 ), .ZN(Output[6]) );
  OR2_X1 \SubCellInst3_LFInst_1_LFInst_2_U7  ( .A1(PermutationOutput3[4]), 
        .A2(PermutationOutput3[7]), .ZN(\SubCellInst3_LFInst_1_LFInst_2_n10 )
         );
  NAND2_X1 \SubCellInst3_LFInst_1_LFInst_2_U6  ( .A1(PermutationOutput3[5]), 
        .A2(\SubCellInst3_LFInst_1_LFInst_2_n9 ), .ZN(
        \SubCellInst3_LFInst_1_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst3_LFInst_1_LFInst_2_U5  ( .A1(
        \SubCellInst3_LFInst_1_LFInst_2_n8 ), .A2(
        \SubCellInst3_LFInst_1_LFInst_2_n7 ), .ZN(
        \SubCellInst3_LFInst_1_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst3_LFInst_1_LFInst_2_U4  ( .A1(PermutationOutput3[4]), 
        .A2(PermutationOutput3[7]), .ZN(\SubCellInst3_LFInst_1_LFInst_2_n7 )
         );
  INV_X1 \SubCellInst3_LFInst_1_LFInst_2_U3  ( .A(PermutationOutput3[6]), .ZN(
        \SubCellInst3_LFInst_1_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst3_LFInst_1_LFInst_3_U6  ( .A1(
        \SubCellInst3_LFInst_1_LFInst_3_n6 ), .A2(
        \SubCellInst3_LFInst_1_LFInst_3_n5 ), .ZN(Output[7]) );
  NOR2_X1 \SubCellInst3_LFInst_1_LFInst_3_U5  ( .A1(PermutationOutput3[7]), 
        .A2(PermutationOutput3[4]), .ZN(\SubCellInst3_LFInst_1_LFInst_3_n5 )
         );
  NOR2_X1 \SubCellInst3_LFInst_1_LFInst_3_U4  ( .A1(PermutationOutput3[5]), 
        .A2(\SubCellInst3_LFInst_1_LFInst_3_n4 ), .ZN(
        \SubCellInst3_LFInst_1_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst3_LFInst_1_LFInst_3_U3  ( .A1(PermutationOutput3[7]), 
        .A2(PermutationOutput3[6]), .ZN(\SubCellInst3_LFInst_1_LFInst_3_n4 )
         );
  NOR2_X1 \SubCellInst3_LFInst_2_LFInst_0_U8  ( .A1(
        \SubCellInst3_LFInst_2_LFInst_0_n11 ), .A2(
        \SubCellInst3_LFInst_2_LFInst_0_n10 ), .ZN(Output[8]) );
  AND2_X1 \SubCellInst3_LFInst_2_LFInst_0_U7  ( .A1(PermutationOutput3[11]), 
        .A2(PermutationOutput3[10]), .ZN(\SubCellInst3_LFInst_2_LFInst_0_n10 )
         );
  NOR2_X1 \SubCellInst3_LFInst_2_LFInst_0_U6  ( .A1(PermutationOutput3[9]), 
        .A2(\SubCellInst3_LFInst_2_LFInst_0_n9 ), .ZN(
        \SubCellInst3_LFInst_2_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst3_LFInst_2_LFInst_0_U5  ( .A1(
        \SubCellInst3_LFInst_2_LFInst_0_n8 ), .A2(
        \SubCellInst3_LFInst_2_LFInst_0_n7 ), .ZN(
        \SubCellInst3_LFInst_2_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst3_LFInst_2_LFInst_0_U4  ( .A1(PermutationOutput3[11]), 
        .A2(PermutationOutput3[10]), .ZN(\SubCellInst3_LFInst_2_LFInst_0_n7 )
         );
  INV_X1 \SubCellInst3_LFInst_2_LFInst_0_U3  ( .A(PermutationOutput3[8]), .ZN(
        \SubCellInst3_LFInst_2_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst3_LFInst_2_LFInst_1_U6  ( .A1(
        \SubCellInst3_LFInst_2_LFInst_1_n6 ), .A2(
        \SubCellInst3_LFInst_2_LFInst_1_n5 ), .ZN(Output[9]) );
  NAND2_X1 \SubCellInst3_LFInst_2_LFInst_1_U5  ( .A1(PermutationOutput3[10]), 
        .A2(PermutationOutput3[8]), .ZN(\SubCellInst3_LFInst_2_LFInst_1_n5 )
         );
  OR2_X1 \SubCellInst3_LFInst_2_LFInst_1_U4  ( .A1(PermutationOutput3[11]), 
        .A2(\SubCellInst3_LFInst_2_LFInst_1_n4 ), .ZN(
        \SubCellInst3_LFInst_2_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst3_LFInst_2_LFInst_1_U3  ( .A1(PermutationOutput3[10]), 
        .A2(PermutationOutput3[8]), .ZN(\SubCellInst3_LFInst_2_LFInst_1_n4 )
         );
  NAND2_X1 \SubCellInst3_LFInst_2_LFInst_2_U8  ( .A1(
        \SubCellInst3_LFInst_2_LFInst_2_n11 ), .A2(
        \SubCellInst3_LFInst_2_LFInst_2_n10 ), .ZN(Output[10]) );
  OR2_X1 \SubCellInst3_LFInst_2_LFInst_2_U7  ( .A1(PermutationOutput3[8]), 
        .A2(PermutationOutput3[11]), .ZN(\SubCellInst3_LFInst_2_LFInst_2_n10 )
         );
  NAND2_X1 \SubCellInst3_LFInst_2_LFInst_2_U6  ( .A1(PermutationOutput3[9]), 
        .A2(\SubCellInst3_LFInst_2_LFInst_2_n9 ), .ZN(
        \SubCellInst3_LFInst_2_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst3_LFInst_2_LFInst_2_U5  ( .A1(
        \SubCellInst3_LFInst_2_LFInst_2_n8 ), .A2(
        \SubCellInst3_LFInst_2_LFInst_2_n7 ), .ZN(
        \SubCellInst3_LFInst_2_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst3_LFInst_2_LFInst_2_U4  ( .A1(PermutationOutput3[8]), 
        .A2(PermutationOutput3[11]), .ZN(\SubCellInst3_LFInst_2_LFInst_2_n7 )
         );
  INV_X1 \SubCellInst3_LFInst_2_LFInst_2_U3  ( .A(PermutationOutput3[10]), 
        .ZN(\SubCellInst3_LFInst_2_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst3_LFInst_2_LFInst_3_U6  ( .A1(
        \SubCellInst3_LFInst_2_LFInst_3_n6 ), .A2(
        \SubCellInst3_LFInst_2_LFInst_3_n5 ), .ZN(Output[11]) );
  NOR2_X1 \SubCellInst3_LFInst_2_LFInst_3_U5  ( .A1(PermutationOutput3[11]), 
        .A2(PermutationOutput3[8]), .ZN(\SubCellInst3_LFInst_2_LFInst_3_n5 )
         );
  NOR2_X1 \SubCellInst3_LFInst_2_LFInst_3_U4  ( .A1(PermutationOutput3[9]), 
        .A2(\SubCellInst3_LFInst_2_LFInst_3_n4 ), .ZN(
        \SubCellInst3_LFInst_2_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst3_LFInst_2_LFInst_3_U3  ( .A1(PermutationOutput3[11]), 
        .A2(PermutationOutput3[10]), .ZN(\SubCellInst3_LFInst_2_LFInst_3_n4 )
         );
  NOR2_X1 \SubCellInst3_LFInst_3_LFInst_0_U8  ( .A1(
        \SubCellInst3_LFInst_3_LFInst_0_n11 ), .A2(
        \SubCellInst3_LFInst_3_LFInst_0_n10 ), .ZN(Output[12]) );
  AND2_X1 \SubCellInst3_LFInst_3_LFInst_0_U7  ( .A1(PermutationOutput3[15]), 
        .A2(PermutationOutput3[14]), .ZN(\SubCellInst3_LFInst_3_LFInst_0_n10 )
         );
  NOR2_X1 \SubCellInst3_LFInst_3_LFInst_0_U6  ( .A1(PermutationOutput3[13]), 
        .A2(\SubCellInst3_LFInst_3_LFInst_0_n9 ), .ZN(
        \SubCellInst3_LFInst_3_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst3_LFInst_3_LFInst_0_U5  ( .A1(
        \SubCellInst3_LFInst_3_LFInst_0_n8 ), .A2(
        \SubCellInst3_LFInst_3_LFInst_0_n7 ), .ZN(
        \SubCellInst3_LFInst_3_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst3_LFInst_3_LFInst_0_U4  ( .A1(PermutationOutput3[15]), 
        .A2(PermutationOutput3[14]), .ZN(\SubCellInst3_LFInst_3_LFInst_0_n7 )
         );
  INV_X1 \SubCellInst3_LFInst_3_LFInst_0_U3  ( .A(PermutationOutput3[12]), 
        .ZN(\SubCellInst3_LFInst_3_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst3_LFInst_3_LFInst_1_U6  ( .A1(
        \SubCellInst3_LFInst_3_LFInst_1_n6 ), .A2(
        \SubCellInst3_LFInst_3_LFInst_1_n5 ), .ZN(Output[13]) );
  NAND2_X1 \SubCellInst3_LFInst_3_LFInst_1_U5  ( .A1(PermutationOutput3[14]), 
        .A2(PermutationOutput3[12]), .ZN(\SubCellInst3_LFInst_3_LFInst_1_n5 )
         );
  OR2_X1 \SubCellInst3_LFInst_3_LFInst_1_U4  ( .A1(PermutationOutput3[15]), 
        .A2(\SubCellInst3_LFInst_3_LFInst_1_n4 ), .ZN(
        \SubCellInst3_LFInst_3_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst3_LFInst_3_LFInst_1_U3  ( .A1(PermutationOutput3[14]), 
        .A2(PermutationOutput3[12]), .ZN(\SubCellInst3_LFInst_3_LFInst_1_n4 )
         );
  NAND2_X1 \SubCellInst3_LFInst_3_LFInst_2_U8  ( .A1(
        \SubCellInst3_LFInst_3_LFInst_2_n11 ), .A2(
        \SubCellInst3_LFInst_3_LFInst_2_n10 ), .ZN(Output[14]) );
  OR2_X1 \SubCellInst3_LFInst_3_LFInst_2_U7  ( .A1(PermutationOutput3[12]), 
        .A2(PermutationOutput3[15]), .ZN(\SubCellInst3_LFInst_3_LFInst_2_n10 )
         );
  NAND2_X1 \SubCellInst3_LFInst_3_LFInst_2_U6  ( .A1(PermutationOutput3[13]), 
        .A2(\SubCellInst3_LFInst_3_LFInst_2_n9 ), .ZN(
        \SubCellInst3_LFInst_3_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst3_LFInst_3_LFInst_2_U5  ( .A1(
        \SubCellInst3_LFInst_3_LFInst_2_n8 ), .A2(
        \SubCellInst3_LFInst_3_LFInst_2_n7 ), .ZN(
        \SubCellInst3_LFInst_3_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst3_LFInst_3_LFInst_2_U4  ( .A1(PermutationOutput3[12]), 
        .A2(PermutationOutput3[15]), .ZN(\SubCellInst3_LFInst_3_LFInst_2_n7 )
         );
  INV_X1 \SubCellInst3_LFInst_3_LFInst_2_U3  ( .A(PermutationOutput3[14]), 
        .ZN(\SubCellInst3_LFInst_3_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst3_LFInst_3_LFInst_3_U6  ( .A1(
        \SubCellInst3_LFInst_3_LFInst_3_n6 ), .A2(
        \SubCellInst3_LFInst_3_LFInst_3_n5 ), .ZN(Output[15]) );
  NOR2_X1 \SubCellInst3_LFInst_3_LFInst_3_U5  ( .A1(PermutationOutput3[15]), 
        .A2(PermutationOutput3[12]), .ZN(\SubCellInst3_LFInst_3_LFInst_3_n5 )
         );
  NOR2_X1 \SubCellInst3_LFInst_3_LFInst_3_U4  ( .A1(PermutationOutput3[13]), 
        .A2(\SubCellInst3_LFInst_3_LFInst_3_n4 ), .ZN(
        \SubCellInst3_LFInst_3_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst3_LFInst_3_LFInst_3_U3  ( .A1(PermutationOutput3[15]), 
        .A2(PermutationOutput3[14]), .ZN(\SubCellInst3_LFInst_3_LFInst_3_n4 )
         );
  NOR2_X1 \SubCellInst3_LFInst_4_LFInst_0_U8  ( .A1(
        \SubCellInst3_LFInst_4_LFInst_0_n11 ), .A2(
        \SubCellInst3_LFInst_4_LFInst_0_n10 ), .ZN(Output[16]) );
  AND2_X1 \SubCellInst3_LFInst_4_LFInst_0_U7  ( .A1(PermutationOutput3[19]), 
        .A2(PermutationOutput3[18]), .ZN(\SubCellInst3_LFInst_4_LFInst_0_n10 )
         );
  NOR2_X1 \SubCellInst3_LFInst_4_LFInst_0_U6  ( .A1(PermutationOutput3[17]), 
        .A2(\SubCellInst3_LFInst_4_LFInst_0_n9 ), .ZN(
        \SubCellInst3_LFInst_4_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst3_LFInst_4_LFInst_0_U5  ( .A1(
        \SubCellInst3_LFInst_4_LFInst_0_n8 ), .A2(
        \SubCellInst3_LFInst_4_LFInst_0_n7 ), .ZN(
        \SubCellInst3_LFInst_4_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst3_LFInst_4_LFInst_0_U4  ( .A1(PermutationOutput3[19]), 
        .A2(PermutationOutput3[18]), .ZN(\SubCellInst3_LFInst_4_LFInst_0_n7 )
         );
  INV_X1 \SubCellInst3_LFInst_4_LFInst_0_U3  ( .A(PermutationOutput3[16]), 
        .ZN(\SubCellInst3_LFInst_4_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst3_LFInst_4_LFInst_1_U6  ( .A1(
        \SubCellInst3_LFInst_4_LFInst_1_n6 ), .A2(
        \SubCellInst3_LFInst_4_LFInst_1_n5 ), .ZN(Output[17]) );
  NAND2_X1 \SubCellInst3_LFInst_4_LFInst_1_U5  ( .A1(PermutationOutput3[18]), 
        .A2(PermutationOutput3[16]), .ZN(\SubCellInst3_LFInst_4_LFInst_1_n5 )
         );
  OR2_X1 \SubCellInst3_LFInst_4_LFInst_1_U4  ( .A1(PermutationOutput3[19]), 
        .A2(\SubCellInst3_LFInst_4_LFInst_1_n4 ), .ZN(
        \SubCellInst3_LFInst_4_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst3_LFInst_4_LFInst_1_U3  ( .A1(PermutationOutput3[18]), 
        .A2(PermutationOutput3[16]), .ZN(\SubCellInst3_LFInst_4_LFInst_1_n4 )
         );
  NAND2_X1 \SubCellInst3_LFInst_4_LFInst_2_U8  ( .A1(
        \SubCellInst3_LFInst_4_LFInst_2_n11 ), .A2(
        \SubCellInst3_LFInst_4_LFInst_2_n10 ), .ZN(Output[18]) );
  OR2_X1 \SubCellInst3_LFInst_4_LFInst_2_U7  ( .A1(PermutationOutput3[16]), 
        .A2(PermutationOutput3[19]), .ZN(\SubCellInst3_LFInst_4_LFInst_2_n10 )
         );
  NAND2_X1 \SubCellInst3_LFInst_4_LFInst_2_U6  ( .A1(PermutationOutput3[17]), 
        .A2(\SubCellInst3_LFInst_4_LFInst_2_n9 ), .ZN(
        \SubCellInst3_LFInst_4_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst3_LFInst_4_LFInst_2_U5  ( .A1(
        \SubCellInst3_LFInst_4_LFInst_2_n8 ), .A2(
        \SubCellInst3_LFInst_4_LFInst_2_n7 ), .ZN(
        \SubCellInst3_LFInst_4_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst3_LFInst_4_LFInst_2_U4  ( .A1(PermutationOutput3[16]), 
        .A2(PermutationOutput3[19]), .ZN(\SubCellInst3_LFInst_4_LFInst_2_n7 )
         );
  INV_X1 \SubCellInst3_LFInst_4_LFInst_2_U3  ( .A(PermutationOutput3[18]), 
        .ZN(\SubCellInst3_LFInst_4_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst3_LFInst_4_LFInst_3_U6  ( .A1(
        \SubCellInst3_LFInst_4_LFInst_3_n6 ), .A2(
        \SubCellInst3_LFInst_4_LFInst_3_n5 ), .ZN(Output[19]) );
  NOR2_X1 \SubCellInst3_LFInst_4_LFInst_3_U5  ( .A1(PermutationOutput3[19]), 
        .A2(PermutationOutput3[16]), .ZN(\SubCellInst3_LFInst_4_LFInst_3_n5 )
         );
  NOR2_X1 \SubCellInst3_LFInst_4_LFInst_3_U4  ( .A1(PermutationOutput3[17]), 
        .A2(\SubCellInst3_LFInst_4_LFInst_3_n4 ), .ZN(
        \SubCellInst3_LFInst_4_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst3_LFInst_4_LFInst_3_U3  ( .A1(PermutationOutput3[19]), 
        .A2(PermutationOutput3[18]), .ZN(\SubCellInst3_LFInst_4_LFInst_3_n4 )
         );
  NOR2_X1 \SubCellInst3_LFInst_5_LFInst_0_U8  ( .A1(
        \SubCellInst3_LFInst_5_LFInst_0_n11 ), .A2(
        \SubCellInst3_LFInst_5_LFInst_0_n10 ), .ZN(Output[20]) );
  AND2_X1 \SubCellInst3_LFInst_5_LFInst_0_U7  ( .A1(PermutationOutput3[23]), 
        .A2(PermutationOutput3[22]), .ZN(\SubCellInst3_LFInst_5_LFInst_0_n10 )
         );
  NOR2_X1 \SubCellInst3_LFInst_5_LFInst_0_U6  ( .A1(PermutationOutput3[21]), 
        .A2(\SubCellInst3_LFInst_5_LFInst_0_n9 ), .ZN(
        \SubCellInst3_LFInst_5_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst3_LFInst_5_LFInst_0_U5  ( .A1(
        \SubCellInst3_LFInst_5_LFInst_0_n8 ), .A2(
        \SubCellInst3_LFInst_5_LFInst_0_n7 ), .ZN(
        \SubCellInst3_LFInst_5_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst3_LFInst_5_LFInst_0_U4  ( .A1(PermutationOutput3[23]), 
        .A2(PermutationOutput3[22]), .ZN(\SubCellInst3_LFInst_5_LFInst_0_n7 )
         );
  INV_X1 \SubCellInst3_LFInst_5_LFInst_0_U3  ( .A(PermutationOutput3[20]), 
        .ZN(\SubCellInst3_LFInst_5_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst3_LFInst_5_LFInst_1_U6  ( .A1(
        \SubCellInst3_LFInst_5_LFInst_1_n6 ), .A2(
        \SubCellInst3_LFInst_5_LFInst_1_n5 ), .ZN(Output[21]) );
  NAND2_X1 \SubCellInst3_LFInst_5_LFInst_1_U5  ( .A1(PermutationOutput3[22]), 
        .A2(PermutationOutput3[20]), .ZN(\SubCellInst3_LFInst_5_LFInst_1_n5 )
         );
  OR2_X1 \SubCellInst3_LFInst_5_LFInst_1_U4  ( .A1(PermutationOutput3[23]), 
        .A2(\SubCellInst3_LFInst_5_LFInst_1_n4 ), .ZN(
        \SubCellInst3_LFInst_5_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst3_LFInst_5_LFInst_1_U3  ( .A1(PermutationOutput3[22]), 
        .A2(PermutationOutput3[20]), .ZN(\SubCellInst3_LFInst_5_LFInst_1_n4 )
         );
  NAND2_X1 \SubCellInst3_LFInst_5_LFInst_2_U8  ( .A1(
        \SubCellInst3_LFInst_5_LFInst_2_n11 ), .A2(
        \SubCellInst3_LFInst_5_LFInst_2_n10 ), .ZN(Output[22]) );
  OR2_X1 \SubCellInst3_LFInst_5_LFInst_2_U7  ( .A1(PermutationOutput3[20]), 
        .A2(PermutationOutput3[23]), .ZN(\SubCellInst3_LFInst_5_LFInst_2_n10 )
         );
  NAND2_X1 \SubCellInst3_LFInst_5_LFInst_2_U6  ( .A1(PermutationOutput3[21]), 
        .A2(\SubCellInst3_LFInst_5_LFInst_2_n9 ), .ZN(
        \SubCellInst3_LFInst_5_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst3_LFInst_5_LFInst_2_U5  ( .A1(
        \SubCellInst3_LFInst_5_LFInst_2_n8 ), .A2(
        \SubCellInst3_LFInst_5_LFInst_2_n7 ), .ZN(
        \SubCellInst3_LFInst_5_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst3_LFInst_5_LFInst_2_U4  ( .A1(PermutationOutput3[20]), 
        .A2(PermutationOutput3[23]), .ZN(\SubCellInst3_LFInst_5_LFInst_2_n7 )
         );
  INV_X1 \SubCellInst3_LFInst_5_LFInst_2_U3  ( .A(PermutationOutput3[22]), 
        .ZN(\SubCellInst3_LFInst_5_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst3_LFInst_5_LFInst_3_U6  ( .A1(
        \SubCellInst3_LFInst_5_LFInst_3_n6 ), .A2(
        \SubCellInst3_LFInst_5_LFInst_3_n5 ), .ZN(Output[23]) );
  NOR2_X1 \SubCellInst3_LFInst_5_LFInst_3_U5  ( .A1(PermutationOutput3[23]), 
        .A2(PermutationOutput3[20]), .ZN(\SubCellInst3_LFInst_5_LFInst_3_n5 )
         );
  NOR2_X1 \SubCellInst3_LFInst_5_LFInst_3_U4  ( .A1(PermutationOutput3[21]), 
        .A2(\SubCellInst3_LFInst_5_LFInst_3_n4 ), .ZN(
        \SubCellInst3_LFInst_5_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst3_LFInst_5_LFInst_3_U3  ( .A1(PermutationOutput3[23]), 
        .A2(PermutationOutput3[22]), .ZN(\SubCellInst3_LFInst_5_LFInst_3_n4 )
         );
  NOR2_X1 \SubCellInst3_LFInst_6_LFInst_0_U8  ( .A1(
        \SubCellInst3_LFInst_6_LFInst_0_n11 ), .A2(
        \SubCellInst3_LFInst_6_LFInst_0_n10 ), .ZN(Output[24]) );
  AND2_X1 \SubCellInst3_LFInst_6_LFInst_0_U7  ( .A1(PermutationOutput3[27]), 
        .A2(PermutationOutput3[26]), .ZN(\SubCellInst3_LFInst_6_LFInst_0_n10 )
         );
  NOR2_X1 \SubCellInst3_LFInst_6_LFInst_0_U6  ( .A1(PermutationOutput3[25]), 
        .A2(\SubCellInst3_LFInst_6_LFInst_0_n9 ), .ZN(
        \SubCellInst3_LFInst_6_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst3_LFInst_6_LFInst_0_U5  ( .A1(
        \SubCellInst3_LFInst_6_LFInst_0_n8 ), .A2(
        \SubCellInst3_LFInst_6_LFInst_0_n7 ), .ZN(
        \SubCellInst3_LFInst_6_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst3_LFInst_6_LFInst_0_U4  ( .A1(PermutationOutput3[27]), 
        .A2(PermutationOutput3[26]), .ZN(\SubCellInst3_LFInst_6_LFInst_0_n7 )
         );
  INV_X1 \SubCellInst3_LFInst_6_LFInst_0_U3  ( .A(PermutationOutput3[24]), 
        .ZN(\SubCellInst3_LFInst_6_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst3_LFInst_6_LFInst_1_U6  ( .A1(
        \SubCellInst3_LFInst_6_LFInst_1_n6 ), .A2(
        \SubCellInst3_LFInst_6_LFInst_1_n5 ), .ZN(Output[25]) );
  NAND2_X1 \SubCellInst3_LFInst_6_LFInst_1_U5  ( .A1(PermutationOutput3[26]), 
        .A2(PermutationOutput3[24]), .ZN(\SubCellInst3_LFInst_6_LFInst_1_n5 )
         );
  OR2_X1 \SubCellInst3_LFInst_6_LFInst_1_U4  ( .A1(PermutationOutput3[27]), 
        .A2(\SubCellInst3_LFInst_6_LFInst_1_n4 ), .ZN(
        \SubCellInst3_LFInst_6_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst3_LFInst_6_LFInst_1_U3  ( .A1(PermutationOutput3[26]), 
        .A2(PermutationOutput3[24]), .ZN(\SubCellInst3_LFInst_6_LFInst_1_n4 )
         );
  NAND2_X1 \SubCellInst3_LFInst_6_LFInst_2_U8  ( .A1(
        \SubCellInst3_LFInst_6_LFInst_2_n11 ), .A2(
        \SubCellInst3_LFInst_6_LFInst_2_n10 ), .ZN(Output[26]) );
  OR2_X1 \SubCellInst3_LFInst_6_LFInst_2_U7  ( .A1(PermutationOutput3[24]), 
        .A2(PermutationOutput3[27]), .ZN(\SubCellInst3_LFInst_6_LFInst_2_n10 )
         );
  NAND2_X1 \SubCellInst3_LFInst_6_LFInst_2_U6  ( .A1(PermutationOutput3[25]), 
        .A2(\SubCellInst3_LFInst_6_LFInst_2_n9 ), .ZN(
        \SubCellInst3_LFInst_6_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst3_LFInst_6_LFInst_2_U5  ( .A1(
        \SubCellInst3_LFInst_6_LFInst_2_n8 ), .A2(
        \SubCellInst3_LFInst_6_LFInst_2_n7 ), .ZN(
        \SubCellInst3_LFInst_6_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst3_LFInst_6_LFInst_2_U4  ( .A1(PermutationOutput3[24]), 
        .A2(PermutationOutput3[27]), .ZN(\SubCellInst3_LFInst_6_LFInst_2_n7 )
         );
  INV_X1 \SubCellInst3_LFInst_6_LFInst_2_U3  ( .A(PermutationOutput3[26]), 
        .ZN(\SubCellInst3_LFInst_6_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst3_LFInst_6_LFInst_3_U6  ( .A1(
        \SubCellInst3_LFInst_6_LFInst_3_n6 ), .A2(
        \SubCellInst3_LFInst_6_LFInst_3_n5 ), .ZN(Output[27]) );
  NOR2_X1 \SubCellInst3_LFInst_6_LFInst_3_U5  ( .A1(PermutationOutput3[27]), 
        .A2(PermutationOutput3[24]), .ZN(\SubCellInst3_LFInst_6_LFInst_3_n5 )
         );
  NOR2_X1 \SubCellInst3_LFInst_6_LFInst_3_U4  ( .A1(PermutationOutput3[25]), 
        .A2(\SubCellInst3_LFInst_6_LFInst_3_n4 ), .ZN(
        \SubCellInst3_LFInst_6_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst3_LFInst_6_LFInst_3_U3  ( .A1(PermutationOutput3[27]), 
        .A2(PermutationOutput3[26]), .ZN(\SubCellInst3_LFInst_6_LFInst_3_n4 )
         );
  NOR2_X1 \SubCellInst3_LFInst_7_LFInst_0_U8  ( .A1(
        \SubCellInst3_LFInst_7_LFInst_0_n11 ), .A2(
        \SubCellInst3_LFInst_7_LFInst_0_n10 ), .ZN(Output[28]) );
  AND2_X1 \SubCellInst3_LFInst_7_LFInst_0_U7  ( .A1(PermutationOutput3[31]), 
        .A2(PermutationOutput3[30]), .ZN(\SubCellInst3_LFInst_7_LFInst_0_n10 )
         );
  NOR2_X1 \SubCellInst3_LFInst_7_LFInst_0_U6  ( .A1(PermutationOutput3[29]), 
        .A2(\SubCellInst3_LFInst_7_LFInst_0_n9 ), .ZN(
        \SubCellInst3_LFInst_7_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst3_LFInst_7_LFInst_0_U5  ( .A1(
        \SubCellInst3_LFInst_7_LFInst_0_n8 ), .A2(
        \SubCellInst3_LFInst_7_LFInst_0_n7 ), .ZN(
        \SubCellInst3_LFInst_7_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst3_LFInst_7_LFInst_0_U4  ( .A1(PermutationOutput3[31]), 
        .A2(PermutationOutput3[30]), .ZN(\SubCellInst3_LFInst_7_LFInst_0_n7 )
         );
  INV_X1 \SubCellInst3_LFInst_7_LFInst_0_U3  ( .A(PermutationOutput3[28]), 
        .ZN(\SubCellInst3_LFInst_7_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst3_LFInst_7_LFInst_1_U6  ( .A1(
        \SubCellInst3_LFInst_7_LFInst_1_n6 ), .A2(
        \SubCellInst3_LFInst_7_LFInst_1_n5 ), .ZN(Output[29]) );
  NAND2_X1 \SubCellInst3_LFInst_7_LFInst_1_U5  ( .A1(PermutationOutput3[30]), 
        .A2(PermutationOutput3[28]), .ZN(\SubCellInst3_LFInst_7_LFInst_1_n5 )
         );
  OR2_X1 \SubCellInst3_LFInst_7_LFInst_1_U4  ( .A1(PermutationOutput3[31]), 
        .A2(\SubCellInst3_LFInst_7_LFInst_1_n4 ), .ZN(
        \SubCellInst3_LFInst_7_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst3_LFInst_7_LFInst_1_U3  ( .A1(PermutationOutput3[30]), 
        .A2(PermutationOutput3[28]), .ZN(\SubCellInst3_LFInst_7_LFInst_1_n4 )
         );
  NAND2_X1 \SubCellInst3_LFInst_7_LFInst_2_U8  ( .A1(
        \SubCellInst3_LFInst_7_LFInst_2_n11 ), .A2(
        \SubCellInst3_LFInst_7_LFInst_2_n10 ), .ZN(Output[30]) );
  OR2_X1 \SubCellInst3_LFInst_7_LFInst_2_U7  ( .A1(PermutationOutput3[28]), 
        .A2(PermutationOutput3[31]), .ZN(\SubCellInst3_LFInst_7_LFInst_2_n10 )
         );
  NAND2_X1 \SubCellInst3_LFInst_7_LFInst_2_U6  ( .A1(PermutationOutput3[29]), 
        .A2(\SubCellInst3_LFInst_7_LFInst_2_n9 ), .ZN(
        \SubCellInst3_LFInst_7_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst3_LFInst_7_LFInst_2_U5  ( .A1(
        \SubCellInst3_LFInst_7_LFInst_2_n8 ), .A2(
        \SubCellInst3_LFInst_7_LFInst_2_n7 ), .ZN(
        \SubCellInst3_LFInst_7_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst3_LFInst_7_LFInst_2_U4  ( .A1(PermutationOutput3[28]), 
        .A2(PermutationOutput3[31]), .ZN(\SubCellInst3_LFInst_7_LFInst_2_n7 )
         );
  INV_X1 \SubCellInst3_LFInst_7_LFInst_2_U3  ( .A(PermutationOutput3[30]), 
        .ZN(\SubCellInst3_LFInst_7_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst3_LFInst_7_LFInst_3_U6  ( .A1(
        \SubCellInst3_LFInst_7_LFInst_3_n6 ), .A2(
        \SubCellInst3_LFInst_7_LFInst_3_n5 ), .ZN(Output[31]) );
  NOR2_X1 \SubCellInst3_LFInst_7_LFInst_3_U5  ( .A1(PermutationOutput3[31]), 
        .A2(PermutationOutput3[28]), .ZN(\SubCellInst3_LFInst_7_LFInst_3_n5 )
         );
  NOR2_X1 \SubCellInst3_LFInst_7_LFInst_3_U4  ( .A1(PermutationOutput3[29]), 
        .A2(\SubCellInst3_LFInst_7_LFInst_3_n4 ), .ZN(
        \SubCellInst3_LFInst_7_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst3_LFInst_7_LFInst_3_U3  ( .A1(PermutationOutput3[31]), 
        .A2(PermutationOutput3[30]), .ZN(\SubCellInst3_LFInst_7_LFInst_3_n4 )
         );
  NOR2_X1 \SubCellInst3_LFInst_8_LFInst_0_U8  ( .A1(
        \SubCellInst3_LFInst_8_LFInst_0_n11 ), .A2(
        \SubCellInst3_LFInst_8_LFInst_0_n10 ), .ZN(Output[32]) );
  AND2_X1 \SubCellInst3_LFInst_8_LFInst_0_U7  ( .A1(PermutationOutput3[35]), 
        .A2(PermutationOutput3[34]), .ZN(\SubCellInst3_LFInst_8_LFInst_0_n10 )
         );
  NOR2_X1 \SubCellInst3_LFInst_8_LFInst_0_U6  ( .A1(PermutationOutput3[33]), 
        .A2(\SubCellInst3_LFInst_8_LFInst_0_n9 ), .ZN(
        \SubCellInst3_LFInst_8_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst3_LFInst_8_LFInst_0_U5  ( .A1(
        \SubCellInst3_LFInst_8_LFInst_0_n8 ), .A2(
        \SubCellInst3_LFInst_8_LFInst_0_n7 ), .ZN(
        \SubCellInst3_LFInst_8_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst3_LFInst_8_LFInst_0_U4  ( .A1(PermutationOutput3[35]), 
        .A2(PermutationOutput3[34]), .ZN(\SubCellInst3_LFInst_8_LFInst_0_n7 )
         );
  INV_X1 \SubCellInst3_LFInst_8_LFInst_0_U3  ( .A(PermutationOutput3[32]), 
        .ZN(\SubCellInst3_LFInst_8_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst3_LFInst_8_LFInst_1_U6  ( .A1(
        \SubCellInst3_LFInst_8_LFInst_1_n6 ), .A2(
        \SubCellInst3_LFInst_8_LFInst_1_n5 ), .ZN(Output[33]) );
  NAND2_X1 \SubCellInst3_LFInst_8_LFInst_1_U5  ( .A1(PermutationOutput3[34]), 
        .A2(PermutationOutput3[32]), .ZN(\SubCellInst3_LFInst_8_LFInst_1_n5 )
         );
  OR2_X1 \SubCellInst3_LFInst_8_LFInst_1_U4  ( .A1(PermutationOutput3[35]), 
        .A2(\SubCellInst3_LFInst_8_LFInst_1_n4 ), .ZN(
        \SubCellInst3_LFInst_8_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst3_LFInst_8_LFInst_1_U3  ( .A1(PermutationOutput3[34]), 
        .A2(PermutationOutput3[32]), .ZN(\SubCellInst3_LFInst_8_LFInst_1_n4 )
         );
  NAND2_X1 \SubCellInst3_LFInst_8_LFInst_2_U8  ( .A1(
        \SubCellInst3_LFInst_8_LFInst_2_n11 ), .A2(
        \SubCellInst3_LFInst_8_LFInst_2_n10 ), .ZN(Output[34]) );
  OR2_X1 \SubCellInst3_LFInst_8_LFInst_2_U7  ( .A1(PermutationOutput3[32]), 
        .A2(PermutationOutput3[35]), .ZN(\SubCellInst3_LFInst_8_LFInst_2_n10 )
         );
  NAND2_X1 \SubCellInst3_LFInst_8_LFInst_2_U6  ( .A1(PermutationOutput3[33]), 
        .A2(\SubCellInst3_LFInst_8_LFInst_2_n9 ), .ZN(
        \SubCellInst3_LFInst_8_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst3_LFInst_8_LFInst_2_U5  ( .A1(
        \SubCellInst3_LFInst_8_LFInst_2_n8 ), .A2(
        \SubCellInst3_LFInst_8_LFInst_2_n7 ), .ZN(
        \SubCellInst3_LFInst_8_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst3_LFInst_8_LFInst_2_U4  ( .A1(PermutationOutput3[32]), 
        .A2(PermutationOutput3[35]), .ZN(\SubCellInst3_LFInst_8_LFInst_2_n7 )
         );
  INV_X1 \SubCellInst3_LFInst_8_LFInst_2_U3  ( .A(PermutationOutput3[34]), 
        .ZN(\SubCellInst3_LFInst_8_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst3_LFInst_8_LFInst_3_U6  ( .A1(
        \SubCellInst3_LFInst_8_LFInst_3_n6 ), .A2(
        \SubCellInst3_LFInst_8_LFInst_3_n5 ), .ZN(Output[35]) );
  NOR2_X1 \SubCellInst3_LFInst_8_LFInst_3_U5  ( .A1(PermutationOutput3[35]), 
        .A2(PermutationOutput3[32]), .ZN(\SubCellInst3_LFInst_8_LFInst_3_n5 )
         );
  NOR2_X1 \SubCellInst3_LFInst_8_LFInst_3_U4  ( .A1(PermutationOutput3[33]), 
        .A2(\SubCellInst3_LFInst_8_LFInst_3_n4 ), .ZN(
        \SubCellInst3_LFInst_8_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst3_LFInst_8_LFInst_3_U3  ( .A1(PermutationOutput3[35]), 
        .A2(PermutationOutput3[34]), .ZN(\SubCellInst3_LFInst_8_LFInst_3_n4 )
         );
  NOR2_X1 \SubCellInst3_LFInst_9_LFInst_0_U8  ( .A1(
        \SubCellInst3_LFInst_9_LFInst_0_n11 ), .A2(
        \SubCellInst3_LFInst_9_LFInst_0_n10 ), .ZN(Output[36]) );
  AND2_X1 \SubCellInst3_LFInst_9_LFInst_0_U7  ( .A1(PermutationOutput3[39]), 
        .A2(PermutationOutput3[38]), .ZN(\SubCellInst3_LFInst_9_LFInst_0_n10 )
         );
  NOR2_X1 \SubCellInst3_LFInst_9_LFInst_0_U6  ( .A1(PermutationOutput3[37]), 
        .A2(\SubCellInst3_LFInst_9_LFInst_0_n9 ), .ZN(
        \SubCellInst3_LFInst_9_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst3_LFInst_9_LFInst_0_U5  ( .A1(
        \SubCellInst3_LFInst_9_LFInst_0_n8 ), .A2(
        \SubCellInst3_LFInst_9_LFInst_0_n7 ), .ZN(
        \SubCellInst3_LFInst_9_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst3_LFInst_9_LFInst_0_U4  ( .A1(PermutationOutput3[39]), 
        .A2(PermutationOutput3[38]), .ZN(\SubCellInst3_LFInst_9_LFInst_0_n7 )
         );
  INV_X1 \SubCellInst3_LFInst_9_LFInst_0_U3  ( .A(PermutationOutput3[36]), 
        .ZN(\SubCellInst3_LFInst_9_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst3_LFInst_9_LFInst_1_U6  ( .A1(
        \SubCellInst3_LFInst_9_LFInst_1_n6 ), .A2(
        \SubCellInst3_LFInst_9_LFInst_1_n5 ), .ZN(Output[37]) );
  NAND2_X1 \SubCellInst3_LFInst_9_LFInst_1_U5  ( .A1(PermutationOutput3[38]), 
        .A2(PermutationOutput3[36]), .ZN(\SubCellInst3_LFInst_9_LFInst_1_n5 )
         );
  OR2_X1 \SubCellInst3_LFInst_9_LFInst_1_U4  ( .A1(PermutationOutput3[39]), 
        .A2(\SubCellInst3_LFInst_9_LFInst_1_n4 ), .ZN(
        \SubCellInst3_LFInst_9_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst3_LFInst_9_LFInst_1_U3  ( .A1(PermutationOutput3[38]), 
        .A2(PermutationOutput3[36]), .ZN(\SubCellInst3_LFInst_9_LFInst_1_n4 )
         );
  NAND2_X1 \SubCellInst3_LFInst_9_LFInst_2_U8  ( .A1(
        \SubCellInst3_LFInst_9_LFInst_2_n11 ), .A2(
        \SubCellInst3_LFInst_9_LFInst_2_n10 ), .ZN(Output[38]) );
  OR2_X1 \SubCellInst3_LFInst_9_LFInst_2_U7  ( .A1(PermutationOutput3[36]), 
        .A2(PermutationOutput3[39]), .ZN(\SubCellInst3_LFInst_9_LFInst_2_n10 )
         );
  NAND2_X1 \SubCellInst3_LFInst_9_LFInst_2_U6  ( .A1(PermutationOutput3[37]), 
        .A2(\SubCellInst3_LFInst_9_LFInst_2_n9 ), .ZN(
        \SubCellInst3_LFInst_9_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst3_LFInst_9_LFInst_2_U5  ( .A1(
        \SubCellInst3_LFInst_9_LFInst_2_n8 ), .A2(
        \SubCellInst3_LFInst_9_LFInst_2_n7 ), .ZN(
        \SubCellInst3_LFInst_9_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst3_LFInst_9_LFInst_2_U4  ( .A1(PermutationOutput3[36]), 
        .A2(PermutationOutput3[39]), .ZN(\SubCellInst3_LFInst_9_LFInst_2_n7 )
         );
  INV_X1 \SubCellInst3_LFInst_9_LFInst_2_U3  ( .A(PermutationOutput3[38]), 
        .ZN(\SubCellInst3_LFInst_9_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst3_LFInst_9_LFInst_3_U6  ( .A1(
        \SubCellInst3_LFInst_9_LFInst_3_n6 ), .A2(
        \SubCellInst3_LFInst_9_LFInst_3_n5 ), .ZN(Output[39]) );
  NOR2_X1 \SubCellInst3_LFInst_9_LFInst_3_U5  ( .A1(PermutationOutput3[39]), 
        .A2(PermutationOutput3[36]), .ZN(\SubCellInst3_LFInst_9_LFInst_3_n5 )
         );
  NOR2_X1 \SubCellInst3_LFInst_9_LFInst_3_U4  ( .A1(PermutationOutput3[37]), 
        .A2(\SubCellInst3_LFInst_9_LFInst_3_n4 ), .ZN(
        \SubCellInst3_LFInst_9_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst3_LFInst_9_LFInst_3_U3  ( .A1(PermutationOutput3[39]), 
        .A2(PermutationOutput3[38]), .ZN(\SubCellInst3_LFInst_9_LFInst_3_n4 )
         );
  NOR2_X1 \SubCellInst3_LFInst_10_LFInst_0_U8  ( .A1(
        \SubCellInst3_LFInst_10_LFInst_0_n11 ), .A2(
        \SubCellInst3_LFInst_10_LFInst_0_n10 ), .ZN(Output[40]) );
  AND2_X1 \SubCellInst3_LFInst_10_LFInst_0_U7  ( .A1(PermutationOutput3[43]), 
        .A2(PermutationOutput3[42]), .ZN(\SubCellInst3_LFInst_10_LFInst_0_n10 ) );
  NOR2_X1 \SubCellInst3_LFInst_10_LFInst_0_U6  ( .A1(PermutationOutput3[41]), 
        .A2(\SubCellInst3_LFInst_10_LFInst_0_n9 ), .ZN(
        \SubCellInst3_LFInst_10_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst3_LFInst_10_LFInst_0_U5  ( .A1(
        \SubCellInst3_LFInst_10_LFInst_0_n8 ), .A2(
        \SubCellInst3_LFInst_10_LFInst_0_n7 ), .ZN(
        \SubCellInst3_LFInst_10_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst3_LFInst_10_LFInst_0_U4  ( .A1(PermutationOutput3[43]), 
        .A2(PermutationOutput3[42]), .ZN(\SubCellInst3_LFInst_10_LFInst_0_n7 )
         );
  INV_X1 \SubCellInst3_LFInst_10_LFInst_0_U3  ( .A(PermutationOutput3[40]), 
        .ZN(\SubCellInst3_LFInst_10_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst3_LFInst_10_LFInst_1_U6  ( .A1(
        \SubCellInst3_LFInst_10_LFInst_1_n6 ), .A2(
        \SubCellInst3_LFInst_10_LFInst_1_n5 ), .ZN(Output[41]) );
  NAND2_X1 \SubCellInst3_LFInst_10_LFInst_1_U5  ( .A1(PermutationOutput3[42]), 
        .A2(PermutationOutput3[40]), .ZN(\SubCellInst3_LFInst_10_LFInst_1_n5 )
         );
  OR2_X1 \SubCellInst3_LFInst_10_LFInst_1_U4  ( .A1(PermutationOutput3[43]), 
        .A2(\SubCellInst3_LFInst_10_LFInst_1_n4 ), .ZN(
        \SubCellInst3_LFInst_10_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst3_LFInst_10_LFInst_1_U3  ( .A1(PermutationOutput3[42]), 
        .A2(PermutationOutput3[40]), .ZN(\SubCellInst3_LFInst_10_LFInst_1_n4 )
         );
  NAND2_X1 \SubCellInst3_LFInst_10_LFInst_2_U8  ( .A1(
        \SubCellInst3_LFInst_10_LFInst_2_n11 ), .A2(
        \SubCellInst3_LFInst_10_LFInst_2_n10 ), .ZN(Output[42]) );
  OR2_X1 \SubCellInst3_LFInst_10_LFInst_2_U7  ( .A1(PermutationOutput3[40]), 
        .A2(PermutationOutput3[43]), .ZN(\SubCellInst3_LFInst_10_LFInst_2_n10 ) );
  NAND2_X1 \SubCellInst3_LFInst_10_LFInst_2_U6  ( .A1(PermutationOutput3[41]), 
        .A2(\SubCellInst3_LFInst_10_LFInst_2_n9 ), .ZN(
        \SubCellInst3_LFInst_10_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst3_LFInst_10_LFInst_2_U5  ( .A1(
        \SubCellInst3_LFInst_10_LFInst_2_n8 ), .A2(
        \SubCellInst3_LFInst_10_LFInst_2_n7 ), .ZN(
        \SubCellInst3_LFInst_10_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst3_LFInst_10_LFInst_2_U4  ( .A1(PermutationOutput3[40]), 
        .A2(PermutationOutput3[43]), .ZN(\SubCellInst3_LFInst_10_LFInst_2_n7 )
         );
  INV_X1 \SubCellInst3_LFInst_10_LFInst_2_U3  ( .A(PermutationOutput3[42]), 
        .ZN(\SubCellInst3_LFInst_10_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst3_LFInst_10_LFInst_3_U6  ( .A1(
        \SubCellInst3_LFInst_10_LFInst_3_n6 ), .A2(
        \SubCellInst3_LFInst_10_LFInst_3_n5 ), .ZN(Output[43]) );
  NOR2_X1 \SubCellInst3_LFInst_10_LFInst_3_U5  ( .A1(PermutationOutput3[43]), 
        .A2(PermutationOutput3[40]), .ZN(\SubCellInst3_LFInst_10_LFInst_3_n5 )
         );
  NOR2_X1 \SubCellInst3_LFInst_10_LFInst_3_U4  ( .A1(PermutationOutput3[41]), 
        .A2(\SubCellInst3_LFInst_10_LFInst_3_n4 ), .ZN(
        \SubCellInst3_LFInst_10_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst3_LFInst_10_LFInst_3_U3  ( .A1(PermutationOutput3[43]), 
        .A2(PermutationOutput3[42]), .ZN(\SubCellInst3_LFInst_10_LFInst_3_n4 )
         );
  NOR2_X1 \SubCellInst3_LFInst_11_LFInst_0_U8  ( .A1(
        \SubCellInst3_LFInst_11_LFInst_0_n11 ), .A2(
        \SubCellInst3_LFInst_11_LFInst_0_n10 ), .ZN(Output[44]) );
  AND2_X1 \SubCellInst3_LFInst_11_LFInst_0_U7  ( .A1(PermutationOutput3[47]), 
        .A2(PermutationOutput3[46]), .ZN(\SubCellInst3_LFInst_11_LFInst_0_n10 ) );
  NOR2_X1 \SubCellInst3_LFInst_11_LFInst_0_U6  ( .A1(PermutationOutput3[45]), 
        .A2(\SubCellInst3_LFInst_11_LFInst_0_n9 ), .ZN(
        \SubCellInst3_LFInst_11_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst3_LFInst_11_LFInst_0_U5  ( .A1(
        \SubCellInst3_LFInst_11_LFInst_0_n8 ), .A2(
        \SubCellInst3_LFInst_11_LFInst_0_n7 ), .ZN(
        \SubCellInst3_LFInst_11_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst3_LFInst_11_LFInst_0_U4  ( .A1(PermutationOutput3[47]), 
        .A2(PermutationOutput3[46]), .ZN(\SubCellInst3_LFInst_11_LFInst_0_n7 )
         );
  INV_X1 \SubCellInst3_LFInst_11_LFInst_0_U3  ( .A(PermutationOutput3[44]), 
        .ZN(\SubCellInst3_LFInst_11_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst3_LFInst_11_LFInst_1_U6  ( .A1(
        \SubCellInst3_LFInst_11_LFInst_1_n6 ), .A2(
        \SubCellInst3_LFInst_11_LFInst_1_n5 ), .ZN(Output[45]) );
  NAND2_X1 \SubCellInst3_LFInst_11_LFInst_1_U5  ( .A1(PermutationOutput3[46]), 
        .A2(PermutationOutput3[44]), .ZN(\SubCellInst3_LFInst_11_LFInst_1_n5 )
         );
  OR2_X1 \SubCellInst3_LFInst_11_LFInst_1_U4  ( .A1(PermutationOutput3[47]), 
        .A2(\SubCellInst3_LFInst_11_LFInst_1_n4 ), .ZN(
        \SubCellInst3_LFInst_11_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst3_LFInst_11_LFInst_1_U3  ( .A1(PermutationOutput3[46]), 
        .A2(PermutationOutput3[44]), .ZN(\SubCellInst3_LFInst_11_LFInst_1_n4 )
         );
  NAND2_X1 \SubCellInst3_LFInst_11_LFInst_2_U8  ( .A1(
        \SubCellInst3_LFInst_11_LFInst_2_n11 ), .A2(
        \SubCellInst3_LFInst_11_LFInst_2_n10 ), .ZN(Output[46]) );
  OR2_X1 \SubCellInst3_LFInst_11_LFInst_2_U7  ( .A1(PermutationOutput3[44]), 
        .A2(PermutationOutput3[47]), .ZN(\SubCellInst3_LFInst_11_LFInst_2_n10 ) );
  NAND2_X1 \SubCellInst3_LFInst_11_LFInst_2_U6  ( .A1(PermutationOutput3[45]), 
        .A2(\SubCellInst3_LFInst_11_LFInst_2_n9 ), .ZN(
        \SubCellInst3_LFInst_11_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst3_LFInst_11_LFInst_2_U5  ( .A1(
        \SubCellInst3_LFInst_11_LFInst_2_n8 ), .A2(
        \SubCellInst3_LFInst_11_LFInst_2_n7 ), .ZN(
        \SubCellInst3_LFInst_11_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst3_LFInst_11_LFInst_2_U4  ( .A1(PermutationOutput3[44]), 
        .A2(PermutationOutput3[47]), .ZN(\SubCellInst3_LFInst_11_LFInst_2_n7 )
         );
  INV_X1 \SubCellInst3_LFInst_11_LFInst_2_U3  ( .A(PermutationOutput3[46]), 
        .ZN(\SubCellInst3_LFInst_11_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst3_LFInst_11_LFInst_3_U6  ( .A1(
        \SubCellInst3_LFInst_11_LFInst_3_n6 ), .A2(
        \SubCellInst3_LFInst_11_LFInst_3_n5 ), .ZN(Output[47]) );
  NOR2_X1 \SubCellInst3_LFInst_11_LFInst_3_U5  ( .A1(PermutationOutput3[47]), 
        .A2(PermutationOutput3[44]), .ZN(\SubCellInst3_LFInst_11_LFInst_3_n5 )
         );
  NOR2_X1 \SubCellInst3_LFInst_11_LFInst_3_U4  ( .A1(PermutationOutput3[45]), 
        .A2(\SubCellInst3_LFInst_11_LFInst_3_n4 ), .ZN(
        \SubCellInst3_LFInst_11_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst3_LFInst_11_LFInst_3_U3  ( .A1(PermutationOutput3[47]), 
        .A2(PermutationOutput3[46]), .ZN(\SubCellInst3_LFInst_11_LFInst_3_n4 )
         );
  NOR2_X1 \SubCellInst3_LFInst_12_LFInst_0_U8  ( .A1(
        \SubCellInst3_LFInst_12_LFInst_0_n11 ), .A2(
        \SubCellInst3_LFInst_12_LFInst_0_n10 ), .ZN(Output[48]) );
  AND2_X1 \SubCellInst3_LFInst_12_LFInst_0_U7  ( .A1(PermutationOutput3[51]), 
        .A2(PermutationOutput3[50]), .ZN(\SubCellInst3_LFInst_12_LFInst_0_n10 ) );
  NOR2_X1 \SubCellInst3_LFInst_12_LFInst_0_U6  ( .A1(PermutationOutput3[49]), 
        .A2(\SubCellInst3_LFInst_12_LFInst_0_n9 ), .ZN(
        \SubCellInst3_LFInst_12_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst3_LFInst_12_LFInst_0_U5  ( .A1(
        \SubCellInst3_LFInst_12_LFInst_0_n8 ), .A2(
        \SubCellInst3_LFInst_12_LFInst_0_n7 ), .ZN(
        \SubCellInst3_LFInst_12_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst3_LFInst_12_LFInst_0_U4  ( .A1(PermutationOutput3[51]), 
        .A2(PermutationOutput3[50]), .ZN(\SubCellInst3_LFInst_12_LFInst_0_n7 )
         );
  INV_X1 \SubCellInst3_LFInst_12_LFInst_0_U3  ( .A(PermutationOutput3[48]), 
        .ZN(\SubCellInst3_LFInst_12_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst3_LFInst_12_LFInst_1_U6  ( .A1(
        \SubCellInst3_LFInst_12_LFInst_1_n6 ), .A2(
        \SubCellInst3_LFInst_12_LFInst_1_n5 ), .ZN(Output[49]) );
  NAND2_X1 \SubCellInst3_LFInst_12_LFInst_1_U5  ( .A1(PermutationOutput3[50]), 
        .A2(PermutationOutput3[48]), .ZN(\SubCellInst3_LFInst_12_LFInst_1_n5 )
         );
  OR2_X1 \SubCellInst3_LFInst_12_LFInst_1_U4  ( .A1(PermutationOutput3[51]), 
        .A2(\SubCellInst3_LFInst_12_LFInst_1_n4 ), .ZN(
        \SubCellInst3_LFInst_12_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst3_LFInst_12_LFInst_1_U3  ( .A1(PermutationOutput3[50]), 
        .A2(PermutationOutput3[48]), .ZN(\SubCellInst3_LFInst_12_LFInst_1_n4 )
         );
  NAND2_X1 \SubCellInst3_LFInst_12_LFInst_2_U8  ( .A1(
        \SubCellInst3_LFInst_12_LFInst_2_n11 ), .A2(
        \SubCellInst3_LFInst_12_LFInst_2_n10 ), .ZN(Output[50]) );
  OR2_X1 \SubCellInst3_LFInst_12_LFInst_2_U7  ( .A1(PermutationOutput3[48]), 
        .A2(PermutationOutput3[51]), .ZN(\SubCellInst3_LFInst_12_LFInst_2_n10 ) );
  NAND2_X1 \SubCellInst3_LFInst_12_LFInst_2_U6  ( .A1(PermutationOutput3[49]), 
        .A2(\SubCellInst3_LFInst_12_LFInst_2_n9 ), .ZN(
        \SubCellInst3_LFInst_12_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst3_LFInst_12_LFInst_2_U5  ( .A1(
        \SubCellInst3_LFInst_12_LFInst_2_n8 ), .A2(
        \SubCellInst3_LFInst_12_LFInst_2_n7 ), .ZN(
        \SubCellInst3_LFInst_12_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst3_LFInst_12_LFInst_2_U4  ( .A1(PermutationOutput3[48]), 
        .A2(PermutationOutput3[51]), .ZN(\SubCellInst3_LFInst_12_LFInst_2_n7 )
         );
  INV_X1 \SubCellInst3_LFInst_12_LFInst_2_U3  ( .A(PermutationOutput3[50]), 
        .ZN(\SubCellInst3_LFInst_12_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst3_LFInst_12_LFInst_3_U6  ( .A1(
        \SubCellInst3_LFInst_12_LFInst_3_n6 ), .A2(
        \SubCellInst3_LFInst_12_LFInst_3_n5 ), .ZN(Output[51]) );
  NOR2_X1 \SubCellInst3_LFInst_12_LFInst_3_U5  ( .A1(PermutationOutput3[51]), 
        .A2(PermutationOutput3[48]), .ZN(\SubCellInst3_LFInst_12_LFInst_3_n5 )
         );
  NOR2_X1 \SubCellInst3_LFInst_12_LFInst_3_U4  ( .A1(PermutationOutput3[49]), 
        .A2(\SubCellInst3_LFInst_12_LFInst_3_n4 ), .ZN(
        \SubCellInst3_LFInst_12_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst3_LFInst_12_LFInst_3_U3  ( .A1(PermutationOutput3[51]), 
        .A2(PermutationOutput3[50]), .ZN(\SubCellInst3_LFInst_12_LFInst_3_n4 )
         );
  NOR2_X1 \SubCellInst3_LFInst_13_LFInst_0_U8  ( .A1(
        \SubCellInst3_LFInst_13_LFInst_0_n11 ), .A2(
        \SubCellInst3_LFInst_13_LFInst_0_n10 ), .ZN(Output[52]) );
  AND2_X1 \SubCellInst3_LFInst_13_LFInst_0_U7  ( .A1(PermutationOutput3[55]), 
        .A2(PermutationOutput3[54]), .ZN(\SubCellInst3_LFInst_13_LFInst_0_n10 ) );
  NOR2_X1 \SubCellInst3_LFInst_13_LFInst_0_U6  ( .A1(PermutationOutput3[53]), 
        .A2(\SubCellInst3_LFInst_13_LFInst_0_n9 ), .ZN(
        \SubCellInst3_LFInst_13_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst3_LFInst_13_LFInst_0_U5  ( .A1(
        \SubCellInst3_LFInst_13_LFInst_0_n8 ), .A2(
        \SubCellInst3_LFInst_13_LFInst_0_n7 ), .ZN(
        \SubCellInst3_LFInst_13_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst3_LFInst_13_LFInst_0_U4  ( .A1(PermutationOutput3[55]), 
        .A2(PermutationOutput3[54]), .ZN(\SubCellInst3_LFInst_13_LFInst_0_n7 )
         );
  INV_X1 \SubCellInst3_LFInst_13_LFInst_0_U3  ( .A(PermutationOutput3[52]), 
        .ZN(\SubCellInst3_LFInst_13_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst3_LFInst_13_LFInst_1_U6  ( .A1(
        \SubCellInst3_LFInst_13_LFInst_1_n6 ), .A2(
        \SubCellInst3_LFInst_13_LFInst_1_n5 ), .ZN(Output[53]) );
  NAND2_X1 \SubCellInst3_LFInst_13_LFInst_1_U5  ( .A1(PermutationOutput3[54]), 
        .A2(PermutationOutput3[52]), .ZN(\SubCellInst3_LFInst_13_LFInst_1_n5 )
         );
  OR2_X1 \SubCellInst3_LFInst_13_LFInst_1_U4  ( .A1(PermutationOutput3[55]), 
        .A2(\SubCellInst3_LFInst_13_LFInst_1_n4 ), .ZN(
        \SubCellInst3_LFInst_13_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst3_LFInst_13_LFInst_1_U3  ( .A1(PermutationOutput3[54]), 
        .A2(PermutationOutput3[52]), .ZN(\SubCellInst3_LFInst_13_LFInst_1_n4 )
         );
  NAND2_X1 \SubCellInst3_LFInst_13_LFInst_2_U8  ( .A1(
        \SubCellInst3_LFInst_13_LFInst_2_n11 ), .A2(
        \SubCellInst3_LFInst_13_LFInst_2_n10 ), .ZN(Output[54]) );
  OR2_X1 \SubCellInst3_LFInst_13_LFInst_2_U7  ( .A1(PermutationOutput3[52]), 
        .A2(PermutationOutput3[55]), .ZN(\SubCellInst3_LFInst_13_LFInst_2_n10 ) );
  NAND2_X1 \SubCellInst3_LFInst_13_LFInst_2_U6  ( .A1(PermutationOutput3[53]), 
        .A2(\SubCellInst3_LFInst_13_LFInst_2_n9 ), .ZN(
        \SubCellInst3_LFInst_13_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst3_LFInst_13_LFInst_2_U5  ( .A1(
        \SubCellInst3_LFInst_13_LFInst_2_n8 ), .A2(
        \SubCellInst3_LFInst_13_LFInst_2_n7 ), .ZN(
        \SubCellInst3_LFInst_13_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst3_LFInst_13_LFInst_2_U4  ( .A1(PermutationOutput3[52]), 
        .A2(PermutationOutput3[55]), .ZN(\SubCellInst3_LFInst_13_LFInst_2_n7 )
         );
  INV_X1 \SubCellInst3_LFInst_13_LFInst_2_U3  ( .A(PermutationOutput3[54]), 
        .ZN(\SubCellInst3_LFInst_13_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst3_LFInst_13_LFInst_3_U6  ( .A1(
        \SubCellInst3_LFInst_13_LFInst_3_n6 ), .A2(
        \SubCellInst3_LFInst_13_LFInst_3_n5 ), .ZN(Output[55]) );
  NOR2_X1 \SubCellInst3_LFInst_13_LFInst_3_U5  ( .A1(PermutationOutput3[55]), 
        .A2(PermutationOutput3[52]), .ZN(\SubCellInst3_LFInst_13_LFInst_3_n5 )
         );
  NOR2_X1 \SubCellInst3_LFInst_13_LFInst_3_U4  ( .A1(PermutationOutput3[53]), 
        .A2(\SubCellInst3_LFInst_13_LFInst_3_n4 ), .ZN(
        \SubCellInst3_LFInst_13_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst3_LFInst_13_LFInst_3_U3  ( .A1(PermutationOutput3[55]), 
        .A2(PermutationOutput3[54]), .ZN(\SubCellInst3_LFInst_13_LFInst_3_n4 )
         );
  NOR2_X1 \SubCellInst3_LFInst_14_LFInst_0_U8  ( .A1(
        \SubCellInst3_LFInst_14_LFInst_0_n11 ), .A2(
        \SubCellInst3_LFInst_14_LFInst_0_n10 ), .ZN(Output[56]) );
  AND2_X1 \SubCellInst3_LFInst_14_LFInst_0_U7  ( .A1(PermutationOutput3[59]), 
        .A2(PermutationOutput3[58]), .ZN(\SubCellInst3_LFInst_14_LFInst_0_n10 ) );
  NOR2_X1 \SubCellInst3_LFInst_14_LFInst_0_U6  ( .A1(PermutationOutput3[57]), 
        .A2(\SubCellInst3_LFInst_14_LFInst_0_n9 ), .ZN(
        \SubCellInst3_LFInst_14_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst3_LFInst_14_LFInst_0_U5  ( .A1(
        \SubCellInst3_LFInst_14_LFInst_0_n8 ), .A2(
        \SubCellInst3_LFInst_14_LFInst_0_n7 ), .ZN(
        \SubCellInst3_LFInst_14_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst3_LFInst_14_LFInst_0_U4  ( .A1(PermutationOutput3[59]), 
        .A2(PermutationOutput3[58]), .ZN(\SubCellInst3_LFInst_14_LFInst_0_n7 )
         );
  INV_X1 \SubCellInst3_LFInst_14_LFInst_0_U3  ( .A(PermutationOutput3[56]), 
        .ZN(\SubCellInst3_LFInst_14_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst3_LFInst_14_LFInst_1_U6  ( .A1(
        \SubCellInst3_LFInst_14_LFInst_1_n6 ), .A2(
        \SubCellInst3_LFInst_14_LFInst_1_n5 ), .ZN(Output[57]) );
  NAND2_X1 \SubCellInst3_LFInst_14_LFInst_1_U5  ( .A1(PermutationOutput3[58]), 
        .A2(PermutationOutput3[56]), .ZN(\SubCellInst3_LFInst_14_LFInst_1_n5 )
         );
  OR2_X1 \SubCellInst3_LFInst_14_LFInst_1_U4  ( .A1(PermutationOutput3[59]), 
        .A2(\SubCellInst3_LFInst_14_LFInst_1_n4 ), .ZN(
        \SubCellInst3_LFInst_14_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst3_LFInst_14_LFInst_1_U3  ( .A1(PermutationOutput3[58]), 
        .A2(PermutationOutput3[56]), .ZN(\SubCellInst3_LFInst_14_LFInst_1_n4 )
         );
  NAND2_X1 \SubCellInst3_LFInst_14_LFInst_2_U8  ( .A1(
        \SubCellInst3_LFInst_14_LFInst_2_n11 ), .A2(
        \SubCellInst3_LFInst_14_LFInst_2_n10 ), .ZN(Output[58]) );
  OR2_X1 \SubCellInst3_LFInst_14_LFInst_2_U7  ( .A1(PermutationOutput3[56]), 
        .A2(PermutationOutput3[59]), .ZN(\SubCellInst3_LFInst_14_LFInst_2_n10 ) );
  NAND2_X1 \SubCellInst3_LFInst_14_LFInst_2_U6  ( .A1(PermutationOutput3[57]), 
        .A2(\SubCellInst3_LFInst_14_LFInst_2_n9 ), .ZN(
        \SubCellInst3_LFInst_14_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst3_LFInst_14_LFInst_2_U5  ( .A1(
        \SubCellInst3_LFInst_14_LFInst_2_n8 ), .A2(
        \SubCellInst3_LFInst_14_LFInst_2_n7 ), .ZN(
        \SubCellInst3_LFInst_14_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst3_LFInst_14_LFInst_2_U4  ( .A1(PermutationOutput3[56]), 
        .A2(PermutationOutput3[59]), .ZN(\SubCellInst3_LFInst_14_LFInst_2_n7 )
         );
  INV_X1 \SubCellInst3_LFInst_14_LFInst_2_U3  ( .A(PermutationOutput3[58]), 
        .ZN(\SubCellInst3_LFInst_14_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst3_LFInst_14_LFInst_3_U6  ( .A1(
        \SubCellInst3_LFInst_14_LFInst_3_n6 ), .A2(
        \SubCellInst3_LFInst_14_LFInst_3_n5 ), .ZN(Output[59]) );
  NOR2_X1 \SubCellInst3_LFInst_14_LFInst_3_U5  ( .A1(PermutationOutput3[59]), 
        .A2(PermutationOutput3[56]), .ZN(\SubCellInst3_LFInst_14_LFInst_3_n5 )
         );
  NOR2_X1 \SubCellInst3_LFInst_14_LFInst_3_U4  ( .A1(PermutationOutput3[57]), 
        .A2(\SubCellInst3_LFInst_14_LFInst_3_n4 ), .ZN(
        \SubCellInst3_LFInst_14_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst3_LFInst_14_LFInst_3_U3  ( .A1(PermutationOutput3[59]), 
        .A2(PermutationOutput3[58]), .ZN(\SubCellInst3_LFInst_14_LFInst_3_n4 )
         );
  NOR2_X1 \SubCellInst3_LFInst_15_LFInst_0_U8  ( .A1(
        \SubCellInst3_LFInst_15_LFInst_0_n11 ), .A2(
        \SubCellInst3_LFInst_15_LFInst_0_n10 ), .ZN(Output[60]) );
  AND2_X1 \SubCellInst3_LFInst_15_LFInst_0_U7  ( .A1(PermutationOutput3[63]), 
        .A2(PermutationOutput3[62]), .ZN(\SubCellInst3_LFInst_15_LFInst_0_n10 ) );
  NOR2_X1 \SubCellInst3_LFInst_15_LFInst_0_U6  ( .A1(PermutationOutput3[61]), 
        .A2(\SubCellInst3_LFInst_15_LFInst_0_n9 ), .ZN(
        \SubCellInst3_LFInst_15_LFInst_0_n11 ) );
  NOR2_X1 \SubCellInst3_LFInst_15_LFInst_0_U5  ( .A1(
        \SubCellInst3_LFInst_15_LFInst_0_n8 ), .A2(
        \SubCellInst3_LFInst_15_LFInst_0_n7 ), .ZN(
        \SubCellInst3_LFInst_15_LFInst_0_n9 ) );
  NOR2_X1 \SubCellInst3_LFInst_15_LFInst_0_U4  ( .A1(PermutationOutput3[63]), 
        .A2(PermutationOutput3[62]), .ZN(\SubCellInst3_LFInst_15_LFInst_0_n7 )
         );
  INV_X1 \SubCellInst3_LFInst_15_LFInst_0_U3  ( .A(PermutationOutput3[60]), 
        .ZN(\SubCellInst3_LFInst_15_LFInst_0_n8 ) );
  NAND2_X1 \SubCellInst3_LFInst_15_LFInst_1_U6  ( .A1(
        \SubCellInst3_LFInst_15_LFInst_1_n6 ), .A2(
        \SubCellInst3_LFInst_15_LFInst_1_n5 ), .ZN(Output[61]) );
  NAND2_X1 \SubCellInst3_LFInst_15_LFInst_1_U5  ( .A1(PermutationOutput3[62]), 
        .A2(PermutationOutput3[60]), .ZN(\SubCellInst3_LFInst_15_LFInst_1_n5 )
         );
  OR2_X1 \SubCellInst3_LFInst_15_LFInst_1_U4  ( .A1(PermutationOutput3[63]), 
        .A2(\SubCellInst3_LFInst_15_LFInst_1_n4 ), .ZN(
        \SubCellInst3_LFInst_15_LFInst_1_n6 ) );
  NOR2_X1 \SubCellInst3_LFInst_15_LFInst_1_U3  ( .A1(PermutationOutput3[62]), 
        .A2(PermutationOutput3[60]), .ZN(\SubCellInst3_LFInst_15_LFInst_1_n4 )
         );
  NAND2_X1 \SubCellInst3_LFInst_15_LFInst_2_U8  ( .A1(
        \SubCellInst3_LFInst_15_LFInst_2_n11 ), .A2(
        \SubCellInst3_LFInst_15_LFInst_2_n10 ), .ZN(Output[62]) );
  OR2_X1 \SubCellInst3_LFInst_15_LFInst_2_U7  ( .A1(PermutationOutput3[60]), 
        .A2(PermutationOutput3[63]), .ZN(\SubCellInst3_LFInst_15_LFInst_2_n10 ) );
  NAND2_X1 \SubCellInst3_LFInst_15_LFInst_2_U6  ( .A1(PermutationOutput3[61]), 
        .A2(\SubCellInst3_LFInst_15_LFInst_2_n9 ), .ZN(
        \SubCellInst3_LFInst_15_LFInst_2_n11 ) );
  NAND2_X1 \SubCellInst3_LFInst_15_LFInst_2_U5  ( .A1(
        \SubCellInst3_LFInst_15_LFInst_2_n8 ), .A2(
        \SubCellInst3_LFInst_15_LFInst_2_n7 ), .ZN(
        \SubCellInst3_LFInst_15_LFInst_2_n9 ) );
  NAND2_X1 \SubCellInst3_LFInst_15_LFInst_2_U4  ( .A1(PermutationOutput3[60]), 
        .A2(PermutationOutput3[63]), .ZN(\SubCellInst3_LFInst_15_LFInst_2_n7 )
         );
  INV_X1 \SubCellInst3_LFInst_15_LFInst_2_U3  ( .A(PermutationOutput3[62]), 
        .ZN(\SubCellInst3_LFInst_15_LFInst_2_n8 ) );
  OR2_X1 \SubCellInst3_LFInst_15_LFInst_3_U6  ( .A1(
        \SubCellInst3_LFInst_15_LFInst_3_n6 ), .A2(
        \SubCellInst3_LFInst_15_LFInst_3_n5 ), .ZN(Output[63]) );
  NOR2_X1 \SubCellInst3_LFInst_15_LFInst_3_U5  ( .A1(PermutationOutput3[63]), 
        .A2(PermutationOutput3[60]), .ZN(\SubCellInst3_LFInst_15_LFInst_3_n5 )
         );
  NOR2_X1 \SubCellInst3_LFInst_15_LFInst_3_U4  ( .A1(PermutationOutput3[61]), 
        .A2(\SubCellInst3_LFInst_15_LFInst_3_n4 ), .ZN(
        \SubCellInst3_LFInst_15_LFInst_3_n6 ) );
  AND2_X1 \SubCellInst3_LFInst_15_LFInst_3_U3  ( .A1(PermutationOutput3[63]), 
        .A2(PermutationOutput3[62]), .ZN(\SubCellInst3_LFInst_15_LFInst_3_n4 )
         );
  XNOR2_X1 \Red_PlaintextInst_LFInst_0_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_0_LFInst_0_n2 ), .B(Input[2]), .ZN(
        Red_MCOutput[0]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_0_LFInst_0_U3  ( .A(Input[3]), .B(
        Input[1]), .ZN(\Red_PlaintextInst_LFInst_0_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_0_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_0_LFInst_1_n2 ), .B(Input[2]), .ZN(
        Red_MCOutput[1]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_0_LFInst_1_U3  ( .A(Input[3]), .B(
        Input[0]), .ZN(\Red_PlaintextInst_LFInst_0_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_0_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_0_LFInst_2_n2 ), .B(Input[1]), .ZN(
        Red_MCOutput[2]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_0_LFInst_2_U3  ( .A(Input[3]), .B(
        Input[0]), .ZN(\Red_PlaintextInst_LFInst_0_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_0_LFInst_3_U4  ( .A(
        \Red_PlaintextInst_LFInst_0_LFInst_3_n2 ), .B(Input[1]), .ZN(
        Red_MCOutput[3]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_0_LFInst_3_U3  ( .A(Input[2]), .B(
        Input[0]), .ZN(\Red_PlaintextInst_LFInst_0_LFInst_3_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_1_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_1_LFInst_0_n2 ), .B(Input[6]), .ZN(
        Red_MCOutput[4]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_1_LFInst_0_U3  ( .A(Input[7]), .B(
        Input[5]), .ZN(\Red_PlaintextInst_LFInst_1_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_1_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_1_LFInst_1_n2 ), .B(Input[6]), .ZN(
        Red_MCOutput[5]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_1_LFInst_1_U3  ( .A(Input[7]), .B(
        Input[4]), .ZN(\Red_PlaintextInst_LFInst_1_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_1_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_1_LFInst_2_n2 ), .B(Input[5]), .ZN(
        Red_MCOutput[6]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_1_LFInst_2_U3  ( .A(Input[7]), .B(
        Input[4]), .ZN(\Red_PlaintextInst_LFInst_1_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_1_LFInst_3_U4  ( .A(
        \Red_PlaintextInst_LFInst_1_LFInst_3_n2 ), .B(Input[5]), .ZN(
        Red_MCOutput[7]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_1_LFInst_3_U3  ( .A(Input[6]), .B(
        Input[4]), .ZN(\Red_PlaintextInst_LFInst_1_LFInst_3_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_2_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_2_LFInst_0_n2 ), .B(Input[10]), .ZN(
        Red_MCOutput[8]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_2_LFInst_0_U3  ( .A(Input[11]), .B(
        Input[9]), .ZN(\Red_PlaintextInst_LFInst_2_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_2_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_2_LFInst_1_n2 ), .B(Input[10]), .ZN(
        Red_MCOutput[9]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_2_LFInst_1_U3  ( .A(Input[11]), .B(
        Input[8]), .ZN(\Red_PlaintextInst_LFInst_2_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_2_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_2_LFInst_2_n2 ), .B(Input[9]), .ZN(
        Red_MCOutput[10]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_2_LFInst_2_U3  ( .A(Input[11]), .B(
        Input[8]), .ZN(\Red_PlaintextInst_LFInst_2_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_2_LFInst_3_U4  ( .A(
        \Red_PlaintextInst_LFInst_2_LFInst_3_n2 ), .B(Input[9]), .ZN(
        Red_MCOutput[11]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_2_LFInst_3_U3  ( .A(Input[10]), .B(
        Input[8]), .ZN(\Red_PlaintextInst_LFInst_2_LFInst_3_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_3_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_3_LFInst_0_n2 ), .B(Input[14]), .ZN(
        Red_MCOutput[12]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_3_LFInst_0_U3  ( .A(Input[15]), .B(
        Input[13]), .ZN(\Red_PlaintextInst_LFInst_3_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_3_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_3_LFInst_1_n2 ), .B(Input[14]), .ZN(
        Red_MCOutput[13]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_3_LFInst_1_U3  ( .A(Input[15]), .B(
        Input[12]), .ZN(\Red_PlaintextInst_LFInst_3_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_3_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_3_LFInst_2_n2 ), .B(Input[13]), .ZN(
        Red_MCOutput[14]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_3_LFInst_2_U3  ( .A(Input[15]), .B(
        Input[12]), .ZN(\Red_PlaintextInst_LFInst_3_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_3_LFInst_3_U4  ( .A(
        \Red_PlaintextInst_LFInst_3_LFInst_3_n2 ), .B(Input[13]), .ZN(
        Red_MCOutput[15]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_3_LFInst_3_U3  ( .A(Input[14]), .B(
        Input[12]), .ZN(\Red_PlaintextInst_LFInst_3_LFInst_3_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_4_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_4_LFInst_0_n2 ), .B(Input[18]), .ZN(
        Red_MCOutput[16]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_4_LFInst_0_U3  ( .A(Input[19]), .B(
        Input[17]), .ZN(\Red_PlaintextInst_LFInst_4_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_4_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_4_LFInst_1_n2 ), .B(Input[18]), .ZN(
        Red_MCOutput[17]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_4_LFInst_1_U3  ( .A(Input[19]), .B(
        Input[16]), .ZN(\Red_PlaintextInst_LFInst_4_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_4_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_4_LFInst_2_n2 ), .B(Input[17]), .ZN(
        Red_MCOutput[18]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_4_LFInst_2_U3  ( .A(Input[19]), .B(
        Input[16]), .ZN(\Red_PlaintextInst_LFInst_4_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_4_LFInst_3_U4  ( .A(
        \Red_PlaintextInst_LFInst_4_LFInst_3_n2 ), .B(Input[17]), .ZN(
        Red_MCOutput[19]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_4_LFInst_3_U3  ( .A(Input[18]), .B(
        Input[16]), .ZN(\Red_PlaintextInst_LFInst_4_LFInst_3_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_5_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_5_LFInst_0_n2 ), .B(Input[22]), .ZN(
        Red_MCOutput[20]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_5_LFInst_0_U3  ( .A(Input[23]), .B(
        Input[21]), .ZN(\Red_PlaintextInst_LFInst_5_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_5_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_5_LFInst_1_n2 ), .B(Input[22]), .ZN(
        Red_MCOutput[21]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_5_LFInst_1_U3  ( .A(Input[23]), .B(
        Input[20]), .ZN(\Red_PlaintextInst_LFInst_5_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_5_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_5_LFInst_2_n2 ), .B(Input[21]), .ZN(
        Red_MCOutput[22]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_5_LFInst_2_U3  ( .A(Input[23]), .B(
        Input[20]), .ZN(\Red_PlaintextInst_LFInst_5_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_5_LFInst_3_U4  ( .A(
        \Red_PlaintextInst_LFInst_5_LFInst_3_n2 ), .B(Input[21]), .ZN(
        Red_MCOutput[23]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_5_LFInst_3_U3  ( .A(Input[22]), .B(
        Input[20]), .ZN(\Red_PlaintextInst_LFInst_5_LFInst_3_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_6_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_6_LFInst_0_n2 ), .B(Input[26]), .ZN(
        Red_MCOutput[24]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_6_LFInst_0_U3  ( .A(Input[27]), .B(
        Input[25]), .ZN(\Red_PlaintextInst_LFInst_6_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_6_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_6_LFInst_1_n2 ), .B(Input[26]), .ZN(
        Red_MCOutput[25]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_6_LFInst_1_U3  ( .A(Input[27]), .B(
        Input[24]), .ZN(\Red_PlaintextInst_LFInst_6_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_6_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_6_LFInst_2_n2 ), .B(Input[25]), .ZN(
        Red_MCOutput[26]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_6_LFInst_2_U3  ( .A(Input[27]), .B(
        Input[24]), .ZN(\Red_PlaintextInst_LFInst_6_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_6_LFInst_3_U4  ( .A(
        \Red_PlaintextInst_LFInst_6_LFInst_3_n2 ), .B(Input[25]), .ZN(
        Red_MCOutput[27]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_6_LFInst_3_U3  ( .A(Input[26]), .B(
        Input[24]), .ZN(\Red_PlaintextInst_LFInst_6_LFInst_3_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_7_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_7_LFInst_0_n2 ), .B(Input[30]), .ZN(
        Red_MCOutput[28]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_7_LFInst_0_U3  ( .A(Input[31]), .B(
        Input[29]), .ZN(\Red_PlaintextInst_LFInst_7_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_7_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_7_LFInst_1_n2 ), .B(Input[30]), .ZN(
        Red_MCOutput[29]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_7_LFInst_1_U3  ( .A(Input[31]), .B(
        Input[28]), .ZN(\Red_PlaintextInst_LFInst_7_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_7_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_7_LFInst_2_n2 ), .B(Input[29]), .ZN(
        Red_MCOutput[30]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_7_LFInst_2_U3  ( .A(Input[31]), .B(
        Input[28]), .ZN(\Red_PlaintextInst_LFInst_7_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_7_LFInst_3_U4  ( .A(
        \Red_PlaintextInst_LFInst_7_LFInst_3_n2 ), .B(Input[29]), .ZN(
        Red_MCOutput[31]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_7_LFInst_3_U3  ( .A(Input[30]), .B(
        Input[28]), .ZN(\Red_PlaintextInst_LFInst_7_LFInst_3_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_8_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_8_LFInst_0_n2 ), .B(Input[34]), .ZN(
        Red_Input[32]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_8_LFInst_0_U3  ( .A(Input[35]), .B(
        Input[33]), .ZN(\Red_PlaintextInst_LFInst_8_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_8_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_8_LFInst_1_n2 ), .B(Input[34]), .ZN(
        Red_Input[33]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_8_LFInst_1_U3  ( .A(Input[35]), .B(
        Input[32]), .ZN(\Red_PlaintextInst_LFInst_8_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_8_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_8_LFInst_2_n2 ), .B(Input[33]), .ZN(
        Red_Input[34]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_8_LFInst_2_U3  ( .A(Input[35]), .B(
        Input[32]), .ZN(\Red_PlaintextInst_LFInst_8_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_8_LFInst_3_U4  ( .A(
        \Red_PlaintextInst_LFInst_8_LFInst_3_n2 ), .B(Input[33]), .ZN(
        Red_Input[35]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_8_LFInst_3_U3  ( .A(Input[34]), .B(
        Input[32]), .ZN(\Red_PlaintextInst_LFInst_8_LFInst_3_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_9_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_9_LFInst_0_n2 ), .B(Input[38]), .ZN(
        Red_Input[36]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_9_LFInst_0_U3  ( .A(Input[39]), .B(
        Input[37]), .ZN(\Red_PlaintextInst_LFInst_9_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_9_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_9_LFInst_1_n2 ), .B(Input[38]), .ZN(
        Red_Input[37]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_9_LFInst_1_U3  ( .A(Input[39]), .B(
        Input[36]), .ZN(\Red_PlaintextInst_LFInst_9_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_9_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_9_LFInst_2_n2 ), .B(Input[37]), .ZN(
        Red_Input[38]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_9_LFInst_2_U3  ( .A(Input[39]), .B(
        Input[36]), .ZN(\Red_PlaintextInst_LFInst_9_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_9_LFInst_3_U4  ( .A(
        \Red_PlaintextInst_LFInst_9_LFInst_3_n2 ), .B(Input[37]), .ZN(
        Red_Input[39]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_9_LFInst_3_U3  ( .A(Input[38]), .B(
        Input[36]), .ZN(\Red_PlaintextInst_LFInst_9_LFInst_3_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_10_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_10_LFInst_0_n2 ), .B(Input[42]), .ZN(
        Red_Input[40]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_10_LFInst_0_U3  ( .A(Input[43]), .B(
        Input[41]), .ZN(\Red_PlaintextInst_LFInst_10_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_10_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_10_LFInst_1_n2 ), .B(Input[42]), .ZN(
        Red_Input[41]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_10_LFInst_1_U3  ( .A(Input[43]), .B(
        Input[40]), .ZN(\Red_PlaintextInst_LFInst_10_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_10_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_10_LFInst_2_n2 ), .B(Input[41]), .ZN(
        Red_Input[42]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_10_LFInst_2_U3  ( .A(Input[43]), .B(
        Input[40]), .ZN(\Red_PlaintextInst_LFInst_10_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_10_LFInst_3_U4  ( .A(
        \Red_PlaintextInst_LFInst_10_LFInst_3_n2 ), .B(Input[41]), .ZN(
        Red_Input[43]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_10_LFInst_3_U3  ( .A(Input[42]), .B(
        Input[40]), .ZN(\Red_PlaintextInst_LFInst_10_LFInst_3_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_11_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_11_LFInst_0_n2 ), .B(Input[46]), .ZN(
        Red_Input[44]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_11_LFInst_0_U3  ( .A(Input[47]), .B(
        Input[45]), .ZN(\Red_PlaintextInst_LFInst_11_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_11_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_11_LFInst_1_n2 ), .B(Input[46]), .ZN(
        Red_Input[45]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_11_LFInst_1_U3  ( .A(Input[47]), .B(
        Input[44]), .ZN(\Red_PlaintextInst_LFInst_11_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_11_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_11_LFInst_2_n2 ), .B(Input[45]), .ZN(
        Red_Input[46]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_11_LFInst_2_U3  ( .A(Input[47]), .B(
        Input[44]), .ZN(\Red_PlaintextInst_LFInst_11_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_11_LFInst_3_U4  ( .A(
        \Red_PlaintextInst_LFInst_11_LFInst_3_n2 ), .B(Input[45]), .ZN(
        Red_Input[47]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_11_LFInst_3_U3  ( .A(Input[46]), .B(
        Input[44]), .ZN(\Red_PlaintextInst_LFInst_11_LFInst_3_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_12_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_12_LFInst_0_n2 ), .B(Input[50]), .ZN(
        Red_Input[48]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_12_LFInst_0_U3  ( .A(Input[51]), .B(
        Input[49]), .ZN(\Red_PlaintextInst_LFInst_12_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_12_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_12_LFInst_1_n2 ), .B(Input[50]), .ZN(
        Red_Input[49]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_12_LFInst_1_U3  ( .A(Input[51]), .B(
        Input[48]), .ZN(\Red_PlaintextInst_LFInst_12_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_12_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_12_LFInst_2_n2 ), .B(Input[49]), .ZN(
        Red_Input[50]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_12_LFInst_2_U3  ( .A(Input[51]), .B(
        Input[48]), .ZN(\Red_PlaintextInst_LFInst_12_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_12_LFInst_3_U4  ( .A(
        \Red_PlaintextInst_LFInst_12_LFInst_3_n2 ), .B(Input[49]), .ZN(
        Red_Input[51]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_12_LFInst_3_U3  ( .A(Input[50]), .B(
        Input[48]), .ZN(\Red_PlaintextInst_LFInst_12_LFInst_3_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_13_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_13_LFInst_0_n2 ), .B(Input[54]), .ZN(
        Red_Input[52]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_13_LFInst_0_U3  ( .A(Input[55]), .B(
        Input[53]), .ZN(\Red_PlaintextInst_LFInst_13_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_13_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_13_LFInst_1_n2 ), .B(Input[54]), .ZN(
        Red_Input[53]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_13_LFInst_1_U3  ( .A(Input[55]), .B(
        Input[52]), .ZN(\Red_PlaintextInst_LFInst_13_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_13_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_13_LFInst_2_n2 ), .B(Input[53]), .ZN(
        Red_Input[54]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_13_LFInst_2_U3  ( .A(Input[55]), .B(
        Input[52]), .ZN(\Red_PlaintextInst_LFInst_13_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_13_LFInst_3_U4  ( .A(
        \Red_PlaintextInst_LFInst_13_LFInst_3_n2 ), .B(Input[53]), .ZN(
        Red_Input[55]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_13_LFInst_3_U3  ( .A(Input[54]), .B(
        Input[52]), .ZN(\Red_PlaintextInst_LFInst_13_LFInst_3_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_14_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_14_LFInst_0_n2 ), .B(Input[58]), .ZN(
        Red_Input[56]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_14_LFInst_0_U3  ( .A(Input[59]), .B(
        Input[57]), .ZN(\Red_PlaintextInst_LFInst_14_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_14_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_14_LFInst_1_n2 ), .B(Input[58]), .ZN(
        Red_Input[57]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_14_LFInst_1_U3  ( .A(Input[59]), .B(
        Input[56]), .ZN(\Red_PlaintextInst_LFInst_14_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_14_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_14_LFInst_2_n2 ), .B(Input[57]), .ZN(
        Red_Input[58]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_14_LFInst_2_U3  ( .A(Input[59]), .B(
        Input[56]), .ZN(\Red_PlaintextInst_LFInst_14_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_14_LFInst_3_U4  ( .A(
        \Red_PlaintextInst_LFInst_14_LFInst_3_n2 ), .B(Input[57]), .ZN(
        Red_Input[59]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_14_LFInst_3_U3  ( .A(Input[58]), .B(
        Input[56]), .ZN(\Red_PlaintextInst_LFInst_14_LFInst_3_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_15_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_15_LFInst_0_n2 ), .B(Input[62]), .ZN(
        Red_Input[60]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_15_LFInst_0_U3  ( .A(Input[63]), .B(
        Input[61]), .ZN(\Red_PlaintextInst_LFInst_15_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_15_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_15_LFInst_1_n2 ), .B(Input[62]), .ZN(
        Red_Input[61]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_15_LFInst_1_U3  ( .A(Input[63]), .B(
        Input[60]), .ZN(\Red_PlaintextInst_LFInst_15_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_15_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_15_LFInst_2_n2 ), .B(Input[61]), .ZN(
        Red_Input[62]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_15_LFInst_2_U3  ( .A(Input[63]), .B(
        Input[60]), .ZN(\Red_PlaintextInst_LFInst_15_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_15_LFInst_3_U4  ( .A(
        \Red_PlaintextInst_LFInst_15_LFInst_3_n2 ), .B(Input[61]), .ZN(
        Red_Input[63]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_15_LFInst_3_U3  ( .A(Input[62]), .B(
        Input[60]), .ZN(\Red_PlaintextInst_LFInst_15_LFInst_3_n2 ) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_0_U2  ( .A(\Red_MCInst_XOR_r0_Inst_0_n3 ), 
        .B(Red_MCOutput[0]), .ZN(Red_MCOutput[48]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_0_U1  ( .A(Red_Input[48]), .B(
        Red_MCOutput[16]), .ZN(\Red_MCInst_XOR_r0_Inst_0_n3 ) );
  XOR2_X1 \Red_MCInst_XOR_r1_Inst_0_U1  ( .A(Red_Input[32]), .B(
        Red_MCOutput[0]), .Z(Red_MCOutput[32]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_1_U2  ( .A(\Red_MCInst_XOR_r0_Inst_1_n3 ), 
        .B(Red_MCOutput[1]), .ZN(Red_MCOutput[49]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_1_U1  ( .A(Red_Input[49]), .B(
        Red_MCOutput[17]), .ZN(\Red_MCInst_XOR_r0_Inst_1_n3 ) );
  XOR2_X1 \Red_MCInst_XOR_r1_Inst_1_U1  ( .A(Red_Input[33]), .B(
        Red_MCOutput[1]), .Z(Red_MCOutput[33]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_2_U2  ( .A(\Red_MCInst_XOR_r0_Inst_2_n3 ), 
        .B(Red_MCOutput[2]), .ZN(Red_MCOutput[50]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_2_U1  ( .A(Red_Input[50]), .B(
        Red_MCOutput[18]), .ZN(\Red_MCInst_XOR_r0_Inst_2_n3 ) );
  XOR2_X1 \Red_MCInst_XOR_r1_Inst_2_U1  ( .A(Red_Input[34]), .B(
        Red_MCOutput[2]), .Z(Red_MCOutput[34]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_3_U2  ( .A(\Red_MCInst_XOR_r0_Inst_3_n3 ), 
        .B(Red_MCOutput[3]), .ZN(Red_MCOutput[51]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_3_U1  ( .A(Red_Input[51]), .B(
        Red_MCOutput[19]), .ZN(\Red_MCInst_XOR_r0_Inst_3_n3 ) );
  XOR2_X1 \Red_MCInst_XOR_r1_Inst_3_U1  ( .A(Red_Input[35]), .B(
        Red_MCOutput[3]), .Z(Red_MCOutput[35]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_4_U2  ( .A(\Red_MCInst_XOR_r0_Inst_4_n3 ), 
        .B(Red_MCOutput[4]), .ZN(Red_MCOutput[52]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_4_U1  ( .A(Red_Input[52]), .B(
        Red_MCOutput[20]), .ZN(\Red_MCInst_XOR_r0_Inst_4_n3 ) );
  XOR2_X1 \Red_MCInst_XOR_r1_Inst_4_U1  ( .A(Red_Input[36]), .B(
        Red_MCOutput[4]), .Z(Red_MCOutput[36]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_5_U2  ( .A(\Red_MCInst_XOR_r0_Inst_5_n3 ), 
        .B(Red_MCOutput[5]), .ZN(Red_MCOutput[53]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_5_U1  ( .A(Red_Input[53]), .B(
        Red_MCOutput[21]), .ZN(\Red_MCInst_XOR_r0_Inst_5_n3 ) );
  XOR2_X1 \Red_MCInst_XOR_r1_Inst_5_U1  ( .A(Red_Input[37]), .B(
        Red_MCOutput[5]), .Z(Red_MCOutput[37]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_6_U2  ( .A(\Red_MCInst_XOR_r0_Inst_6_n3 ), 
        .B(Red_MCOutput[6]), .ZN(Red_MCOutput[54]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_6_U1  ( .A(Red_Input[54]), .B(
        Red_MCOutput[22]), .ZN(\Red_MCInst_XOR_r0_Inst_6_n3 ) );
  XOR2_X1 \Red_MCInst_XOR_r1_Inst_6_U1  ( .A(Red_Input[38]), .B(
        Red_MCOutput[6]), .Z(Red_MCOutput[38]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_7_U2  ( .A(\Red_MCInst_XOR_r0_Inst_7_n3 ), 
        .B(Red_MCOutput[7]), .ZN(Red_MCOutput[55]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_7_U1  ( .A(Red_Input[55]), .B(
        Red_MCOutput[23]), .ZN(\Red_MCInst_XOR_r0_Inst_7_n3 ) );
  XOR2_X1 \Red_MCInst_XOR_r1_Inst_7_U1  ( .A(Red_Input[39]), .B(
        Red_MCOutput[7]), .Z(Red_MCOutput[39]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_8_U2  ( .A(\Red_MCInst_XOR_r0_Inst_8_n3 ), 
        .B(Red_MCOutput[8]), .ZN(Red_MCOutput[56]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_8_U1  ( .A(Red_Input[56]), .B(
        Red_MCOutput[24]), .ZN(\Red_MCInst_XOR_r0_Inst_8_n3 ) );
  XOR2_X1 \Red_MCInst_XOR_r1_Inst_8_U1  ( .A(Red_Input[40]), .B(
        Red_MCOutput[8]), .Z(Red_MCOutput[40]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_9_U2  ( .A(\Red_MCInst_XOR_r0_Inst_9_n3 ), 
        .B(Red_MCOutput[9]), .ZN(Red_MCOutput[57]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_9_U1  ( .A(Red_Input[57]), .B(
        Red_MCOutput[25]), .ZN(\Red_MCInst_XOR_r0_Inst_9_n3 ) );
  XOR2_X1 \Red_MCInst_XOR_r1_Inst_9_U1  ( .A(Red_Input[41]), .B(
        Red_MCOutput[9]), .Z(Red_MCOutput[41]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_10_U2  ( .A(\Red_MCInst_XOR_r0_Inst_10_n3 ), 
        .B(Red_MCOutput[10]), .ZN(Red_MCOutput[58]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_10_U1  ( .A(Red_Input[58]), .B(
        Red_MCOutput[26]), .ZN(\Red_MCInst_XOR_r0_Inst_10_n3 ) );
  XOR2_X1 \Red_MCInst_XOR_r1_Inst_10_U1  ( .A(Red_Input[42]), .B(
        Red_MCOutput[10]), .Z(Red_MCOutput[42]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_11_U2  ( .A(\Red_MCInst_XOR_r0_Inst_11_n3 ), 
        .B(Red_MCOutput[11]), .ZN(Red_MCOutput[59]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_11_U1  ( .A(Red_Input[59]), .B(
        Red_MCOutput[27]), .ZN(\Red_MCInst_XOR_r0_Inst_11_n3 ) );
  XOR2_X1 \Red_MCInst_XOR_r1_Inst_11_U1  ( .A(Red_Input[43]), .B(
        Red_MCOutput[11]), .Z(Red_MCOutput[43]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_12_U2  ( .A(\Red_MCInst_XOR_r0_Inst_12_n3 ), 
        .B(Red_MCOutput[12]), .ZN(Red_MCOutput[60]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_12_U1  ( .A(Red_Input[60]), .B(
        Red_MCOutput[28]), .ZN(\Red_MCInst_XOR_r0_Inst_12_n3 ) );
  XOR2_X1 \Red_MCInst_XOR_r1_Inst_12_U1  ( .A(Red_Input[44]), .B(
        Red_MCOutput[12]), .Z(Red_MCOutput[44]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_13_U2  ( .A(\Red_MCInst_XOR_r0_Inst_13_n3 ), 
        .B(Red_MCOutput[13]), .ZN(Red_MCOutput[61]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_13_U1  ( .A(Red_Input[61]), .B(
        Red_MCOutput[29]), .ZN(\Red_MCInst_XOR_r0_Inst_13_n3 ) );
  XOR2_X1 \Red_MCInst_XOR_r1_Inst_13_U1  ( .A(Red_Input[45]), .B(
        Red_MCOutput[13]), .Z(Red_MCOutput[45]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_14_U2  ( .A(\Red_MCInst_XOR_r0_Inst_14_n3 ), 
        .B(Red_MCOutput[14]), .ZN(Red_MCOutput[62]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_14_U1  ( .A(Red_Input[62]), .B(
        Red_MCOutput[30]), .ZN(\Red_MCInst_XOR_r0_Inst_14_n3 ) );
  XOR2_X1 \Red_MCInst_XOR_r1_Inst_14_U1  ( .A(Red_Input[46]), .B(
        Red_MCOutput[14]), .Z(Red_MCOutput[46]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_15_U2  ( .A(\Red_MCInst_XOR_r0_Inst_15_n3 ), 
        .B(Red_MCOutput[15]), .ZN(Red_MCOutput[63]) );
  XNOR2_X1 \Red_MCInst_XOR_r0_Inst_15_U1  ( .A(Red_Input[63]), .B(
        Red_MCOutput[31]), .ZN(\Red_MCInst_XOR_r0_Inst_15_n3 ) );
  XOR2_X1 \Red_MCInst_XOR_r1_Inst_15_U1  ( .A(Red_Input[47]), .B(
        Red_MCOutput[15]), .Z(Red_MCOutput[47]) );
  XOR2_X1 \Red_AddKeyXOR1_XORInst_0_0_U1  ( .A(Red_MCOutput[48]), .B(
        Red_K0[48]), .Z(Red_AddRoundKeyOutput[48]) );
  XOR2_X1 \Red_AddKeyXOR1_XORInst_0_1_U1  ( .A(Red_MCOutput[49]), .B(
        Red_K0[49]), .Z(Red_AddRoundKeyOutput[49]) );
  XOR2_X1 \Red_AddKeyXOR1_XORInst_0_2_U1  ( .A(Red_MCOutput[50]), .B(
        Red_K0[50]), .Z(Red_AddRoundKeyOutput[50]) );
  XOR2_X1 \Red_AddKeyXOR1_XORInst_0_3_U1  ( .A(Red_MCOutput[51]), .B(
        Red_K0[51]), .Z(Red_AddRoundKeyOutput[51]) );
  XOR2_X1 \Red_AddKeyXOR1_XORInst_1_0_U1  ( .A(Red_MCOutput[52]), .B(
        Red_K0[52]), .Z(Red_AddRoundKeyOutput[52]) );
  XOR2_X1 \Red_AddKeyXOR1_XORInst_1_1_U1  ( .A(Red_MCOutput[53]), .B(
        Red_K0[53]), .Z(Red_AddRoundKeyOutput[53]) );
  XOR2_X1 \Red_AddKeyXOR1_XORInst_1_2_U1  ( .A(Red_MCOutput[54]), .B(
        Red_K0[54]), .Z(Red_AddRoundKeyOutput[54]) );
  XOR2_X1 \Red_AddKeyXOR1_XORInst_1_3_U1  ( .A(Red_MCOutput[55]), .B(
        Red_K0[55]), .Z(Red_AddRoundKeyOutput[55]) );
  XOR2_X1 \Red_AddKeyXOR1_XORInst_2_0_U1  ( .A(Red_MCOutput[56]), .B(
        Red_K0[56]), .Z(Red_AddRoundKeyOutput[56]) );
  XOR2_X1 \Red_AddKeyXOR1_XORInst_2_1_U1  ( .A(Red_MCOutput[57]), .B(
        Red_K0[57]), .Z(Red_AddRoundKeyOutput[57]) );
  XOR2_X1 \Red_AddKeyXOR1_XORInst_2_2_U1  ( .A(Red_MCOutput[58]), .B(
        Red_K0[58]), .Z(Red_AddRoundKeyOutput[58]) );
  XOR2_X1 \Red_AddKeyXOR1_XORInst_2_3_U1  ( .A(Red_MCOutput[59]), .B(
        Red_K0[59]), .Z(Red_AddRoundKeyOutput[59]) );
  XOR2_X1 \Red_AddKeyXOR1_XORInst_3_0_U1  ( .A(Red_MCOutput[60]), .B(
        Red_K0[60]), .Z(Red_AddRoundKeyOutput[60]) );
  XOR2_X1 \Red_AddKeyXOR1_XORInst_3_1_U1  ( .A(Red_MCOutput[61]), .B(
        Red_K0[61]), .Z(Red_AddRoundKeyOutput[61]) );
  XOR2_X1 \Red_AddKeyXOR1_XORInst_3_2_U1  ( .A(Red_MCOutput[62]), .B(
        Red_K0[62]), .Z(Red_AddRoundKeyOutput[62]) );
  XOR2_X1 \Red_AddKeyXOR1_XORInst_3_3_U1  ( .A(Red_MCOutput[63]), .B(
        Red_K0[63]), .Z(Red_AddRoundKeyOutput[63]) );
  XOR2_X1 \Red_AddKeyConstXOR_XORInst_0_0_U1  ( .A(Red_K0[40]), .B(
        Red_MCOutput[40]), .Z(Red_AddRoundKeyOutput[40]) );
  XOR2_X1 \Red_AddKeyConstXOR_XORInst_0_1_U1  ( .A(Red_K0[41]), .B(
        Red_MCOutput[41]), .Z(Red_AddRoundKeyOutput[41]) );
  XOR2_X1 \Red_AddKeyConstXOR_XORInst_0_2_U1  ( .A(Red_K0[42]), .B(
        Red_MCOutput[42]), .Z(Red_AddRoundKeyOutput[42]) );
  XOR2_X1 \Red_AddKeyConstXOR_XORInst_0_3_U1  ( .A(Red_K0[43]), .B(
        Red_MCOutput[43]), .Z(Red_AddRoundKeyOutput[43]) );
  XOR2_X1 \Red_AddKeyConstXOR_XORInst_1_0_U1  ( .A(Red_K0[44]), .B(
        Red_MCOutput[44]), .Z(Red_AddRoundKeyOutput[44]) );
  XOR2_X1 \Red_AddKeyConstXOR_XORInst_1_1_U1  ( .A(Red_K0[45]), .B(
        Red_MCOutput[45]), .Z(Red_AddRoundKeyOutput[45]) );
  XOR2_X1 \Red_AddKeyConstXOR_XORInst_1_2_U1  ( .A(Red_K0[46]), .B(
        Red_MCOutput[46]), .Z(Red_AddRoundKeyOutput[46]) );
  XOR2_X1 \Red_AddKeyConstXOR_XORInst_1_3_U1  ( .A(Red_K0[47]), .B(
        Red_MCOutput[47]), .Z(Red_AddRoundKeyOutput[47]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_0_0_U1  ( .A(Red_MCOutput[0]), .B(Red_K0[0]), 
        .Z(Red_AddRoundKeyOutput[0]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_0_1_U1  ( .A(Red_MCOutput[1]), .B(Red_K0[1]), 
        .Z(Red_AddRoundKeyOutput[1]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_0_2_U1  ( .A(Red_MCOutput[2]), .B(Red_K0[2]), 
        .Z(Red_AddRoundKeyOutput[2]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_0_3_U1  ( .A(Red_MCOutput[3]), .B(Red_K0[3]), 
        .Z(Red_AddRoundKeyOutput[3]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_1_0_U1  ( .A(Red_MCOutput[4]), .B(Red_K0[4]), 
        .Z(Red_AddRoundKeyOutput[4]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_1_1_U1  ( .A(Red_MCOutput[5]), .B(Red_K0[5]), 
        .Z(Red_AddRoundKeyOutput[5]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_1_2_U1  ( .A(Red_MCOutput[6]), .B(Red_K0[6]), 
        .Z(Red_AddRoundKeyOutput[6]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_1_3_U1  ( .A(Red_MCOutput[7]), .B(Red_K0[7]), 
        .Z(Red_AddRoundKeyOutput[7]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_2_0_U1  ( .A(Red_MCOutput[8]), .B(Red_K0[8]), 
        .Z(Red_AddRoundKeyOutput[8]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_2_1_U1  ( .A(Red_MCOutput[9]), .B(Red_K0[9]), 
        .Z(Red_AddRoundKeyOutput[9]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_2_2_U1  ( .A(Red_MCOutput[10]), .B(
        Red_K0[10]), .Z(Red_AddRoundKeyOutput[10]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_2_3_U1  ( .A(Red_MCOutput[11]), .B(
        Red_K0[11]), .Z(Red_AddRoundKeyOutput[11]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_3_0_U1  ( .A(Red_MCOutput[12]), .B(
        Red_K0[12]), .Z(Red_AddRoundKeyOutput[12]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_3_1_U1  ( .A(Red_MCOutput[13]), .B(
        Red_K0[13]), .Z(Red_AddRoundKeyOutput[13]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_3_2_U1  ( .A(Red_MCOutput[14]), .B(
        Red_K0[14]), .Z(Red_AddRoundKeyOutput[14]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_3_3_U1  ( .A(Red_MCOutput[15]), .B(
        Red_K0[15]), .Z(Red_AddRoundKeyOutput[15]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_4_0_U1  ( .A(Red_MCOutput[16]), .B(
        Red_K0[16]), .Z(Red_AddRoundKeyOutput[16]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_4_1_U1  ( .A(Red_MCOutput[17]), .B(
        Red_K0[17]), .Z(Red_AddRoundKeyOutput[17]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_4_2_U1  ( .A(Red_MCOutput[18]), .B(
        Red_K0[18]), .Z(Red_AddRoundKeyOutput[18]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_4_3_U1  ( .A(Red_MCOutput[19]), .B(
        Red_K0[19]), .Z(Red_AddRoundKeyOutput[19]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_5_0_U1  ( .A(Red_MCOutput[20]), .B(
        Red_K0[20]), .Z(Red_AddRoundKeyOutput[20]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_5_1_U1  ( .A(Red_MCOutput[21]), .B(
        Red_K0[21]), .Z(Red_AddRoundKeyOutput[21]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_5_2_U1  ( .A(Red_MCOutput[22]), .B(
        Red_K0[22]), .Z(Red_AddRoundKeyOutput[22]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_5_3_U1  ( .A(Red_MCOutput[23]), .B(
        Red_K0[23]), .Z(Red_AddRoundKeyOutput[23]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_6_0_U1  ( .A(Red_MCOutput[24]), .B(
        Red_K0[24]), .Z(Red_AddRoundKeyOutput[24]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_6_1_U1  ( .A(Red_MCOutput[25]), .B(
        Red_K0[25]), .Z(Red_AddRoundKeyOutput[25]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_6_2_U1  ( .A(Red_MCOutput[26]), .B(
        Red_K0[26]), .Z(Red_AddRoundKeyOutput[26]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_6_3_U1  ( .A(Red_MCOutput[27]), .B(
        Red_K0[27]), .Z(Red_AddRoundKeyOutput[27]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_7_0_U1  ( .A(Red_MCOutput[28]), .B(
        Red_K0[28]), .Z(Red_AddRoundKeyOutput[28]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_7_1_U1  ( .A(Red_MCOutput[29]), .B(
        Red_K0[29]), .Z(Red_AddRoundKeyOutput[29]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_7_2_U1  ( .A(Red_MCOutput[30]), .B(
        Red_K0[30]), .Z(Red_AddRoundKeyOutput[30]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_7_3_U1  ( .A(Red_MCOutput[31]), .B(
        Red_K0[31]), .Z(Red_AddRoundKeyOutput[31]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_8_0_U1  ( .A(Red_MCOutput[32]), .B(
        Red_K0[32]), .Z(Red_AddRoundKeyOutput[32]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_8_1_U1  ( .A(Red_MCOutput[33]), .B(
        Red_K0[33]), .Z(Red_AddRoundKeyOutput[33]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_8_2_U1  ( .A(Red_MCOutput[34]), .B(
        Red_K0[34]), .Z(Red_AddRoundKeyOutput[34]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_8_3_U1  ( .A(Red_MCOutput[35]), .B(
        Red_K0[35]), .Z(Red_AddRoundKeyOutput[35]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_9_0_U1  ( .A(Red_MCOutput[36]), .B(
        Red_K0[36]), .Z(Red_AddRoundKeyOutput[36]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_9_1_U1  ( .A(Red_MCOutput[37]), .B(
        Red_K0[37]), .Z(Red_AddRoundKeyOutput[37]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_9_2_U1  ( .A(Red_MCOutput[38]), .B(
        Red_K0[38]), .Z(Red_AddRoundKeyOutput[38]) );
  XOR2_X1 \Red_AddKeyXOR2_XORInst_9_3_U1  ( .A(Red_MCOutput[39]), .B(
        Red_K0[39]), .Z(Red_AddRoundKeyOutput[39]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[0]  ( .D(Red_AddRoundKeyOutput[0]), 
        .CK(clk), .Q(Red_StateRegOutput[0]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[1]  ( .D(Red_AddRoundKeyOutput[1]), 
        .CK(clk), .Q(Red_StateRegOutput[1]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[2]  ( .D(Red_AddRoundKeyOutput[2]), 
        .CK(clk), .Q(Red_StateRegOutput[2]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[3]  ( .D(Red_AddRoundKeyOutput[3]), 
        .CK(clk), .Q(Red_StateRegOutput[3]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[4]  ( .D(Red_AddRoundKeyOutput[4]), 
        .CK(clk), .Q(Red_StateRegOutput[4]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[5]  ( .D(Red_AddRoundKeyOutput[5]), 
        .CK(clk), .Q(Red_StateRegOutput[5]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[6]  ( .D(Red_AddRoundKeyOutput[6]), 
        .CK(clk), .Q(Red_StateRegOutput[6]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[7]  ( .D(Red_AddRoundKeyOutput[7]), 
        .CK(clk), .Q(Red_StateRegOutput[7]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[8]  ( .D(Red_AddRoundKeyOutput[8]), 
        .CK(clk), .Q(Red_StateRegOutput[8]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[9]  ( .D(Red_AddRoundKeyOutput[9]), 
        .CK(clk), .Q(Red_StateRegOutput[9]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[10]  ( .D(Red_AddRoundKeyOutput[10]), .CK(clk), .Q(Red_StateRegOutput[10]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[11]  ( .D(Red_AddRoundKeyOutput[11]), .CK(clk), .Q(Red_StateRegOutput[11]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[12]  ( .D(Red_AddRoundKeyOutput[12]), .CK(clk), .Q(Red_StateRegOutput[12]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[13]  ( .D(Red_AddRoundKeyOutput[13]), .CK(clk), .Q(Red_StateRegOutput[13]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[14]  ( .D(Red_AddRoundKeyOutput[14]), .CK(clk), .Q(Red_StateRegOutput[14]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[15]  ( .D(Red_AddRoundKeyOutput[15]), .CK(clk), .Q(Red_StateRegOutput[15]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[16]  ( .D(Red_AddRoundKeyOutput[16]), .CK(clk), .Q(Red_StateRegOutput[16]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[17]  ( .D(Red_AddRoundKeyOutput[17]), .CK(clk), .Q(Red_StateRegOutput[17]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[18]  ( .D(Red_AddRoundKeyOutput[18]), .CK(clk), .Q(Red_StateRegOutput[18]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[19]  ( .D(Red_AddRoundKeyOutput[19]), .CK(clk), .Q(Red_StateRegOutput[19]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[20]  ( .D(Red_AddRoundKeyOutput[20]), .CK(clk), .Q(Red_StateRegOutput[20]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[21]  ( .D(Red_AddRoundKeyOutput[21]), .CK(clk), .Q(Red_StateRegOutput[21]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[22]  ( .D(Red_AddRoundKeyOutput[22]), .CK(clk), .Q(Red_StateRegOutput[22]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[23]  ( .D(Red_AddRoundKeyOutput[23]), .CK(clk), .Q(Red_StateRegOutput[23]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[24]  ( .D(Red_AddRoundKeyOutput[24]), .CK(clk), .Q(Red_StateRegOutput[24]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[25]  ( .D(Red_AddRoundKeyOutput[25]), .CK(clk), .Q(Red_StateRegOutput[25]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[26]  ( .D(Red_AddRoundKeyOutput[26]), .CK(clk), .Q(Red_StateRegOutput[26]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[27]  ( .D(Red_AddRoundKeyOutput[27]), .CK(clk), .Q(Red_StateRegOutput[27]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[28]  ( .D(Red_AddRoundKeyOutput[28]), .CK(clk), .Q(Red_StateRegOutput[28]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[29]  ( .D(Red_AddRoundKeyOutput[29]), .CK(clk), .Q(Red_StateRegOutput[29]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[30]  ( .D(Red_AddRoundKeyOutput[30]), .CK(clk), .Q(Red_StateRegOutput[30]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[31]  ( .D(Red_AddRoundKeyOutput[31]), .CK(clk), .Q(Red_StateRegOutput[31]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[32]  ( .D(Red_AddRoundKeyOutput[32]), .CK(clk), .Q(Red_StateRegOutput[32]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[33]  ( .D(Red_AddRoundKeyOutput[33]), .CK(clk), .Q(Red_StateRegOutput[33]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[34]  ( .D(Red_AddRoundKeyOutput[34]), .CK(clk), .Q(Red_StateRegOutput[34]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[35]  ( .D(Red_AddRoundKeyOutput[35]), .CK(clk), .Q(Red_StateRegOutput[35]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[36]  ( .D(Red_AddRoundKeyOutput[36]), .CK(clk), .Q(Red_StateRegOutput[36]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[37]  ( .D(Red_AddRoundKeyOutput[37]), .CK(clk), .Q(Red_StateRegOutput[37]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[38]  ( .D(Red_AddRoundKeyOutput[38]), .CK(clk), .Q(Red_StateRegOutput[38]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[39]  ( .D(Red_AddRoundKeyOutput[39]), .CK(clk), .Q(Red_StateRegOutput[39]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[40]  ( .D(Red_AddRoundKeyOutput[40]), .CK(clk), .Q(Red_StateRegOutput[40]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[41]  ( .D(Red_AddRoundKeyOutput[41]), .CK(clk), .Q(Red_StateRegOutput[41]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[42]  ( .D(Red_AddRoundKeyOutput[42]), .CK(clk), .Q(Red_StateRegOutput[42]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[43]  ( .D(Red_AddRoundKeyOutput[43]), .CK(clk), .Q(Red_StateRegOutput[43]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[44]  ( .D(Red_AddRoundKeyOutput[44]), .CK(clk), .Q(Red_StateRegOutput[44]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[45]  ( .D(Red_AddRoundKeyOutput[45]), .CK(clk), .Q(Red_StateRegOutput[45]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[46]  ( .D(Red_AddRoundKeyOutput[46]), .CK(clk), .Q(Red_StateRegOutput[46]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[47]  ( .D(Red_AddRoundKeyOutput[47]), .CK(clk), .Q(Red_StateRegOutput[47]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[48]  ( .D(Red_AddRoundKeyOutput[48]), .CK(clk), .Q(Red_StateRegOutput[48]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[49]  ( .D(Red_AddRoundKeyOutput[49]), .CK(clk), .Q(Red_StateRegOutput[49]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[50]  ( .D(Red_AddRoundKeyOutput[50]), .CK(clk), .Q(Red_StateRegOutput[50]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[51]  ( .D(Red_AddRoundKeyOutput[51]), .CK(clk), .Q(Red_StateRegOutput[51]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[52]  ( .D(Red_AddRoundKeyOutput[52]), .CK(clk), .Q(Red_StateRegOutput[52]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[53]  ( .D(Red_AddRoundKeyOutput[53]), .CK(clk), .Q(Red_StateRegOutput[53]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[54]  ( .D(Red_AddRoundKeyOutput[54]), .CK(clk), .Q(Red_StateRegOutput[54]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[55]  ( .D(Red_AddRoundKeyOutput[55]), .CK(clk), .Q(Red_StateRegOutput[55]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[56]  ( .D(Red_AddRoundKeyOutput[56]), .CK(clk), .Q(Red_StateRegOutput[56]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[57]  ( .D(Red_AddRoundKeyOutput[57]), .CK(clk), .Q(Red_StateRegOutput[57]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[58]  ( .D(Red_AddRoundKeyOutput[58]), .CK(clk), .Q(Red_StateRegOutput[58]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[59]  ( .D(Red_AddRoundKeyOutput[59]), .CK(clk), .Q(Red_StateRegOutput[59]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[60]  ( .D(Red_AddRoundKeyOutput[60]), .CK(clk), .Q(Red_StateRegOutput[60]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[61]  ( .D(Red_AddRoundKeyOutput[61]), .CK(clk), .Q(Red_StateRegOutput[61]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[62]  ( .D(Red_AddRoundKeyOutput[62]), .CK(clk), .Q(Red_StateRegOutput[62]) );
  DFF_X1 \Red_StateReg_s_current_state_reg[63]  ( .D(Red_AddRoundKeyOutput[63]), .CK(clk), .Q(Red_StateRegOutput[63]) );
  NAND2_X1 \Red_SubCellInst_LFInst_0_LFInst_0_U10  ( .A1(
        \Red_SubCellInst_LFInst_0_LFInst_0_n14 ), .A2(
        \Red_SubCellInst_LFInst_0_LFInst_0_n13 ), .ZN(Red_MCOutput2[0]) );
  NAND2_X1 \Red_SubCellInst_LFInst_0_LFInst_0_U9  ( .A1(PermutationOutput[0]), 
        .A2(\Red_SubCellInst_LFInst_0_LFInst_0_n12 ), .ZN(
        \Red_SubCellInst_LFInst_0_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_0_LFInst_0_U8  ( .A1(
        \Red_SubCellInst_LFInst_0_LFInst_0_n11 ), .A2(PermutationOutput[2]), 
        .ZN(\Red_SubCellInst_LFInst_0_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_0_LFInst_0_U7  ( .A(
        \Red_SubCellInst_LFInst_0_LFInst_0_n10 ), .B(
        \Red_SubCellInst_LFInst_0_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst_LFInst_0_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_0_LFInst_0_U6  ( .A1(PermutationOutput[3]), 
        .A2(\Red_SubCellInst_LFInst_0_LFInst_0_n11 ), .ZN(
        \Red_SubCellInst_LFInst_0_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst_LFInst_0_LFInst_0_U5  ( .A(PermutationOutput[1]), 
        .ZN(\Red_SubCellInst_LFInst_0_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_0_LFInst_0_U4  ( .A1(PermutationOutput[2]), 
        .A2(\Red_SubCellInst_LFInst_0_LFInst_0_n8 ), .ZN(
        \Red_SubCellInst_LFInst_0_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst_LFInst_0_LFInst_0_U3  ( .A(PermutationOutput[0]), 
        .ZN(\Red_SubCellInst_LFInst_0_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_0_LFInst_1_U8  ( .A1(
        \Red_SubCellInst_LFInst_0_LFInst_1_n15 ), .A2(
        \Red_SubCellInst_LFInst_0_LFInst_1_n14 ), .ZN(Red_MCOutput2[1]) );
  NAND2_X1 \Red_SubCellInst_LFInst_0_LFInst_1_U7  ( .A1(
        \Red_SubCellInst_LFInst_0_LFInst_1_n13 ), .A2(PermutationOutput[1]), 
        .ZN(\Red_SubCellInst_LFInst_0_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_0_LFInst_1_U6  ( .A1(
        \Red_SubCellInst_LFInst_0_LFInst_1_n12 ), .A2(PermutationOutput[0]), 
        .ZN(\Red_SubCellInst_LFInst_0_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_0_LFInst_1_U5  ( .A1(PermutationOutput[3]), 
        .A2(PermutationOutput[2]), .ZN(\Red_SubCellInst_LFInst_0_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst_LFInst_0_LFInst_1_U4  ( .A1(PermutationOutput[2]), 
        .A2(\Red_SubCellInst_LFInst_0_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst_LFInst_0_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_0_LFInst_1_U3  ( .A(PermutationOutput[0]), 
        .B(PermutationOutput[3]), .ZN(\Red_SubCellInst_LFInst_0_LFInst_1_n11 )
         );
  NOR2_X1 \Red_SubCellInst_LFInst_0_LFInst_2_U10  ( .A1(
        \Red_SubCellInst_LFInst_0_LFInst_2_n19 ), .A2(
        \Red_SubCellInst_LFInst_0_LFInst_2_n18 ), .ZN(Red_MCOutput2[2]) );
  AND2_X1 \Red_SubCellInst_LFInst_0_LFInst_2_U9  ( .A1(
        \Red_SubCellInst_LFInst_0_LFInst_2_n17 ), .A2(PermutationOutput[0]), 
        .ZN(\Red_SubCellInst_LFInst_0_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_0_LFInst_2_U8  ( .A1(PermutationOutput[2]), 
        .A2(PermutationOutput[1]), .ZN(\Red_SubCellInst_LFInst_0_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_0_LFInst_2_U7  ( .A(
        \Red_SubCellInst_LFInst_0_LFInst_2_n16 ), .B(
        \Red_SubCellInst_LFInst_0_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst_LFInst_0_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_0_LFInst_2_U6  ( .A1(PermutationOutput[3]), 
        .A2(\Red_SubCellInst_LFInst_0_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst_LFInst_0_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst_LFInst_0_LFInst_2_U5  ( .A(PermutationOutput[1]), 
        .ZN(\Red_SubCellInst_LFInst_0_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_0_LFInst_2_U4  ( .A1(PermutationOutput[2]), 
        .A2(\Red_SubCellInst_LFInst_0_LFInst_2_n13 ), .ZN(
        \Red_SubCellInst_LFInst_0_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst_LFInst_0_LFInst_2_U3  ( .A(PermutationOutput[0]), 
        .ZN(\Red_SubCellInst_LFInst_0_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_0_LFInst_3_U6  ( .A(PermutationOutput[1]), 
        .B(\Red_SubCellInst_LFInst_0_LFInst_3_n8 ), .ZN(Red_MCOutput2[3]) );
  NOR2_X1 \Red_SubCellInst_LFInst_0_LFInst_3_U5  ( .A1(
        \Red_SubCellInst_LFInst_0_LFInst_3_n7 ), .A2(
        \Red_SubCellInst_LFInst_0_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst_LFInst_0_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_0_LFInst_3_U4  ( .A1(PermutationOutput[2]), 
        .A2(PermutationOutput[3]), .ZN(\Red_SubCellInst_LFInst_0_LFInst_3_n6 )
         );
  AND2_X1 \Red_SubCellInst_LFInst_0_LFInst_3_U3  ( .A1(PermutationOutput[3]), 
        .A2(PermutationOutput[0]), .ZN(\Red_SubCellInst_LFInst_0_LFInst_3_n7 )
         );
  NAND2_X1 \Red_SubCellInst_LFInst_1_LFInst_0_U10  ( .A1(
        \Red_SubCellInst_LFInst_1_LFInst_0_n14 ), .A2(
        \Red_SubCellInst_LFInst_1_LFInst_0_n13 ), .ZN(Red_MCOutput2[4]) );
  NAND2_X1 \Red_SubCellInst_LFInst_1_LFInst_0_U9  ( .A1(PermutationOutput[4]), 
        .A2(\Red_SubCellInst_LFInst_1_LFInst_0_n12 ), .ZN(
        \Red_SubCellInst_LFInst_1_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_1_LFInst_0_U8  ( .A1(
        \Red_SubCellInst_LFInst_1_LFInst_0_n11 ), .A2(PermutationOutput[6]), 
        .ZN(\Red_SubCellInst_LFInst_1_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_1_LFInst_0_U7  ( .A(
        \Red_SubCellInst_LFInst_1_LFInst_0_n10 ), .B(
        \Red_SubCellInst_LFInst_1_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst_LFInst_1_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_1_LFInst_0_U6  ( .A1(PermutationOutput[7]), 
        .A2(\Red_SubCellInst_LFInst_1_LFInst_0_n11 ), .ZN(
        \Red_SubCellInst_LFInst_1_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst_LFInst_1_LFInst_0_U5  ( .A(PermutationOutput[5]), 
        .ZN(\Red_SubCellInst_LFInst_1_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_1_LFInst_0_U4  ( .A1(PermutationOutput[6]), 
        .A2(\Red_SubCellInst_LFInst_1_LFInst_0_n8 ), .ZN(
        \Red_SubCellInst_LFInst_1_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst_LFInst_1_LFInst_0_U3  ( .A(PermutationOutput[4]), 
        .ZN(\Red_SubCellInst_LFInst_1_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_1_LFInst_1_U8  ( .A1(
        \Red_SubCellInst_LFInst_1_LFInst_1_n15 ), .A2(
        \Red_SubCellInst_LFInst_1_LFInst_1_n14 ), .ZN(Red_MCOutput2[5]) );
  NAND2_X1 \Red_SubCellInst_LFInst_1_LFInst_1_U7  ( .A1(
        \Red_SubCellInst_LFInst_1_LFInst_1_n13 ), .A2(PermutationOutput[5]), 
        .ZN(\Red_SubCellInst_LFInst_1_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_1_LFInst_1_U6  ( .A1(
        \Red_SubCellInst_LFInst_1_LFInst_1_n12 ), .A2(PermutationOutput[4]), 
        .ZN(\Red_SubCellInst_LFInst_1_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_1_LFInst_1_U5  ( .A1(PermutationOutput[7]), 
        .A2(PermutationOutput[6]), .ZN(\Red_SubCellInst_LFInst_1_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst_LFInst_1_LFInst_1_U4  ( .A1(PermutationOutput[6]), 
        .A2(\Red_SubCellInst_LFInst_1_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst_LFInst_1_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_1_LFInst_1_U3  ( .A(PermutationOutput[4]), 
        .B(PermutationOutput[7]), .ZN(\Red_SubCellInst_LFInst_1_LFInst_1_n11 )
         );
  NOR2_X1 \Red_SubCellInst_LFInst_1_LFInst_2_U10  ( .A1(
        \Red_SubCellInst_LFInst_1_LFInst_2_n19 ), .A2(
        \Red_SubCellInst_LFInst_1_LFInst_2_n18 ), .ZN(Red_MCOutput2[6]) );
  AND2_X1 \Red_SubCellInst_LFInst_1_LFInst_2_U9  ( .A1(
        \Red_SubCellInst_LFInst_1_LFInst_2_n17 ), .A2(PermutationOutput[4]), 
        .ZN(\Red_SubCellInst_LFInst_1_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_1_LFInst_2_U8  ( .A1(PermutationOutput[6]), 
        .A2(PermutationOutput[5]), .ZN(\Red_SubCellInst_LFInst_1_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_1_LFInst_2_U7  ( .A(
        \Red_SubCellInst_LFInst_1_LFInst_2_n16 ), .B(
        \Red_SubCellInst_LFInst_1_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst_LFInst_1_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_1_LFInst_2_U6  ( .A1(PermutationOutput[7]), 
        .A2(\Red_SubCellInst_LFInst_1_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst_LFInst_1_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst_LFInst_1_LFInst_2_U5  ( .A(PermutationOutput[5]), 
        .ZN(\Red_SubCellInst_LFInst_1_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_1_LFInst_2_U4  ( .A1(PermutationOutput[6]), 
        .A2(\Red_SubCellInst_LFInst_1_LFInst_2_n13 ), .ZN(
        \Red_SubCellInst_LFInst_1_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst_LFInst_1_LFInst_2_U3  ( .A(PermutationOutput[4]), 
        .ZN(\Red_SubCellInst_LFInst_1_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_1_LFInst_3_U6  ( .A(PermutationOutput[5]), 
        .B(\Red_SubCellInst_LFInst_1_LFInst_3_n8 ), .ZN(Red_MCOutput2[7]) );
  NOR2_X1 \Red_SubCellInst_LFInst_1_LFInst_3_U5  ( .A1(
        \Red_SubCellInst_LFInst_1_LFInst_3_n7 ), .A2(
        \Red_SubCellInst_LFInst_1_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst_LFInst_1_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_1_LFInst_3_U4  ( .A1(PermutationOutput[6]), 
        .A2(PermutationOutput[7]), .ZN(\Red_SubCellInst_LFInst_1_LFInst_3_n6 )
         );
  AND2_X1 \Red_SubCellInst_LFInst_1_LFInst_3_U3  ( .A1(PermutationOutput[7]), 
        .A2(PermutationOutput[4]), .ZN(\Red_SubCellInst_LFInst_1_LFInst_3_n7 )
         );
  NAND2_X1 \Red_SubCellInst_LFInst_2_LFInst_0_U10  ( .A1(
        \Red_SubCellInst_LFInst_2_LFInst_0_n14 ), .A2(
        \Red_SubCellInst_LFInst_2_LFInst_0_n13 ), .ZN(Red_MCOutput2[8]) );
  NAND2_X1 \Red_SubCellInst_LFInst_2_LFInst_0_U9  ( .A1(PermutationOutput[8]), 
        .A2(\Red_SubCellInst_LFInst_2_LFInst_0_n12 ), .ZN(
        \Red_SubCellInst_LFInst_2_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_2_LFInst_0_U8  ( .A1(
        \Red_SubCellInst_LFInst_2_LFInst_0_n11 ), .A2(PermutationOutput[10]), 
        .ZN(\Red_SubCellInst_LFInst_2_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_2_LFInst_0_U7  ( .A(
        \Red_SubCellInst_LFInst_2_LFInst_0_n10 ), .B(
        \Red_SubCellInst_LFInst_2_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst_LFInst_2_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_2_LFInst_0_U6  ( .A1(PermutationOutput[11]), 
        .A2(\Red_SubCellInst_LFInst_2_LFInst_0_n11 ), .ZN(
        \Red_SubCellInst_LFInst_2_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst_LFInst_2_LFInst_0_U5  ( .A(PermutationOutput[9]), 
        .ZN(\Red_SubCellInst_LFInst_2_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_2_LFInst_0_U4  ( .A1(PermutationOutput[10]), 
        .A2(\Red_SubCellInst_LFInst_2_LFInst_0_n8 ), .ZN(
        \Red_SubCellInst_LFInst_2_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst_LFInst_2_LFInst_0_U3  ( .A(PermutationOutput[8]), 
        .ZN(\Red_SubCellInst_LFInst_2_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_2_LFInst_1_U8  ( .A1(
        \Red_SubCellInst_LFInst_2_LFInst_1_n15 ), .A2(
        \Red_SubCellInst_LFInst_2_LFInst_1_n14 ), .ZN(Red_MCOutput2[9]) );
  NAND2_X1 \Red_SubCellInst_LFInst_2_LFInst_1_U7  ( .A1(
        \Red_SubCellInst_LFInst_2_LFInst_1_n13 ), .A2(PermutationOutput[9]), 
        .ZN(\Red_SubCellInst_LFInst_2_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_2_LFInst_1_U6  ( .A1(
        \Red_SubCellInst_LFInst_2_LFInst_1_n12 ), .A2(PermutationOutput[8]), 
        .ZN(\Red_SubCellInst_LFInst_2_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_2_LFInst_1_U5  ( .A1(PermutationOutput[11]), 
        .A2(PermutationOutput[10]), .ZN(
        \Red_SubCellInst_LFInst_2_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst_LFInst_2_LFInst_1_U4  ( .A1(PermutationOutput[10]), 
        .A2(\Red_SubCellInst_LFInst_2_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst_LFInst_2_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_2_LFInst_1_U3  ( .A(PermutationOutput[8]), 
        .B(PermutationOutput[11]), .ZN(\Red_SubCellInst_LFInst_2_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_2_LFInst_2_U10  ( .A1(
        \Red_SubCellInst_LFInst_2_LFInst_2_n19 ), .A2(
        \Red_SubCellInst_LFInst_2_LFInst_2_n18 ), .ZN(Red_MCOutput2[10]) );
  AND2_X1 \Red_SubCellInst_LFInst_2_LFInst_2_U9  ( .A1(
        \Red_SubCellInst_LFInst_2_LFInst_2_n17 ), .A2(PermutationOutput[8]), 
        .ZN(\Red_SubCellInst_LFInst_2_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_2_LFInst_2_U8  ( .A1(PermutationOutput[10]), 
        .A2(PermutationOutput[9]), .ZN(\Red_SubCellInst_LFInst_2_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_2_LFInst_2_U7  ( .A(
        \Red_SubCellInst_LFInst_2_LFInst_2_n16 ), .B(
        \Red_SubCellInst_LFInst_2_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst_LFInst_2_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_2_LFInst_2_U6  ( .A1(PermutationOutput[11]), 
        .A2(\Red_SubCellInst_LFInst_2_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst_LFInst_2_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst_LFInst_2_LFInst_2_U5  ( .A(PermutationOutput[9]), 
        .ZN(\Red_SubCellInst_LFInst_2_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_2_LFInst_2_U4  ( .A1(PermutationOutput[10]), 
        .A2(\Red_SubCellInst_LFInst_2_LFInst_2_n13 ), .ZN(
        \Red_SubCellInst_LFInst_2_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst_LFInst_2_LFInst_2_U3  ( .A(PermutationOutput[8]), 
        .ZN(\Red_SubCellInst_LFInst_2_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_2_LFInst_3_U6  ( .A(PermutationOutput[9]), 
        .B(\Red_SubCellInst_LFInst_2_LFInst_3_n8 ), .ZN(Red_MCOutput2[11]) );
  NOR2_X1 \Red_SubCellInst_LFInst_2_LFInst_3_U5  ( .A1(
        \Red_SubCellInst_LFInst_2_LFInst_3_n7 ), .A2(
        \Red_SubCellInst_LFInst_2_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst_LFInst_2_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_2_LFInst_3_U4  ( .A1(PermutationOutput[10]), 
        .A2(PermutationOutput[11]), .ZN(\Red_SubCellInst_LFInst_2_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst_LFInst_2_LFInst_3_U3  ( .A1(PermutationOutput[11]), 
        .A2(PermutationOutput[8]), .ZN(\Red_SubCellInst_LFInst_2_LFInst_3_n7 )
         );
  NAND2_X1 \Red_SubCellInst_LFInst_3_LFInst_0_U10  ( .A1(
        \Red_SubCellInst_LFInst_3_LFInst_0_n14 ), .A2(
        \Red_SubCellInst_LFInst_3_LFInst_0_n13 ), .ZN(Red_MCOutput2[12]) );
  NAND2_X1 \Red_SubCellInst_LFInst_3_LFInst_0_U9  ( .A1(PermutationOutput[12]), 
        .A2(\Red_SubCellInst_LFInst_3_LFInst_0_n12 ), .ZN(
        \Red_SubCellInst_LFInst_3_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_3_LFInst_0_U8  ( .A1(
        \Red_SubCellInst_LFInst_3_LFInst_0_n11 ), .A2(PermutationOutput[14]), 
        .ZN(\Red_SubCellInst_LFInst_3_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_3_LFInst_0_U7  ( .A(
        \Red_SubCellInst_LFInst_3_LFInst_0_n10 ), .B(
        \Red_SubCellInst_LFInst_3_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst_LFInst_3_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_3_LFInst_0_U6  ( .A1(PermutationOutput[15]), 
        .A2(\Red_SubCellInst_LFInst_3_LFInst_0_n11 ), .ZN(
        \Red_SubCellInst_LFInst_3_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst_LFInst_3_LFInst_0_U5  ( .A(PermutationOutput[13]), 
        .ZN(\Red_SubCellInst_LFInst_3_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_3_LFInst_0_U4  ( .A1(PermutationOutput[14]), 
        .A2(\Red_SubCellInst_LFInst_3_LFInst_0_n8 ), .ZN(
        \Red_SubCellInst_LFInst_3_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst_LFInst_3_LFInst_0_U3  ( .A(PermutationOutput[12]), 
        .ZN(\Red_SubCellInst_LFInst_3_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_3_LFInst_1_U8  ( .A1(
        \Red_SubCellInst_LFInst_3_LFInst_1_n15 ), .A2(
        \Red_SubCellInst_LFInst_3_LFInst_1_n14 ), .ZN(Red_MCOutput2[13]) );
  NAND2_X1 \Red_SubCellInst_LFInst_3_LFInst_1_U7  ( .A1(
        \Red_SubCellInst_LFInst_3_LFInst_1_n13 ), .A2(PermutationOutput[13]), 
        .ZN(\Red_SubCellInst_LFInst_3_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_3_LFInst_1_U6  ( .A1(
        \Red_SubCellInst_LFInst_3_LFInst_1_n12 ), .A2(PermutationOutput[12]), 
        .ZN(\Red_SubCellInst_LFInst_3_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_3_LFInst_1_U5  ( .A1(PermutationOutput[15]), 
        .A2(PermutationOutput[14]), .ZN(
        \Red_SubCellInst_LFInst_3_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst_LFInst_3_LFInst_1_U4  ( .A1(PermutationOutput[14]), 
        .A2(\Red_SubCellInst_LFInst_3_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst_LFInst_3_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_3_LFInst_1_U3  ( .A(PermutationOutput[12]), 
        .B(PermutationOutput[15]), .ZN(\Red_SubCellInst_LFInst_3_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_3_LFInst_2_U10  ( .A1(
        \Red_SubCellInst_LFInst_3_LFInst_2_n19 ), .A2(
        \Red_SubCellInst_LFInst_3_LFInst_2_n18 ), .ZN(Red_MCOutput2[14]) );
  AND2_X1 \Red_SubCellInst_LFInst_3_LFInst_2_U9  ( .A1(
        \Red_SubCellInst_LFInst_3_LFInst_2_n17 ), .A2(PermutationOutput[12]), 
        .ZN(\Red_SubCellInst_LFInst_3_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_3_LFInst_2_U8  ( .A1(PermutationOutput[14]), 
        .A2(PermutationOutput[13]), .ZN(
        \Red_SubCellInst_LFInst_3_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_3_LFInst_2_U7  ( .A(
        \Red_SubCellInst_LFInst_3_LFInst_2_n16 ), .B(
        \Red_SubCellInst_LFInst_3_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst_LFInst_3_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_3_LFInst_2_U6  ( .A1(PermutationOutput[15]), 
        .A2(\Red_SubCellInst_LFInst_3_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst_LFInst_3_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst_LFInst_3_LFInst_2_U5  ( .A(PermutationOutput[13]), 
        .ZN(\Red_SubCellInst_LFInst_3_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_3_LFInst_2_U4  ( .A1(PermutationOutput[14]), 
        .A2(\Red_SubCellInst_LFInst_3_LFInst_2_n13 ), .ZN(
        \Red_SubCellInst_LFInst_3_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst_LFInst_3_LFInst_2_U3  ( .A(PermutationOutput[12]), 
        .ZN(\Red_SubCellInst_LFInst_3_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_3_LFInst_3_U6  ( .A(PermutationOutput[13]), 
        .B(\Red_SubCellInst_LFInst_3_LFInst_3_n8 ), .ZN(Red_MCOutput2[15]) );
  NOR2_X1 \Red_SubCellInst_LFInst_3_LFInst_3_U5  ( .A1(
        \Red_SubCellInst_LFInst_3_LFInst_3_n7 ), .A2(
        \Red_SubCellInst_LFInst_3_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst_LFInst_3_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_3_LFInst_3_U4  ( .A1(PermutationOutput[14]), 
        .A2(PermutationOutput[15]), .ZN(\Red_SubCellInst_LFInst_3_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst_LFInst_3_LFInst_3_U3  ( .A1(PermutationOutput[15]), 
        .A2(PermutationOutput[12]), .ZN(\Red_SubCellInst_LFInst_3_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_4_LFInst_0_U10  ( .A1(
        \Red_SubCellInst_LFInst_4_LFInst_0_n14 ), .A2(
        \Red_SubCellInst_LFInst_4_LFInst_0_n13 ), .ZN(Red_MCOutput2[16]) );
  NAND2_X1 \Red_SubCellInst_LFInst_4_LFInst_0_U9  ( .A1(PermutationOutput[16]), 
        .A2(\Red_SubCellInst_LFInst_4_LFInst_0_n12 ), .ZN(
        \Red_SubCellInst_LFInst_4_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_4_LFInst_0_U8  ( .A1(
        \Red_SubCellInst_LFInst_4_LFInst_0_n11 ), .A2(PermutationOutput[18]), 
        .ZN(\Red_SubCellInst_LFInst_4_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_4_LFInst_0_U7  ( .A(
        \Red_SubCellInst_LFInst_4_LFInst_0_n10 ), .B(
        \Red_SubCellInst_LFInst_4_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst_LFInst_4_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_4_LFInst_0_U6  ( .A1(PermutationOutput[19]), 
        .A2(\Red_SubCellInst_LFInst_4_LFInst_0_n11 ), .ZN(
        \Red_SubCellInst_LFInst_4_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst_LFInst_4_LFInst_0_U5  ( .A(PermutationOutput[17]), 
        .ZN(\Red_SubCellInst_LFInst_4_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_4_LFInst_0_U4  ( .A1(PermutationOutput[18]), 
        .A2(\Red_SubCellInst_LFInst_4_LFInst_0_n8 ), .ZN(
        \Red_SubCellInst_LFInst_4_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst_LFInst_4_LFInst_0_U3  ( .A(PermutationOutput[16]), 
        .ZN(\Red_SubCellInst_LFInst_4_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_4_LFInst_1_U8  ( .A1(
        \Red_SubCellInst_LFInst_4_LFInst_1_n15 ), .A2(
        \Red_SubCellInst_LFInst_4_LFInst_1_n14 ), .ZN(Red_MCOutput2[17]) );
  NAND2_X1 \Red_SubCellInst_LFInst_4_LFInst_1_U7  ( .A1(
        \Red_SubCellInst_LFInst_4_LFInst_1_n13 ), .A2(PermutationOutput[17]), 
        .ZN(\Red_SubCellInst_LFInst_4_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_4_LFInst_1_U6  ( .A1(
        \Red_SubCellInst_LFInst_4_LFInst_1_n12 ), .A2(PermutationOutput[16]), 
        .ZN(\Red_SubCellInst_LFInst_4_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_4_LFInst_1_U5  ( .A1(PermutationOutput[19]), 
        .A2(PermutationOutput[18]), .ZN(
        \Red_SubCellInst_LFInst_4_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst_LFInst_4_LFInst_1_U4  ( .A1(PermutationOutput[18]), 
        .A2(\Red_SubCellInst_LFInst_4_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst_LFInst_4_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_4_LFInst_1_U3  ( .A(PermutationOutput[16]), 
        .B(PermutationOutput[19]), .ZN(\Red_SubCellInst_LFInst_4_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_4_LFInst_2_U10  ( .A1(
        \Red_SubCellInst_LFInst_4_LFInst_2_n19 ), .A2(
        \Red_SubCellInst_LFInst_4_LFInst_2_n18 ), .ZN(Red_MCOutput2[18]) );
  AND2_X1 \Red_SubCellInst_LFInst_4_LFInst_2_U9  ( .A1(
        \Red_SubCellInst_LFInst_4_LFInst_2_n17 ), .A2(PermutationOutput[16]), 
        .ZN(\Red_SubCellInst_LFInst_4_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_4_LFInst_2_U8  ( .A1(PermutationOutput[18]), 
        .A2(PermutationOutput[17]), .ZN(
        \Red_SubCellInst_LFInst_4_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_4_LFInst_2_U7  ( .A(
        \Red_SubCellInst_LFInst_4_LFInst_2_n16 ), .B(
        \Red_SubCellInst_LFInst_4_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst_LFInst_4_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_4_LFInst_2_U6  ( .A1(PermutationOutput[19]), 
        .A2(\Red_SubCellInst_LFInst_4_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst_LFInst_4_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst_LFInst_4_LFInst_2_U5  ( .A(PermutationOutput[17]), 
        .ZN(\Red_SubCellInst_LFInst_4_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_4_LFInst_2_U4  ( .A1(PermutationOutput[18]), 
        .A2(\Red_SubCellInst_LFInst_4_LFInst_2_n13 ), .ZN(
        \Red_SubCellInst_LFInst_4_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst_LFInst_4_LFInst_2_U3  ( .A(PermutationOutput[16]), 
        .ZN(\Red_SubCellInst_LFInst_4_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_4_LFInst_3_U6  ( .A(PermutationOutput[17]), 
        .B(\Red_SubCellInst_LFInst_4_LFInst_3_n8 ), .ZN(Red_MCOutput2[19]) );
  NOR2_X1 \Red_SubCellInst_LFInst_4_LFInst_3_U5  ( .A1(
        \Red_SubCellInst_LFInst_4_LFInst_3_n7 ), .A2(
        \Red_SubCellInst_LFInst_4_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst_LFInst_4_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_4_LFInst_3_U4  ( .A1(PermutationOutput[18]), 
        .A2(PermutationOutput[19]), .ZN(\Red_SubCellInst_LFInst_4_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst_LFInst_4_LFInst_3_U3  ( .A1(PermutationOutput[19]), 
        .A2(PermutationOutput[16]), .ZN(\Red_SubCellInst_LFInst_4_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_5_LFInst_0_U10  ( .A1(
        \Red_SubCellInst_LFInst_5_LFInst_0_n14 ), .A2(
        \Red_SubCellInst_LFInst_5_LFInst_0_n13 ), .ZN(Red_MCOutput2[20]) );
  NAND2_X1 \Red_SubCellInst_LFInst_5_LFInst_0_U9  ( .A1(PermutationOutput[20]), 
        .A2(\Red_SubCellInst_LFInst_5_LFInst_0_n12 ), .ZN(
        \Red_SubCellInst_LFInst_5_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_5_LFInst_0_U8  ( .A1(
        \Red_SubCellInst_LFInst_5_LFInst_0_n11 ), .A2(PermutationOutput[22]), 
        .ZN(\Red_SubCellInst_LFInst_5_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_5_LFInst_0_U7  ( .A(
        \Red_SubCellInst_LFInst_5_LFInst_0_n10 ), .B(
        \Red_SubCellInst_LFInst_5_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst_LFInst_5_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_5_LFInst_0_U6  ( .A1(PermutationOutput[23]), 
        .A2(\Red_SubCellInst_LFInst_5_LFInst_0_n11 ), .ZN(
        \Red_SubCellInst_LFInst_5_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst_LFInst_5_LFInst_0_U5  ( .A(PermutationOutput[21]), 
        .ZN(\Red_SubCellInst_LFInst_5_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_5_LFInst_0_U4  ( .A1(PermutationOutput[22]), 
        .A2(\Red_SubCellInst_LFInst_5_LFInst_0_n8 ), .ZN(
        \Red_SubCellInst_LFInst_5_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst_LFInst_5_LFInst_0_U3  ( .A(PermutationOutput[20]), 
        .ZN(\Red_SubCellInst_LFInst_5_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_5_LFInst_1_U8  ( .A1(
        \Red_SubCellInst_LFInst_5_LFInst_1_n15 ), .A2(
        \Red_SubCellInst_LFInst_5_LFInst_1_n14 ), .ZN(Red_MCOutput2[21]) );
  NAND2_X1 \Red_SubCellInst_LFInst_5_LFInst_1_U7  ( .A1(
        \Red_SubCellInst_LFInst_5_LFInst_1_n13 ), .A2(PermutationOutput[21]), 
        .ZN(\Red_SubCellInst_LFInst_5_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_5_LFInst_1_U6  ( .A1(
        \Red_SubCellInst_LFInst_5_LFInst_1_n12 ), .A2(PermutationOutput[20]), 
        .ZN(\Red_SubCellInst_LFInst_5_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_5_LFInst_1_U5  ( .A1(PermutationOutput[23]), 
        .A2(PermutationOutput[22]), .ZN(
        \Red_SubCellInst_LFInst_5_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst_LFInst_5_LFInst_1_U4  ( .A1(PermutationOutput[22]), 
        .A2(\Red_SubCellInst_LFInst_5_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst_LFInst_5_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_5_LFInst_1_U3  ( .A(PermutationOutput[20]), 
        .B(PermutationOutput[23]), .ZN(\Red_SubCellInst_LFInst_5_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_5_LFInst_2_U10  ( .A1(
        \Red_SubCellInst_LFInst_5_LFInst_2_n19 ), .A2(
        \Red_SubCellInst_LFInst_5_LFInst_2_n18 ), .ZN(Red_MCOutput2[22]) );
  AND2_X1 \Red_SubCellInst_LFInst_5_LFInst_2_U9  ( .A1(
        \Red_SubCellInst_LFInst_5_LFInst_2_n17 ), .A2(PermutationOutput[20]), 
        .ZN(\Red_SubCellInst_LFInst_5_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_5_LFInst_2_U8  ( .A1(PermutationOutput[22]), 
        .A2(PermutationOutput[21]), .ZN(
        \Red_SubCellInst_LFInst_5_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_5_LFInst_2_U7  ( .A(
        \Red_SubCellInst_LFInst_5_LFInst_2_n16 ), .B(
        \Red_SubCellInst_LFInst_5_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst_LFInst_5_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_5_LFInst_2_U6  ( .A1(PermutationOutput[23]), 
        .A2(\Red_SubCellInst_LFInst_5_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst_LFInst_5_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst_LFInst_5_LFInst_2_U5  ( .A(PermutationOutput[21]), 
        .ZN(\Red_SubCellInst_LFInst_5_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_5_LFInst_2_U4  ( .A1(PermutationOutput[22]), 
        .A2(\Red_SubCellInst_LFInst_5_LFInst_2_n13 ), .ZN(
        \Red_SubCellInst_LFInst_5_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst_LFInst_5_LFInst_2_U3  ( .A(PermutationOutput[20]), 
        .ZN(\Red_SubCellInst_LFInst_5_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_5_LFInst_3_U6  ( .A(PermutationOutput[21]), 
        .B(\Red_SubCellInst_LFInst_5_LFInst_3_n8 ), .ZN(Red_MCOutput2[23]) );
  NOR2_X1 \Red_SubCellInst_LFInst_5_LFInst_3_U5  ( .A1(
        \Red_SubCellInst_LFInst_5_LFInst_3_n7 ), .A2(
        \Red_SubCellInst_LFInst_5_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst_LFInst_5_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_5_LFInst_3_U4  ( .A1(PermutationOutput[22]), 
        .A2(PermutationOutput[23]), .ZN(\Red_SubCellInst_LFInst_5_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst_LFInst_5_LFInst_3_U3  ( .A1(PermutationOutput[23]), 
        .A2(PermutationOutput[20]), .ZN(\Red_SubCellInst_LFInst_5_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_6_LFInst_0_U10  ( .A1(
        \Red_SubCellInst_LFInst_6_LFInst_0_n14 ), .A2(
        \Red_SubCellInst_LFInst_6_LFInst_0_n13 ), .ZN(Red_MCOutput2[24]) );
  NAND2_X1 \Red_SubCellInst_LFInst_6_LFInst_0_U9  ( .A1(PermutationOutput[24]), 
        .A2(\Red_SubCellInst_LFInst_6_LFInst_0_n12 ), .ZN(
        \Red_SubCellInst_LFInst_6_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_6_LFInst_0_U8  ( .A1(
        \Red_SubCellInst_LFInst_6_LFInst_0_n11 ), .A2(PermutationOutput[26]), 
        .ZN(\Red_SubCellInst_LFInst_6_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_6_LFInst_0_U7  ( .A(
        \Red_SubCellInst_LFInst_6_LFInst_0_n10 ), .B(
        \Red_SubCellInst_LFInst_6_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst_LFInst_6_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_6_LFInst_0_U6  ( .A1(PermutationOutput[27]), 
        .A2(\Red_SubCellInst_LFInst_6_LFInst_0_n11 ), .ZN(
        \Red_SubCellInst_LFInst_6_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst_LFInst_6_LFInst_0_U5  ( .A(PermutationOutput[25]), 
        .ZN(\Red_SubCellInst_LFInst_6_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_6_LFInst_0_U4  ( .A1(PermutationOutput[26]), 
        .A2(\Red_SubCellInst_LFInst_6_LFInst_0_n8 ), .ZN(
        \Red_SubCellInst_LFInst_6_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst_LFInst_6_LFInst_0_U3  ( .A(PermutationOutput[24]), 
        .ZN(\Red_SubCellInst_LFInst_6_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_6_LFInst_1_U8  ( .A1(
        \Red_SubCellInst_LFInst_6_LFInst_1_n15 ), .A2(
        \Red_SubCellInst_LFInst_6_LFInst_1_n14 ), .ZN(Red_MCOutput2[25]) );
  NAND2_X1 \Red_SubCellInst_LFInst_6_LFInst_1_U7  ( .A1(
        \Red_SubCellInst_LFInst_6_LFInst_1_n13 ), .A2(PermutationOutput[25]), 
        .ZN(\Red_SubCellInst_LFInst_6_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_6_LFInst_1_U6  ( .A1(
        \Red_SubCellInst_LFInst_6_LFInst_1_n12 ), .A2(PermutationOutput[24]), 
        .ZN(\Red_SubCellInst_LFInst_6_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_6_LFInst_1_U5  ( .A1(PermutationOutput[27]), 
        .A2(PermutationOutput[26]), .ZN(
        \Red_SubCellInst_LFInst_6_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst_LFInst_6_LFInst_1_U4  ( .A1(PermutationOutput[26]), 
        .A2(\Red_SubCellInst_LFInst_6_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst_LFInst_6_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_6_LFInst_1_U3  ( .A(PermutationOutput[24]), 
        .B(PermutationOutput[27]), .ZN(\Red_SubCellInst_LFInst_6_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_6_LFInst_2_U10  ( .A1(
        \Red_SubCellInst_LFInst_6_LFInst_2_n19 ), .A2(
        \Red_SubCellInst_LFInst_6_LFInst_2_n18 ), .ZN(Red_MCOutput2[26]) );
  AND2_X1 \Red_SubCellInst_LFInst_6_LFInst_2_U9  ( .A1(
        \Red_SubCellInst_LFInst_6_LFInst_2_n17 ), .A2(PermutationOutput[24]), 
        .ZN(\Red_SubCellInst_LFInst_6_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_6_LFInst_2_U8  ( .A1(PermutationOutput[26]), 
        .A2(PermutationOutput[25]), .ZN(
        \Red_SubCellInst_LFInst_6_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_6_LFInst_2_U7  ( .A(
        \Red_SubCellInst_LFInst_6_LFInst_2_n16 ), .B(
        \Red_SubCellInst_LFInst_6_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst_LFInst_6_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_6_LFInst_2_U6  ( .A1(PermutationOutput[27]), 
        .A2(\Red_SubCellInst_LFInst_6_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst_LFInst_6_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst_LFInst_6_LFInst_2_U5  ( .A(PermutationOutput[25]), 
        .ZN(\Red_SubCellInst_LFInst_6_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_6_LFInst_2_U4  ( .A1(PermutationOutput[26]), 
        .A2(\Red_SubCellInst_LFInst_6_LFInst_2_n13 ), .ZN(
        \Red_SubCellInst_LFInst_6_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst_LFInst_6_LFInst_2_U3  ( .A(PermutationOutput[24]), 
        .ZN(\Red_SubCellInst_LFInst_6_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_6_LFInst_3_U6  ( .A(PermutationOutput[25]), 
        .B(\Red_SubCellInst_LFInst_6_LFInst_3_n8 ), .ZN(Red_MCOutput2[27]) );
  NOR2_X1 \Red_SubCellInst_LFInst_6_LFInst_3_U5  ( .A1(
        \Red_SubCellInst_LFInst_6_LFInst_3_n7 ), .A2(
        \Red_SubCellInst_LFInst_6_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst_LFInst_6_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_6_LFInst_3_U4  ( .A1(PermutationOutput[26]), 
        .A2(PermutationOutput[27]), .ZN(\Red_SubCellInst_LFInst_6_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst_LFInst_6_LFInst_3_U3  ( .A1(PermutationOutput[27]), 
        .A2(PermutationOutput[24]), .ZN(\Red_SubCellInst_LFInst_6_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_7_LFInst_0_U10  ( .A1(
        \Red_SubCellInst_LFInst_7_LFInst_0_n14 ), .A2(
        \Red_SubCellInst_LFInst_7_LFInst_0_n13 ), .ZN(Red_MCOutput2[28]) );
  NAND2_X1 \Red_SubCellInst_LFInst_7_LFInst_0_U9  ( .A1(PermutationOutput[28]), 
        .A2(\Red_SubCellInst_LFInst_7_LFInst_0_n12 ), .ZN(
        \Red_SubCellInst_LFInst_7_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_7_LFInst_0_U8  ( .A1(
        \Red_SubCellInst_LFInst_7_LFInst_0_n11 ), .A2(PermutationOutput[30]), 
        .ZN(\Red_SubCellInst_LFInst_7_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_7_LFInst_0_U7  ( .A(
        \Red_SubCellInst_LFInst_7_LFInst_0_n10 ), .B(
        \Red_SubCellInst_LFInst_7_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst_LFInst_7_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_7_LFInst_0_U6  ( .A1(PermutationOutput[31]), 
        .A2(\Red_SubCellInst_LFInst_7_LFInst_0_n11 ), .ZN(
        \Red_SubCellInst_LFInst_7_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst_LFInst_7_LFInst_0_U5  ( .A(PermutationOutput[29]), 
        .ZN(\Red_SubCellInst_LFInst_7_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_7_LFInst_0_U4  ( .A1(PermutationOutput[30]), 
        .A2(\Red_SubCellInst_LFInst_7_LFInst_0_n8 ), .ZN(
        \Red_SubCellInst_LFInst_7_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst_LFInst_7_LFInst_0_U3  ( .A(PermutationOutput[28]), 
        .ZN(\Red_SubCellInst_LFInst_7_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_7_LFInst_1_U8  ( .A1(
        \Red_SubCellInst_LFInst_7_LFInst_1_n15 ), .A2(
        \Red_SubCellInst_LFInst_7_LFInst_1_n14 ), .ZN(Red_MCOutput2[29]) );
  NAND2_X1 \Red_SubCellInst_LFInst_7_LFInst_1_U7  ( .A1(
        \Red_SubCellInst_LFInst_7_LFInst_1_n13 ), .A2(PermutationOutput[29]), 
        .ZN(\Red_SubCellInst_LFInst_7_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_7_LFInst_1_U6  ( .A1(
        \Red_SubCellInst_LFInst_7_LFInst_1_n12 ), .A2(PermutationOutput[28]), 
        .ZN(\Red_SubCellInst_LFInst_7_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_7_LFInst_1_U5  ( .A1(PermutationOutput[31]), 
        .A2(PermutationOutput[30]), .ZN(
        \Red_SubCellInst_LFInst_7_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst_LFInst_7_LFInst_1_U4  ( .A1(PermutationOutput[30]), 
        .A2(\Red_SubCellInst_LFInst_7_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst_LFInst_7_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_7_LFInst_1_U3  ( .A(PermutationOutput[28]), 
        .B(PermutationOutput[31]), .ZN(\Red_SubCellInst_LFInst_7_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_7_LFInst_2_U10  ( .A1(
        \Red_SubCellInst_LFInst_7_LFInst_2_n19 ), .A2(
        \Red_SubCellInst_LFInst_7_LFInst_2_n18 ), .ZN(Red_MCOutput2[30]) );
  AND2_X1 \Red_SubCellInst_LFInst_7_LFInst_2_U9  ( .A1(
        \Red_SubCellInst_LFInst_7_LFInst_2_n17 ), .A2(PermutationOutput[28]), 
        .ZN(\Red_SubCellInst_LFInst_7_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_7_LFInst_2_U8  ( .A1(PermutationOutput[30]), 
        .A2(PermutationOutput[29]), .ZN(
        \Red_SubCellInst_LFInst_7_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_7_LFInst_2_U7  ( .A(
        \Red_SubCellInst_LFInst_7_LFInst_2_n16 ), .B(
        \Red_SubCellInst_LFInst_7_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst_LFInst_7_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_7_LFInst_2_U6  ( .A1(PermutationOutput[31]), 
        .A2(\Red_SubCellInst_LFInst_7_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst_LFInst_7_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst_LFInst_7_LFInst_2_U5  ( .A(PermutationOutput[29]), 
        .ZN(\Red_SubCellInst_LFInst_7_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_7_LFInst_2_U4  ( .A1(PermutationOutput[30]), 
        .A2(\Red_SubCellInst_LFInst_7_LFInst_2_n13 ), .ZN(
        \Red_SubCellInst_LFInst_7_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst_LFInst_7_LFInst_2_U3  ( .A(PermutationOutput[28]), 
        .ZN(\Red_SubCellInst_LFInst_7_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_7_LFInst_3_U6  ( .A(PermutationOutput[29]), 
        .B(\Red_SubCellInst_LFInst_7_LFInst_3_n8 ), .ZN(Red_MCOutput2[31]) );
  NOR2_X1 \Red_SubCellInst_LFInst_7_LFInst_3_U5  ( .A1(
        \Red_SubCellInst_LFInst_7_LFInst_3_n7 ), .A2(
        \Red_SubCellInst_LFInst_7_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst_LFInst_7_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_7_LFInst_3_U4  ( .A1(PermutationOutput[30]), 
        .A2(PermutationOutput[31]), .ZN(\Red_SubCellInst_LFInst_7_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst_LFInst_7_LFInst_3_U3  ( .A1(PermutationOutput[31]), 
        .A2(PermutationOutput[28]), .ZN(\Red_SubCellInst_LFInst_7_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_8_LFInst_0_U10  ( .A1(
        \Red_SubCellInst_LFInst_8_LFInst_0_n14 ), .A2(
        \Red_SubCellInst_LFInst_8_LFInst_0_n13 ), .ZN(Red_Feedback[32]) );
  NAND2_X1 \Red_SubCellInst_LFInst_8_LFInst_0_U9  ( .A1(PermutationOutput[32]), 
        .A2(\Red_SubCellInst_LFInst_8_LFInst_0_n12 ), .ZN(
        \Red_SubCellInst_LFInst_8_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_8_LFInst_0_U8  ( .A1(
        \Red_SubCellInst_LFInst_8_LFInst_0_n11 ), .A2(PermutationOutput[34]), 
        .ZN(\Red_SubCellInst_LFInst_8_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_8_LFInst_0_U7  ( .A(
        \Red_SubCellInst_LFInst_8_LFInst_0_n10 ), .B(
        \Red_SubCellInst_LFInst_8_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst_LFInst_8_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_8_LFInst_0_U6  ( .A1(PermutationOutput[35]), 
        .A2(\Red_SubCellInst_LFInst_8_LFInst_0_n11 ), .ZN(
        \Red_SubCellInst_LFInst_8_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst_LFInst_8_LFInst_0_U5  ( .A(PermutationOutput[33]), 
        .ZN(\Red_SubCellInst_LFInst_8_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_8_LFInst_0_U4  ( .A1(PermutationOutput[34]), 
        .A2(\Red_SubCellInst_LFInst_8_LFInst_0_n8 ), .ZN(
        \Red_SubCellInst_LFInst_8_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst_LFInst_8_LFInst_0_U3  ( .A(PermutationOutput[32]), 
        .ZN(\Red_SubCellInst_LFInst_8_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_8_LFInst_1_U8  ( .A1(
        \Red_SubCellInst_LFInst_8_LFInst_1_n15 ), .A2(
        \Red_SubCellInst_LFInst_8_LFInst_1_n14 ), .ZN(Red_Feedback[33]) );
  NAND2_X1 \Red_SubCellInst_LFInst_8_LFInst_1_U7  ( .A1(
        \Red_SubCellInst_LFInst_8_LFInst_1_n13 ), .A2(PermutationOutput[33]), 
        .ZN(\Red_SubCellInst_LFInst_8_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_8_LFInst_1_U6  ( .A1(
        \Red_SubCellInst_LFInst_8_LFInst_1_n12 ), .A2(PermutationOutput[32]), 
        .ZN(\Red_SubCellInst_LFInst_8_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_8_LFInst_1_U5  ( .A1(PermutationOutput[35]), 
        .A2(PermutationOutput[34]), .ZN(
        \Red_SubCellInst_LFInst_8_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst_LFInst_8_LFInst_1_U4  ( .A1(PermutationOutput[34]), 
        .A2(\Red_SubCellInst_LFInst_8_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst_LFInst_8_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_8_LFInst_1_U3  ( .A(PermutationOutput[32]), 
        .B(PermutationOutput[35]), .ZN(\Red_SubCellInst_LFInst_8_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_8_LFInst_2_U10  ( .A1(
        \Red_SubCellInst_LFInst_8_LFInst_2_n19 ), .A2(
        \Red_SubCellInst_LFInst_8_LFInst_2_n18 ), .ZN(Red_Feedback[34]) );
  AND2_X1 \Red_SubCellInst_LFInst_8_LFInst_2_U9  ( .A1(
        \Red_SubCellInst_LFInst_8_LFInst_2_n17 ), .A2(PermutationOutput[32]), 
        .ZN(\Red_SubCellInst_LFInst_8_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_8_LFInst_2_U8  ( .A1(PermutationOutput[34]), 
        .A2(PermutationOutput[33]), .ZN(
        \Red_SubCellInst_LFInst_8_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_8_LFInst_2_U7  ( .A(
        \Red_SubCellInst_LFInst_8_LFInst_2_n16 ), .B(
        \Red_SubCellInst_LFInst_8_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst_LFInst_8_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_8_LFInst_2_U6  ( .A1(PermutationOutput[35]), 
        .A2(\Red_SubCellInst_LFInst_8_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst_LFInst_8_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst_LFInst_8_LFInst_2_U5  ( .A(PermutationOutput[33]), 
        .ZN(\Red_SubCellInst_LFInst_8_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_8_LFInst_2_U4  ( .A1(PermutationOutput[34]), 
        .A2(\Red_SubCellInst_LFInst_8_LFInst_2_n13 ), .ZN(
        \Red_SubCellInst_LFInst_8_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst_LFInst_8_LFInst_2_U3  ( .A(PermutationOutput[32]), 
        .ZN(\Red_SubCellInst_LFInst_8_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_8_LFInst_3_U6  ( .A(PermutationOutput[33]), 
        .B(\Red_SubCellInst_LFInst_8_LFInst_3_n8 ), .ZN(Red_Feedback[35]) );
  NOR2_X1 \Red_SubCellInst_LFInst_8_LFInst_3_U5  ( .A1(
        \Red_SubCellInst_LFInst_8_LFInst_3_n7 ), .A2(
        \Red_SubCellInst_LFInst_8_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst_LFInst_8_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_8_LFInst_3_U4  ( .A1(PermutationOutput[34]), 
        .A2(PermutationOutput[35]), .ZN(\Red_SubCellInst_LFInst_8_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst_LFInst_8_LFInst_3_U3  ( .A1(PermutationOutput[35]), 
        .A2(PermutationOutput[32]), .ZN(\Red_SubCellInst_LFInst_8_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_9_LFInst_0_U10  ( .A1(
        \Red_SubCellInst_LFInst_9_LFInst_0_n14 ), .A2(
        \Red_SubCellInst_LFInst_9_LFInst_0_n13 ), .ZN(Red_Feedback[36]) );
  NAND2_X1 \Red_SubCellInst_LFInst_9_LFInst_0_U9  ( .A1(PermutationOutput[36]), 
        .A2(\Red_SubCellInst_LFInst_9_LFInst_0_n12 ), .ZN(
        \Red_SubCellInst_LFInst_9_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_9_LFInst_0_U8  ( .A1(
        \Red_SubCellInst_LFInst_9_LFInst_0_n11 ), .A2(PermutationOutput[38]), 
        .ZN(\Red_SubCellInst_LFInst_9_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_9_LFInst_0_U7  ( .A(
        \Red_SubCellInst_LFInst_9_LFInst_0_n10 ), .B(
        \Red_SubCellInst_LFInst_9_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst_LFInst_9_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_9_LFInst_0_U6  ( .A1(PermutationOutput[39]), 
        .A2(\Red_SubCellInst_LFInst_9_LFInst_0_n11 ), .ZN(
        \Red_SubCellInst_LFInst_9_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst_LFInst_9_LFInst_0_U5  ( .A(PermutationOutput[37]), 
        .ZN(\Red_SubCellInst_LFInst_9_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_9_LFInst_0_U4  ( .A1(PermutationOutput[38]), 
        .A2(\Red_SubCellInst_LFInst_9_LFInst_0_n8 ), .ZN(
        \Red_SubCellInst_LFInst_9_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst_LFInst_9_LFInst_0_U3  ( .A(PermutationOutput[36]), 
        .ZN(\Red_SubCellInst_LFInst_9_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_9_LFInst_1_U8  ( .A1(
        \Red_SubCellInst_LFInst_9_LFInst_1_n15 ), .A2(
        \Red_SubCellInst_LFInst_9_LFInst_1_n14 ), .ZN(Red_Feedback[37]) );
  NAND2_X1 \Red_SubCellInst_LFInst_9_LFInst_1_U7  ( .A1(
        \Red_SubCellInst_LFInst_9_LFInst_1_n13 ), .A2(PermutationOutput[37]), 
        .ZN(\Red_SubCellInst_LFInst_9_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_9_LFInst_1_U6  ( .A1(
        \Red_SubCellInst_LFInst_9_LFInst_1_n12 ), .A2(PermutationOutput[36]), 
        .ZN(\Red_SubCellInst_LFInst_9_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_9_LFInst_1_U5  ( .A1(PermutationOutput[39]), 
        .A2(PermutationOutput[38]), .ZN(
        \Red_SubCellInst_LFInst_9_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst_LFInst_9_LFInst_1_U4  ( .A1(PermutationOutput[38]), 
        .A2(\Red_SubCellInst_LFInst_9_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst_LFInst_9_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_9_LFInst_1_U3  ( .A(PermutationOutput[36]), 
        .B(PermutationOutput[39]), .ZN(\Red_SubCellInst_LFInst_9_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_9_LFInst_2_U10  ( .A1(
        \Red_SubCellInst_LFInst_9_LFInst_2_n19 ), .A2(
        \Red_SubCellInst_LFInst_9_LFInst_2_n18 ), .ZN(Red_Feedback[38]) );
  AND2_X1 \Red_SubCellInst_LFInst_9_LFInst_2_U9  ( .A1(
        \Red_SubCellInst_LFInst_9_LFInst_2_n17 ), .A2(PermutationOutput[36]), 
        .ZN(\Red_SubCellInst_LFInst_9_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_9_LFInst_2_U8  ( .A1(PermutationOutput[38]), 
        .A2(PermutationOutput[37]), .ZN(
        \Red_SubCellInst_LFInst_9_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_9_LFInst_2_U7  ( .A(
        \Red_SubCellInst_LFInst_9_LFInst_2_n16 ), .B(
        \Red_SubCellInst_LFInst_9_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst_LFInst_9_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_9_LFInst_2_U6  ( .A1(PermutationOutput[39]), 
        .A2(\Red_SubCellInst_LFInst_9_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst_LFInst_9_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst_LFInst_9_LFInst_2_U5  ( .A(PermutationOutput[37]), 
        .ZN(\Red_SubCellInst_LFInst_9_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_9_LFInst_2_U4  ( .A1(PermutationOutput[38]), 
        .A2(\Red_SubCellInst_LFInst_9_LFInst_2_n13 ), .ZN(
        \Red_SubCellInst_LFInst_9_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst_LFInst_9_LFInst_2_U3  ( .A(PermutationOutput[36]), 
        .ZN(\Red_SubCellInst_LFInst_9_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_9_LFInst_3_U6  ( .A(PermutationOutput[37]), 
        .B(\Red_SubCellInst_LFInst_9_LFInst_3_n8 ), .ZN(Red_Feedback[39]) );
  NOR2_X1 \Red_SubCellInst_LFInst_9_LFInst_3_U5  ( .A1(
        \Red_SubCellInst_LFInst_9_LFInst_3_n7 ), .A2(
        \Red_SubCellInst_LFInst_9_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst_LFInst_9_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_9_LFInst_3_U4  ( .A1(PermutationOutput[38]), 
        .A2(PermutationOutput[39]), .ZN(\Red_SubCellInst_LFInst_9_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst_LFInst_9_LFInst_3_U3  ( .A1(PermutationOutput[39]), 
        .A2(PermutationOutput[36]), .ZN(\Red_SubCellInst_LFInst_9_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_10_LFInst_0_U10  ( .A1(
        \Red_SubCellInst_LFInst_10_LFInst_0_n14 ), .A2(
        \Red_SubCellInst_LFInst_10_LFInst_0_n13 ), .ZN(Red_Feedback[40]) );
  NAND2_X1 \Red_SubCellInst_LFInst_10_LFInst_0_U9  ( .A1(PermutationOutput[40]), .A2(\Red_SubCellInst_LFInst_10_LFInst_0_n12 ), .ZN(
        \Red_SubCellInst_LFInst_10_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_10_LFInst_0_U8  ( .A1(
        \Red_SubCellInst_LFInst_10_LFInst_0_n11 ), .A2(PermutationOutput[42]), 
        .ZN(\Red_SubCellInst_LFInst_10_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_10_LFInst_0_U7  ( .A(
        \Red_SubCellInst_LFInst_10_LFInst_0_n10 ), .B(
        \Red_SubCellInst_LFInst_10_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst_LFInst_10_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_10_LFInst_0_U6  ( .A1(PermutationOutput[43]), .A2(\Red_SubCellInst_LFInst_10_LFInst_0_n11 ), .ZN(
        \Red_SubCellInst_LFInst_10_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst_LFInst_10_LFInst_0_U5  ( .A(PermutationOutput[41]), 
        .ZN(\Red_SubCellInst_LFInst_10_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_10_LFInst_0_U4  ( .A1(PermutationOutput[42]), .A2(\Red_SubCellInst_LFInst_10_LFInst_0_n8 ), .ZN(
        \Red_SubCellInst_LFInst_10_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst_LFInst_10_LFInst_0_U3  ( .A(PermutationOutput[40]), 
        .ZN(\Red_SubCellInst_LFInst_10_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_10_LFInst_1_U8  ( .A1(
        \Red_SubCellInst_LFInst_10_LFInst_1_n15 ), .A2(
        \Red_SubCellInst_LFInst_10_LFInst_1_n14 ), .ZN(Red_Feedback[41]) );
  NAND2_X1 \Red_SubCellInst_LFInst_10_LFInst_1_U7  ( .A1(
        \Red_SubCellInst_LFInst_10_LFInst_1_n13 ), .A2(PermutationOutput[41]), 
        .ZN(\Red_SubCellInst_LFInst_10_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_10_LFInst_1_U6  ( .A1(
        \Red_SubCellInst_LFInst_10_LFInst_1_n12 ), .A2(PermutationOutput[40]), 
        .ZN(\Red_SubCellInst_LFInst_10_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_10_LFInst_1_U5  ( .A1(PermutationOutput[43]), .A2(PermutationOutput[42]), .ZN(\Red_SubCellInst_LFInst_10_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst_LFInst_10_LFInst_1_U4  ( .A1(PermutationOutput[42]), 
        .A2(\Red_SubCellInst_LFInst_10_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst_LFInst_10_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_10_LFInst_1_U3  ( .A(PermutationOutput[40]), 
        .B(PermutationOutput[43]), .ZN(
        \Red_SubCellInst_LFInst_10_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_10_LFInst_2_U10  ( .A1(
        \Red_SubCellInst_LFInst_10_LFInst_2_n19 ), .A2(
        \Red_SubCellInst_LFInst_10_LFInst_2_n18 ), .ZN(Red_Feedback[42]) );
  AND2_X1 \Red_SubCellInst_LFInst_10_LFInst_2_U9  ( .A1(
        \Red_SubCellInst_LFInst_10_LFInst_2_n17 ), .A2(PermutationOutput[40]), 
        .ZN(\Red_SubCellInst_LFInst_10_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_10_LFInst_2_U8  ( .A1(PermutationOutput[42]), 
        .A2(PermutationOutput[41]), .ZN(
        \Red_SubCellInst_LFInst_10_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_10_LFInst_2_U7  ( .A(
        \Red_SubCellInst_LFInst_10_LFInst_2_n16 ), .B(
        \Red_SubCellInst_LFInst_10_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst_LFInst_10_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_10_LFInst_2_U6  ( .A1(PermutationOutput[43]), 
        .A2(\Red_SubCellInst_LFInst_10_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst_LFInst_10_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst_LFInst_10_LFInst_2_U5  ( .A(PermutationOutput[41]), 
        .ZN(\Red_SubCellInst_LFInst_10_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_10_LFInst_2_U4  ( .A1(PermutationOutput[42]), .A2(\Red_SubCellInst_LFInst_10_LFInst_2_n13 ), .ZN(
        \Red_SubCellInst_LFInst_10_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst_LFInst_10_LFInst_2_U3  ( .A(PermutationOutput[40]), 
        .ZN(\Red_SubCellInst_LFInst_10_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_10_LFInst_3_U6  ( .A(PermutationOutput[41]), 
        .B(\Red_SubCellInst_LFInst_10_LFInst_3_n8 ), .ZN(Red_Feedback[43]) );
  NOR2_X1 \Red_SubCellInst_LFInst_10_LFInst_3_U5  ( .A1(
        \Red_SubCellInst_LFInst_10_LFInst_3_n7 ), .A2(
        \Red_SubCellInst_LFInst_10_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst_LFInst_10_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_10_LFInst_3_U4  ( .A1(PermutationOutput[42]), 
        .A2(PermutationOutput[43]), .ZN(
        \Red_SubCellInst_LFInst_10_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst_LFInst_10_LFInst_3_U3  ( .A1(PermutationOutput[43]), 
        .A2(PermutationOutput[40]), .ZN(
        \Red_SubCellInst_LFInst_10_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_11_LFInst_0_U10  ( .A1(
        \Red_SubCellInst_LFInst_11_LFInst_0_n14 ), .A2(
        \Red_SubCellInst_LFInst_11_LFInst_0_n13 ), .ZN(Red_Feedback[44]) );
  NAND2_X1 \Red_SubCellInst_LFInst_11_LFInst_0_U9  ( .A1(PermutationOutput[44]), .A2(\Red_SubCellInst_LFInst_11_LFInst_0_n12 ), .ZN(
        \Red_SubCellInst_LFInst_11_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_11_LFInst_0_U8  ( .A1(
        \Red_SubCellInst_LFInst_11_LFInst_0_n11 ), .A2(PermutationOutput[46]), 
        .ZN(\Red_SubCellInst_LFInst_11_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_11_LFInst_0_U7  ( .A(
        \Red_SubCellInst_LFInst_11_LFInst_0_n10 ), .B(
        \Red_SubCellInst_LFInst_11_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst_LFInst_11_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_11_LFInst_0_U6  ( .A1(PermutationOutput[47]), .A2(\Red_SubCellInst_LFInst_11_LFInst_0_n11 ), .ZN(
        \Red_SubCellInst_LFInst_11_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst_LFInst_11_LFInst_0_U5  ( .A(PermutationOutput[45]), 
        .ZN(\Red_SubCellInst_LFInst_11_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_11_LFInst_0_U4  ( .A1(PermutationOutput[46]), .A2(\Red_SubCellInst_LFInst_11_LFInst_0_n8 ), .ZN(
        \Red_SubCellInst_LFInst_11_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst_LFInst_11_LFInst_0_U3  ( .A(PermutationOutput[44]), 
        .ZN(\Red_SubCellInst_LFInst_11_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_11_LFInst_1_U8  ( .A1(
        \Red_SubCellInst_LFInst_11_LFInst_1_n15 ), .A2(
        \Red_SubCellInst_LFInst_11_LFInst_1_n14 ), .ZN(Red_Feedback[45]) );
  NAND2_X1 \Red_SubCellInst_LFInst_11_LFInst_1_U7  ( .A1(
        \Red_SubCellInst_LFInst_11_LFInst_1_n13 ), .A2(PermutationOutput[45]), 
        .ZN(\Red_SubCellInst_LFInst_11_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_11_LFInst_1_U6  ( .A1(
        \Red_SubCellInst_LFInst_11_LFInst_1_n12 ), .A2(PermutationOutput[44]), 
        .ZN(\Red_SubCellInst_LFInst_11_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_11_LFInst_1_U5  ( .A1(PermutationOutput[47]), .A2(PermutationOutput[46]), .ZN(\Red_SubCellInst_LFInst_11_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst_LFInst_11_LFInst_1_U4  ( .A1(PermutationOutput[46]), 
        .A2(\Red_SubCellInst_LFInst_11_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst_LFInst_11_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_11_LFInst_1_U3  ( .A(PermutationOutput[44]), 
        .B(PermutationOutput[47]), .ZN(
        \Red_SubCellInst_LFInst_11_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_11_LFInst_2_U10  ( .A1(
        \Red_SubCellInst_LFInst_11_LFInst_2_n19 ), .A2(
        \Red_SubCellInst_LFInst_11_LFInst_2_n18 ), .ZN(Red_Feedback[46]) );
  AND2_X1 \Red_SubCellInst_LFInst_11_LFInst_2_U9  ( .A1(
        \Red_SubCellInst_LFInst_11_LFInst_2_n17 ), .A2(PermutationOutput[44]), 
        .ZN(\Red_SubCellInst_LFInst_11_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_11_LFInst_2_U8  ( .A1(PermutationOutput[46]), 
        .A2(PermutationOutput[45]), .ZN(
        \Red_SubCellInst_LFInst_11_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_11_LFInst_2_U7  ( .A(
        \Red_SubCellInst_LFInst_11_LFInst_2_n16 ), .B(
        \Red_SubCellInst_LFInst_11_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst_LFInst_11_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_11_LFInst_2_U6  ( .A1(PermutationOutput[47]), 
        .A2(\Red_SubCellInst_LFInst_11_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst_LFInst_11_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst_LFInst_11_LFInst_2_U5  ( .A(PermutationOutput[45]), 
        .ZN(\Red_SubCellInst_LFInst_11_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_11_LFInst_2_U4  ( .A1(PermutationOutput[46]), .A2(\Red_SubCellInst_LFInst_11_LFInst_2_n13 ), .ZN(
        \Red_SubCellInst_LFInst_11_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst_LFInst_11_LFInst_2_U3  ( .A(PermutationOutput[44]), 
        .ZN(\Red_SubCellInst_LFInst_11_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_11_LFInst_3_U6  ( .A(PermutationOutput[45]), 
        .B(\Red_SubCellInst_LFInst_11_LFInst_3_n8 ), .ZN(Red_Feedback[47]) );
  NOR2_X1 \Red_SubCellInst_LFInst_11_LFInst_3_U5  ( .A1(
        \Red_SubCellInst_LFInst_11_LFInst_3_n7 ), .A2(
        \Red_SubCellInst_LFInst_11_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst_LFInst_11_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_11_LFInst_3_U4  ( .A1(PermutationOutput[46]), 
        .A2(PermutationOutput[47]), .ZN(
        \Red_SubCellInst_LFInst_11_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst_LFInst_11_LFInst_3_U3  ( .A1(PermutationOutput[47]), 
        .A2(PermutationOutput[44]), .ZN(
        \Red_SubCellInst_LFInst_11_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_12_LFInst_0_U10  ( .A1(
        \Red_SubCellInst_LFInst_12_LFInst_0_n14 ), .A2(
        \Red_SubCellInst_LFInst_12_LFInst_0_n13 ), .ZN(Red_Feedback[48]) );
  NAND2_X1 \Red_SubCellInst_LFInst_12_LFInst_0_U9  ( .A1(PermutationOutput[48]), .A2(\Red_SubCellInst_LFInst_12_LFInst_0_n12 ), .ZN(
        \Red_SubCellInst_LFInst_12_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_12_LFInst_0_U8  ( .A1(
        \Red_SubCellInst_LFInst_12_LFInst_0_n11 ), .A2(PermutationOutput[50]), 
        .ZN(\Red_SubCellInst_LFInst_12_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_12_LFInst_0_U7  ( .A(
        \Red_SubCellInst_LFInst_12_LFInst_0_n10 ), .B(
        \Red_SubCellInst_LFInst_12_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst_LFInst_12_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_12_LFInst_0_U6  ( .A1(PermutationOutput[51]), .A2(\Red_SubCellInst_LFInst_12_LFInst_0_n11 ), .ZN(
        \Red_SubCellInst_LFInst_12_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst_LFInst_12_LFInst_0_U5  ( .A(PermutationOutput[49]), 
        .ZN(\Red_SubCellInst_LFInst_12_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_12_LFInst_0_U4  ( .A1(PermutationOutput[50]), .A2(\Red_SubCellInst_LFInst_12_LFInst_0_n8 ), .ZN(
        \Red_SubCellInst_LFInst_12_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst_LFInst_12_LFInst_0_U3  ( .A(PermutationOutput[48]), 
        .ZN(\Red_SubCellInst_LFInst_12_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_12_LFInst_1_U8  ( .A1(
        \Red_SubCellInst_LFInst_12_LFInst_1_n15 ), .A2(
        \Red_SubCellInst_LFInst_12_LFInst_1_n14 ), .ZN(Red_Feedback[49]) );
  NAND2_X1 \Red_SubCellInst_LFInst_12_LFInst_1_U7  ( .A1(
        \Red_SubCellInst_LFInst_12_LFInst_1_n13 ), .A2(PermutationOutput[49]), 
        .ZN(\Red_SubCellInst_LFInst_12_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_12_LFInst_1_U6  ( .A1(
        \Red_SubCellInst_LFInst_12_LFInst_1_n12 ), .A2(PermutationOutput[48]), 
        .ZN(\Red_SubCellInst_LFInst_12_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_12_LFInst_1_U5  ( .A1(PermutationOutput[51]), .A2(PermutationOutput[50]), .ZN(\Red_SubCellInst_LFInst_12_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst_LFInst_12_LFInst_1_U4  ( .A1(PermutationOutput[50]), 
        .A2(\Red_SubCellInst_LFInst_12_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst_LFInst_12_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_12_LFInst_1_U3  ( .A(PermutationOutput[48]), 
        .B(PermutationOutput[51]), .ZN(
        \Red_SubCellInst_LFInst_12_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_12_LFInst_2_U10  ( .A1(
        \Red_SubCellInst_LFInst_12_LFInst_2_n19 ), .A2(
        \Red_SubCellInst_LFInst_12_LFInst_2_n18 ), .ZN(Red_Feedback[50]) );
  AND2_X1 \Red_SubCellInst_LFInst_12_LFInst_2_U9  ( .A1(
        \Red_SubCellInst_LFInst_12_LFInst_2_n17 ), .A2(PermutationOutput[48]), 
        .ZN(\Red_SubCellInst_LFInst_12_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_12_LFInst_2_U8  ( .A1(PermutationOutput[50]), 
        .A2(PermutationOutput[49]), .ZN(
        \Red_SubCellInst_LFInst_12_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_12_LFInst_2_U7  ( .A(
        \Red_SubCellInst_LFInst_12_LFInst_2_n16 ), .B(
        \Red_SubCellInst_LFInst_12_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst_LFInst_12_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_12_LFInst_2_U6  ( .A1(PermutationOutput[51]), 
        .A2(\Red_SubCellInst_LFInst_12_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst_LFInst_12_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst_LFInst_12_LFInst_2_U5  ( .A(PermutationOutput[49]), 
        .ZN(\Red_SubCellInst_LFInst_12_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_12_LFInst_2_U4  ( .A1(PermutationOutput[50]), .A2(\Red_SubCellInst_LFInst_12_LFInst_2_n13 ), .ZN(
        \Red_SubCellInst_LFInst_12_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst_LFInst_12_LFInst_2_U3  ( .A(PermutationOutput[48]), 
        .ZN(\Red_SubCellInst_LFInst_12_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_12_LFInst_3_U6  ( .A(PermutationOutput[49]), 
        .B(\Red_SubCellInst_LFInst_12_LFInst_3_n8 ), .ZN(Red_Feedback[51]) );
  NOR2_X1 \Red_SubCellInst_LFInst_12_LFInst_3_U5  ( .A1(
        \Red_SubCellInst_LFInst_12_LFInst_3_n7 ), .A2(
        \Red_SubCellInst_LFInst_12_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst_LFInst_12_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_12_LFInst_3_U4  ( .A1(PermutationOutput[50]), 
        .A2(PermutationOutput[51]), .ZN(
        \Red_SubCellInst_LFInst_12_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst_LFInst_12_LFInst_3_U3  ( .A1(PermutationOutput[51]), 
        .A2(PermutationOutput[48]), .ZN(
        \Red_SubCellInst_LFInst_12_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_13_LFInst_0_U10  ( .A1(
        \Red_SubCellInst_LFInst_13_LFInst_0_n14 ), .A2(
        \Red_SubCellInst_LFInst_13_LFInst_0_n13 ), .ZN(Red_Feedback[52]) );
  NAND2_X1 \Red_SubCellInst_LFInst_13_LFInst_0_U9  ( .A1(PermutationOutput[52]), .A2(\Red_SubCellInst_LFInst_13_LFInst_0_n12 ), .ZN(
        \Red_SubCellInst_LFInst_13_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_13_LFInst_0_U8  ( .A1(
        \Red_SubCellInst_LFInst_13_LFInst_0_n11 ), .A2(PermutationOutput[54]), 
        .ZN(\Red_SubCellInst_LFInst_13_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_13_LFInst_0_U7  ( .A(
        \Red_SubCellInst_LFInst_13_LFInst_0_n10 ), .B(
        \Red_SubCellInst_LFInst_13_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst_LFInst_13_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_13_LFInst_0_U6  ( .A1(PermutationOutput[55]), .A2(\Red_SubCellInst_LFInst_13_LFInst_0_n11 ), .ZN(
        \Red_SubCellInst_LFInst_13_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst_LFInst_13_LFInst_0_U5  ( .A(PermutationOutput[53]), 
        .ZN(\Red_SubCellInst_LFInst_13_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_13_LFInst_0_U4  ( .A1(PermutationOutput[54]), .A2(\Red_SubCellInst_LFInst_13_LFInst_0_n8 ), .ZN(
        \Red_SubCellInst_LFInst_13_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst_LFInst_13_LFInst_0_U3  ( .A(PermutationOutput[52]), 
        .ZN(\Red_SubCellInst_LFInst_13_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_13_LFInst_1_U8  ( .A1(
        \Red_SubCellInst_LFInst_13_LFInst_1_n15 ), .A2(
        \Red_SubCellInst_LFInst_13_LFInst_1_n14 ), .ZN(Red_Feedback[53]) );
  NAND2_X1 \Red_SubCellInst_LFInst_13_LFInst_1_U7  ( .A1(
        \Red_SubCellInst_LFInst_13_LFInst_1_n13 ), .A2(PermutationOutput[53]), 
        .ZN(\Red_SubCellInst_LFInst_13_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_13_LFInst_1_U6  ( .A1(
        \Red_SubCellInst_LFInst_13_LFInst_1_n12 ), .A2(PermutationOutput[52]), 
        .ZN(\Red_SubCellInst_LFInst_13_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_13_LFInst_1_U5  ( .A1(PermutationOutput[55]), .A2(PermutationOutput[54]), .ZN(\Red_SubCellInst_LFInst_13_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst_LFInst_13_LFInst_1_U4  ( .A1(PermutationOutput[54]), 
        .A2(\Red_SubCellInst_LFInst_13_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst_LFInst_13_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_13_LFInst_1_U3  ( .A(PermutationOutput[52]), 
        .B(PermutationOutput[55]), .ZN(
        \Red_SubCellInst_LFInst_13_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_13_LFInst_2_U10  ( .A1(
        \Red_SubCellInst_LFInst_13_LFInst_2_n19 ), .A2(
        \Red_SubCellInst_LFInst_13_LFInst_2_n18 ), .ZN(Red_Feedback[54]) );
  AND2_X1 \Red_SubCellInst_LFInst_13_LFInst_2_U9  ( .A1(
        \Red_SubCellInst_LFInst_13_LFInst_2_n17 ), .A2(PermutationOutput[52]), 
        .ZN(\Red_SubCellInst_LFInst_13_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_13_LFInst_2_U8  ( .A1(PermutationOutput[54]), 
        .A2(PermutationOutput[53]), .ZN(
        \Red_SubCellInst_LFInst_13_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_13_LFInst_2_U7  ( .A(
        \Red_SubCellInst_LFInst_13_LFInst_2_n16 ), .B(
        \Red_SubCellInst_LFInst_13_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst_LFInst_13_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_13_LFInst_2_U6  ( .A1(PermutationOutput[55]), 
        .A2(\Red_SubCellInst_LFInst_13_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst_LFInst_13_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst_LFInst_13_LFInst_2_U5  ( .A(PermutationOutput[53]), 
        .ZN(\Red_SubCellInst_LFInst_13_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_13_LFInst_2_U4  ( .A1(PermutationOutput[54]), .A2(\Red_SubCellInst_LFInst_13_LFInst_2_n13 ), .ZN(
        \Red_SubCellInst_LFInst_13_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst_LFInst_13_LFInst_2_U3  ( .A(PermutationOutput[52]), 
        .ZN(\Red_SubCellInst_LFInst_13_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_13_LFInst_3_U6  ( .A(PermutationOutput[53]), 
        .B(\Red_SubCellInst_LFInst_13_LFInst_3_n8 ), .ZN(Red_Feedback[55]) );
  NOR2_X1 \Red_SubCellInst_LFInst_13_LFInst_3_U5  ( .A1(
        \Red_SubCellInst_LFInst_13_LFInst_3_n7 ), .A2(
        \Red_SubCellInst_LFInst_13_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst_LFInst_13_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_13_LFInst_3_U4  ( .A1(PermutationOutput[54]), 
        .A2(PermutationOutput[55]), .ZN(
        \Red_SubCellInst_LFInst_13_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst_LFInst_13_LFInst_3_U3  ( .A1(PermutationOutput[55]), 
        .A2(PermutationOutput[52]), .ZN(
        \Red_SubCellInst_LFInst_13_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_14_LFInst_0_U10  ( .A1(
        \Red_SubCellInst_LFInst_14_LFInst_0_n14 ), .A2(
        \Red_SubCellInst_LFInst_14_LFInst_0_n13 ), .ZN(Red_Feedback[56]) );
  NAND2_X1 \Red_SubCellInst_LFInst_14_LFInst_0_U9  ( .A1(PermutationOutput[56]), .A2(\Red_SubCellInst_LFInst_14_LFInst_0_n12 ), .ZN(
        \Red_SubCellInst_LFInst_14_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_14_LFInst_0_U8  ( .A1(
        \Red_SubCellInst_LFInst_14_LFInst_0_n11 ), .A2(PermutationOutput[58]), 
        .ZN(\Red_SubCellInst_LFInst_14_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_14_LFInst_0_U7  ( .A(
        \Red_SubCellInst_LFInst_14_LFInst_0_n10 ), .B(
        \Red_SubCellInst_LFInst_14_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst_LFInst_14_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_14_LFInst_0_U6  ( .A1(PermutationOutput[59]), .A2(\Red_SubCellInst_LFInst_14_LFInst_0_n11 ), .ZN(
        \Red_SubCellInst_LFInst_14_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst_LFInst_14_LFInst_0_U5  ( .A(PermutationOutput[57]), 
        .ZN(\Red_SubCellInst_LFInst_14_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_14_LFInst_0_U4  ( .A1(PermutationOutput[58]), .A2(\Red_SubCellInst_LFInst_14_LFInst_0_n8 ), .ZN(
        \Red_SubCellInst_LFInst_14_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst_LFInst_14_LFInst_0_U3  ( .A(PermutationOutput[56]), 
        .ZN(\Red_SubCellInst_LFInst_14_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_14_LFInst_1_U8  ( .A1(
        \Red_SubCellInst_LFInst_14_LFInst_1_n15 ), .A2(
        \Red_SubCellInst_LFInst_14_LFInst_1_n14 ), .ZN(Red_Feedback[57]) );
  NAND2_X1 \Red_SubCellInst_LFInst_14_LFInst_1_U7  ( .A1(
        \Red_SubCellInst_LFInst_14_LFInst_1_n13 ), .A2(PermutationOutput[57]), 
        .ZN(\Red_SubCellInst_LFInst_14_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_14_LFInst_1_U6  ( .A1(
        \Red_SubCellInst_LFInst_14_LFInst_1_n12 ), .A2(PermutationOutput[56]), 
        .ZN(\Red_SubCellInst_LFInst_14_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_14_LFInst_1_U5  ( .A1(PermutationOutput[59]), .A2(PermutationOutput[58]), .ZN(\Red_SubCellInst_LFInst_14_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst_LFInst_14_LFInst_1_U4  ( .A1(PermutationOutput[58]), 
        .A2(\Red_SubCellInst_LFInst_14_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst_LFInst_14_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_14_LFInst_1_U3  ( .A(PermutationOutput[56]), 
        .B(PermutationOutput[59]), .ZN(
        \Red_SubCellInst_LFInst_14_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_14_LFInst_2_U10  ( .A1(
        \Red_SubCellInst_LFInst_14_LFInst_2_n19 ), .A2(
        \Red_SubCellInst_LFInst_14_LFInst_2_n18 ), .ZN(Red_Feedback[58]) );
  AND2_X1 \Red_SubCellInst_LFInst_14_LFInst_2_U9  ( .A1(
        \Red_SubCellInst_LFInst_14_LFInst_2_n17 ), .A2(PermutationOutput[56]), 
        .ZN(\Red_SubCellInst_LFInst_14_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_14_LFInst_2_U8  ( .A1(PermutationOutput[58]), 
        .A2(PermutationOutput[57]), .ZN(
        \Red_SubCellInst_LFInst_14_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_14_LFInst_2_U7  ( .A(
        \Red_SubCellInst_LFInst_14_LFInst_2_n16 ), .B(
        \Red_SubCellInst_LFInst_14_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst_LFInst_14_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_14_LFInst_2_U6  ( .A1(PermutationOutput[59]), 
        .A2(\Red_SubCellInst_LFInst_14_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst_LFInst_14_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst_LFInst_14_LFInst_2_U5  ( .A(PermutationOutput[57]), 
        .ZN(\Red_SubCellInst_LFInst_14_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_14_LFInst_2_U4  ( .A1(PermutationOutput[58]), .A2(\Red_SubCellInst_LFInst_14_LFInst_2_n13 ), .ZN(
        \Red_SubCellInst_LFInst_14_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst_LFInst_14_LFInst_2_U3  ( .A(PermutationOutput[56]), 
        .ZN(\Red_SubCellInst_LFInst_14_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_14_LFInst_3_U6  ( .A(PermutationOutput[57]), 
        .B(\Red_SubCellInst_LFInst_14_LFInst_3_n8 ), .ZN(Red_Feedback[59]) );
  NOR2_X1 \Red_SubCellInst_LFInst_14_LFInst_3_U5  ( .A1(
        \Red_SubCellInst_LFInst_14_LFInst_3_n7 ), .A2(
        \Red_SubCellInst_LFInst_14_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst_LFInst_14_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_14_LFInst_3_U4  ( .A1(PermutationOutput[58]), 
        .A2(PermutationOutput[59]), .ZN(
        \Red_SubCellInst_LFInst_14_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst_LFInst_14_LFInst_3_U3  ( .A1(PermutationOutput[59]), 
        .A2(PermutationOutput[56]), .ZN(
        \Red_SubCellInst_LFInst_14_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_15_LFInst_0_U10  ( .A1(
        \Red_SubCellInst_LFInst_15_LFInst_0_n14 ), .A2(
        \Red_SubCellInst_LFInst_15_LFInst_0_n13 ), .ZN(Red_Feedback[60]) );
  NAND2_X1 \Red_SubCellInst_LFInst_15_LFInst_0_U9  ( .A1(PermutationOutput[60]), .A2(\Red_SubCellInst_LFInst_15_LFInst_0_n12 ), .ZN(
        \Red_SubCellInst_LFInst_15_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_15_LFInst_0_U8  ( .A1(
        \Red_SubCellInst_LFInst_15_LFInst_0_n11 ), .A2(PermutationOutput[62]), 
        .ZN(\Red_SubCellInst_LFInst_15_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_15_LFInst_0_U7  ( .A(
        \Red_SubCellInst_LFInst_15_LFInst_0_n10 ), .B(
        \Red_SubCellInst_LFInst_15_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst_LFInst_15_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_15_LFInst_0_U6  ( .A1(PermutationOutput[63]), .A2(\Red_SubCellInst_LFInst_15_LFInst_0_n11 ), .ZN(
        \Red_SubCellInst_LFInst_15_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst_LFInst_15_LFInst_0_U5  ( .A(PermutationOutput[61]), 
        .ZN(\Red_SubCellInst_LFInst_15_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_15_LFInst_0_U4  ( .A1(PermutationOutput[62]), .A2(\Red_SubCellInst_LFInst_15_LFInst_0_n8 ), .ZN(
        \Red_SubCellInst_LFInst_15_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst_LFInst_15_LFInst_0_U3  ( .A(PermutationOutput[60]), 
        .ZN(\Red_SubCellInst_LFInst_15_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_15_LFInst_1_U8  ( .A1(
        \Red_SubCellInst_LFInst_15_LFInst_1_n15 ), .A2(
        \Red_SubCellInst_LFInst_15_LFInst_1_n14 ), .ZN(Red_Feedback[61]) );
  NAND2_X1 \Red_SubCellInst_LFInst_15_LFInst_1_U7  ( .A1(
        \Red_SubCellInst_LFInst_15_LFInst_1_n13 ), .A2(PermutationOutput[61]), 
        .ZN(\Red_SubCellInst_LFInst_15_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_15_LFInst_1_U6  ( .A1(
        \Red_SubCellInst_LFInst_15_LFInst_1_n12 ), .A2(PermutationOutput[60]), 
        .ZN(\Red_SubCellInst_LFInst_15_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_15_LFInst_1_U5  ( .A1(PermutationOutput[63]), .A2(PermutationOutput[62]), .ZN(\Red_SubCellInst_LFInst_15_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst_LFInst_15_LFInst_1_U4  ( .A1(PermutationOutput[62]), 
        .A2(\Red_SubCellInst_LFInst_15_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst_LFInst_15_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_15_LFInst_1_U3  ( .A(PermutationOutput[60]), 
        .B(PermutationOutput[63]), .ZN(
        \Red_SubCellInst_LFInst_15_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_15_LFInst_2_U10  ( .A1(
        \Red_SubCellInst_LFInst_15_LFInst_2_n19 ), .A2(
        \Red_SubCellInst_LFInst_15_LFInst_2_n18 ), .ZN(Red_Feedback[62]) );
  AND2_X1 \Red_SubCellInst_LFInst_15_LFInst_2_U9  ( .A1(
        \Red_SubCellInst_LFInst_15_LFInst_2_n17 ), .A2(PermutationOutput[60]), 
        .ZN(\Red_SubCellInst_LFInst_15_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_15_LFInst_2_U8  ( .A1(PermutationOutput[62]), 
        .A2(PermutationOutput[61]), .ZN(
        \Red_SubCellInst_LFInst_15_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_15_LFInst_2_U7  ( .A(
        \Red_SubCellInst_LFInst_15_LFInst_2_n16 ), .B(
        \Red_SubCellInst_LFInst_15_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst_LFInst_15_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_15_LFInst_2_U6  ( .A1(PermutationOutput[63]), 
        .A2(\Red_SubCellInst_LFInst_15_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst_LFInst_15_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst_LFInst_15_LFInst_2_U5  ( .A(PermutationOutput[61]), 
        .ZN(\Red_SubCellInst_LFInst_15_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst_LFInst_15_LFInst_2_U4  ( .A1(PermutationOutput[62]), .A2(\Red_SubCellInst_LFInst_15_LFInst_2_n13 ), .ZN(
        \Red_SubCellInst_LFInst_15_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst_LFInst_15_LFInst_2_U3  ( .A(PermutationOutput[60]), 
        .ZN(\Red_SubCellInst_LFInst_15_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst_LFInst_15_LFInst_3_U6  ( .A(PermutationOutput[61]), 
        .B(\Red_SubCellInst_LFInst_15_LFInst_3_n8 ), .ZN(Red_Feedback[63]) );
  NOR2_X1 \Red_SubCellInst_LFInst_15_LFInst_3_U5  ( .A1(
        \Red_SubCellInst_LFInst_15_LFInst_3_n7 ), .A2(
        \Red_SubCellInst_LFInst_15_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst_LFInst_15_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst_LFInst_15_LFInst_3_U4  ( .A1(PermutationOutput[62]), 
        .A2(PermutationOutput[63]), .ZN(
        \Red_SubCellInst_LFInst_15_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst_LFInst_15_LFInst_3_U3  ( .A1(PermutationOutput[63]), 
        .A2(PermutationOutput[60]), .ZN(
        \Red_SubCellInst_LFInst_15_LFInst_3_n7 ) );
  XNOR2_X1 \Red_MCInst2_XOR_r0_Inst_0_U2  ( .A(\Red_MCInst2_XOR_r0_Inst_0_n3 ), 
        .B(Red_MCOutput2[0]), .ZN(Red_MCOutput2[48]) );
  XNOR2_X1 \Red_MCInst2_XOR_r0_Inst_0_U1  ( .A(Red_Feedback[48]), .B(
        Red_MCOutput2[16]), .ZN(\Red_MCInst2_XOR_r0_Inst_0_n3 ) );
  XOR2_X1 \Red_MCInst2_XOR_r1_Inst_0_U1  ( .A(Red_Feedback[32]), .B(
        Red_MCOutput2[0]), .Z(Red_MCOutput2[32]) );
  XNOR2_X1 \Red_MCInst2_XOR_r0_Inst_1_U2  ( .A(\Red_MCInst2_XOR_r0_Inst_1_n3 ), 
        .B(Red_MCOutput2[1]), .ZN(Red_MCOutput2[49]) );
  XNOR2_X1 \Red_MCInst2_XOR_r0_Inst_1_U1  ( .A(Red_Feedback[49]), .B(
        Red_MCOutput2[17]), .ZN(\Red_MCInst2_XOR_r0_Inst_1_n3 ) );
  XOR2_X1 \Red_MCInst2_XOR_r1_Inst_1_U1  ( .A(Red_Feedback[33]), .B(
        Red_MCOutput2[1]), .Z(Red_MCOutput2[33]) );
  XNOR2_X1 \Red_MCInst2_XOR_r0_Inst_2_U2  ( .A(\Red_MCInst2_XOR_r0_Inst_2_n3 ), 
        .B(Red_MCOutput2[2]), .ZN(Red_MCOutput2[50]) );
  XNOR2_X1 \Red_MCInst2_XOR_r0_Inst_2_U1  ( .A(Red_Feedback[50]), .B(
        Red_MCOutput2[18]), .ZN(\Red_MCInst2_XOR_r0_Inst_2_n3 ) );
  XOR2_X1 \Red_MCInst2_XOR_r1_Inst_2_U1  ( .A(Red_Feedback[34]), .B(
        Red_MCOutput2[2]), .Z(Red_MCOutput2[34]) );
  XNOR2_X1 \Red_MCInst2_XOR_r0_Inst_3_U2  ( .A(\Red_MCInst2_XOR_r0_Inst_3_n3 ), 
        .B(Red_MCOutput2[3]), .ZN(Red_MCOutput2[51]) );
  XNOR2_X1 \Red_MCInst2_XOR_r0_Inst_3_U1  ( .A(Red_Feedback[51]), .B(
        Red_MCOutput2[19]), .ZN(\Red_MCInst2_XOR_r0_Inst_3_n3 ) );
  XOR2_X1 \Red_MCInst2_XOR_r1_Inst_3_U1  ( .A(Red_Feedback[35]), .B(
        Red_MCOutput2[3]), .Z(Red_MCOutput2[35]) );
  XNOR2_X1 \Red_MCInst2_XOR_r0_Inst_4_U2  ( .A(\Red_MCInst2_XOR_r0_Inst_4_n3 ), 
        .B(Red_MCOutput2[4]), .ZN(Red_MCOutput2[52]) );
  XNOR2_X1 \Red_MCInst2_XOR_r0_Inst_4_U1  ( .A(Red_Feedback[52]), .B(
        Red_MCOutput2[20]), .ZN(\Red_MCInst2_XOR_r0_Inst_4_n3 ) );
  XOR2_X1 \Red_MCInst2_XOR_r1_Inst_4_U1  ( .A(Red_Feedback[36]), .B(
        Red_MCOutput2[4]), .Z(Red_MCOutput2[36]) );
  XNOR2_X1 \Red_MCInst2_XOR_r0_Inst_5_U2  ( .A(\Red_MCInst2_XOR_r0_Inst_5_n3 ), 
        .B(Red_MCOutput2[5]), .ZN(Red_MCOutput2[53]) );
  XNOR2_X1 \Red_MCInst2_XOR_r0_Inst_5_U1  ( .A(Red_Feedback[53]), .B(
        Red_MCOutput2[21]), .ZN(\Red_MCInst2_XOR_r0_Inst_5_n3 ) );
  XOR2_X1 \Red_MCInst2_XOR_r1_Inst_5_U1  ( .A(Red_Feedback[37]), .B(
        Red_MCOutput2[5]), .Z(Red_MCOutput2[37]) );
  XNOR2_X1 \Red_MCInst2_XOR_r0_Inst_6_U2  ( .A(\Red_MCInst2_XOR_r0_Inst_6_n3 ), 
        .B(Red_MCOutput2[6]), .ZN(Red_MCOutput2[54]) );
  XNOR2_X1 \Red_MCInst2_XOR_r0_Inst_6_U1  ( .A(Red_Feedback[54]), .B(
        Red_MCOutput2[22]), .ZN(\Red_MCInst2_XOR_r0_Inst_6_n3 ) );
  XOR2_X1 \Red_MCInst2_XOR_r1_Inst_6_U1  ( .A(Red_Feedback[38]), .B(
        Red_MCOutput2[6]), .Z(Red_MCOutput2[38]) );
  XNOR2_X1 \Red_MCInst2_XOR_r0_Inst_7_U2  ( .A(\Red_MCInst2_XOR_r0_Inst_7_n3 ), 
        .B(Red_MCOutput2[7]), .ZN(Red_MCOutput2[55]) );
  XNOR2_X1 \Red_MCInst2_XOR_r0_Inst_7_U1  ( .A(Red_Feedback[55]), .B(
        Red_MCOutput2[23]), .ZN(\Red_MCInst2_XOR_r0_Inst_7_n3 ) );
  XOR2_X1 \Red_MCInst2_XOR_r1_Inst_7_U1  ( .A(Red_Feedback[39]), .B(
        Red_MCOutput2[7]), .Z(Red_MCOutput2[39]) );
  XNOR2_X1 \Red_MCInst2_XOR_r0_Inst_8_U2  ( .A(\Red_MCInst2_XOR_r0_Inst_8_n3 ), 
        .B(Red_MCOutput2[8]), .ZN(Red_MCOutput2[56]) );
  XNOR2_X1 \Red_MCInst2_XOR_r0_Inst_8_U1  ( .A(Red_Feedback[56]), .B(
        Red_MCOutput2[24]), .ZN(\Red_MCInst2_XOR_r0_Inst_8_n3 ) );
  XOR2_X1 \Red_MCInst2_XOR_r1_Inst_8_U1  ( .A(Red_Feedback[40]), .B(
        Red_MCOutput2[8]), .Z(Red_MCOutput2[40]) );
  XNOR2_X1 \Red_MCInst2_XOR_r0_Inst_9_U2  ( .A(\Red_MCInst2_XOR_r0_Inst_9_n3 ), 
        .B(Red_MCOutput2[9]), .ZN(Red_MCOutput2[57]) );
  XNOR2_X1 \Red_MCInst2_XOR_r0_Inst_9_U1  ( .A(Red_Feedback[57]), .B(
        Red_MCOutput2[25]), .ZN(\Red_MCInst2_XOR_r0_Inst_9_n3 ) );
  XOR2_X1 \Red_MCInst2_XOR_r1_Inst_9_U1  ( .A(Red_Feedback[41]), .B(
        Red_MCOutput2[9]), .Z(Red_MCOutput2[41]) );
  XNOR2_X1 \Red_MCInst2_XOR_r0_Inst_10_U2  ( .A(
        \Red_MCInst2_XOR_r0_Inst_10_n3 ), .B(Red_MCOutput2[10]), .ZN(
        Red_MCOutput2[58]) );
  XNOR2_X1 \Red_MCInst2_XOR_r0_Inst_10_U1  ( .A(Red_Feedback[58]), .B(
        Red_MCOutput2[26]), .ZN(\Red_MCInst2_XOR_r0_Inst_10_n3 ) );
  XOR2_X1 \Red_MCInst2_XOR_r1_Inst_10_U1  ( .A(Red_Feedback[42]), .B(
        Red_MCOutput2[10]), .Z(Red_MCOutput2[42]) );
  XNOR2_X1 \Red_MCInst2_XOR_r0_Inst_11_U2  ( .A(
        \Red_MCInst2_XOR_r0_Inst_11_n3 ), .B(Red_MCOutput2[11]), .ZN(
        Red_MCOutput2[59]) );
  XNOR2_X1 \Red_MCInst2_XOR_r0_Inst_11_U1  ( .A(Red_Feedback[59]), .B(
        Red_MCOutput2[27]), .ZN(\Red_MCInst2_XOR_r0_Inst_11_n3 ) );
  XOR2_X1 \Red_MCInst2_XOR_r1_Inst_11_U1  ( .A(Red_Feedback[43]), .B(
        Red_MCOutput2[11]), .Z(Red_MCOutput2[43]) );
  XNOR2_X1 \Red_MCInst2_XOR_r0_Inst_12_U2  ( .A(
        \Red_MCInst2_XOR_r0_Inst_12_n3 ), .B(Red_MCOutput2[12]), .ZN(
        Red_MCOutput2[60]) );
  XNOR2_X1 \Red_MCInst2_XOR_r0_Inst_12_U1  ( .A(Red_Feedback[60]), .B(
        Red_MCOutput2[28]), .ZN(\Red_MCInst2_XOR_r0_Inst_12_n3 ) );
  XOR2_X1 \Red_MCInst2_XOR_r1_Inst_12_U1  ( .A(Red_Feedback[44]), .B(
        Red_MCOutput2[12]), .Z(Red_MCOutput2[44]) );
  XNOR2_X1 \Red_MCInst2_XOR_r0_Inst_13_U2  ( .A(
        \Red_MCInst2_XOR_r0_Inst_13_n3 ), .B(Red_MCOutput2[13]), .ZN(
        Red_MCOutput2[61]) );
  XNOR2_X1 \Red_MCInst2_XOR_r0_Inst_13_U1  ( .A(Red_Feedback[61]), .B(
        Red_MCOutput2[29]), .ZN(\Red_MCInst2_XOR_r0_Inst_13_n3 ) );
  XOR2_X1 \Red_MCInst2_XOR_r1_Inst_13_U1  ( .A(Red_Feedback[45]), .B(
        Red_MCOutput2[13]), .Z(Red_MCOutput2[45]) );
  XNOR2_X1 \Red_MCInst2_XOR_r0_Inst_14_U2  ( .A(
        \Red_MCInst2_XOR_r0_Inst_14_n3 ), .B(Red_MCOutput2[14]), .ZN(
        Red_MCOutput2[62]) );
  XNOR2_X1 \Red_MCInst2_XOR_r0_Inst_14_U1  ( .A(Red_Feedback[62]), .B(
        Red_MCOutput2[30]), .ZN(\Red_MCInst2_XOR_r0_Inst_14_n3 ) );
  XOR2_X1 \Red_MCInst2_XOR_r1_Inst_14_U1  ( .A(Red_Feedback[46]), .B(
        Red_MCOutput2[14]), .Z(Red_MCOutput2[46]) );
  XNOR2_X1 \Red_MCInst2_XOR_r0_Inst_15_U2  ( .A(
        \Red_MCInst2_XOR_r0_Inst_15_n3 ), .B(Red_MCOutput2[15]), .ZN(
        Red_MCOutput2[63]) );
  XNOR2_X1 \Red_MCInst2_XOR_r0_Inst_15_U1  ( .A(Red_Feedback[63]), .B(
        Red_MCOutput2[31]), .ZN(\Red_MCInst2_XOR_r0_Inst_15_n3 ) );
  XOR2_X1 \Red_MCInst2_XOR_r1_Inst_15_U1  ( .A(Red_Feedback[47]), .B(
        Red_MCOutput2[15]), .Z(Red_MCOutput2[47]) );
  XOR2_X1 \Red_AddKeyXOR12_XORInst_0_0_U1  ( .A(Red_MCOutput2[48]), .B(
        Red_K1[48]), .Z(Red_AddRoundKeyOutput2[48]) );
  XOR2_X1 \Red_AddKeyXOR12_XORInst_0_1_U1  ( .A(Red_MCOutput2[49]), .B(
        Red_K1[49]), .Z(Red_AddRoundKeyOutput2[49]) );
  XOR2_X1 \Red_AddKeyXOR12_XORInst_0_2_U1  ( .A(Red_MCOutput2[50]), .B(
        Red_K1[50]), .Z(Red_AddRoundKeyOutput2[50]) );
  XOR2_X1 \Red_AddKeyXOR12_XORInst_0_3_U1  ( .A(Red_MCOutput2[51]), .B(
        Red_K1[51]), .Z(Red_AddRoundKeyOutput2[51]) );
  XOR2_X1 \Red_AddKeyXOR12_XORInst_1_0_U1  ( .A(Red_MCOutput2[52]), .B(
        Red_K1[52]), .Z(Red_AddRoundKeyOutput2[52]) );
  XOR2_X1 \Red_AddKeyXOR12_XORInst_1_1_U1  ( .A(Red_MCOutput2[53]), .B(
        Red_K1[53]), .Z(Red_AddRoundKeyOutput2[53]) );
  XOR2_X1 \Red_AddKeyXOR12_XORInst_1_2_U1  ( .A(Red_MCOutput2[54]), .B(
        Red_K1[54]), .Z(Red_AddRoundKeyOutput2[54]) );
  XOR2_X1 \Red_AddKeyXOR12_XORInst_1_3_U1  ( .A(Red_MCOutput2[55]), .B(
        Red_K1[55]), .Z(Red_AddRoundKeyOutput2[55]) );
  XOR2_X1 \Red_AddKeyXOR12_XORInst_2_0_U1  ( .A(Red_MCOutput2[56]), .B(
        Red_K1[56]), .Z(Red_AddRoundKeyOutput2[56]) );
  XOR2_X1 \Red_AddKeyXOR12_XORInst_2_1_U1  ( .A(Red_MCOutput2[57]), .B(
        Red_K1[57]), .Z(Red_AddRoundKeyOutput2[57]) );
  XOR2_X1 \Red_AddKeyXOR12_XORInst_2_2_U1  ( .A(Red_MCOutput2[58]), .B(
        Red_K1[58]), .Z(Red_AddRoundKeyOutput2[58]) );
  XOR2_X1 \Red_AddKeyXOR12_XORInst_2_3_U1  ( .A(Red_MCOutput2[59]), .B(
        Red_K1[59]), .Z(Red_AddRoundKeyOutput2[59]) );
  XOR2_X1 \Red_AddKeyXOR12_XORInst_3_0_U1  ( .A(Red_MCOutput2[60]), .B(
        Red_K1[60]), .Z(Red_AddRoundKeyOutput2[60]) );
  XOR2_X1 \Red_AddKeyXOR12_XORInst_3_1_U1  ( .A(Red_MCOutput2[61]), .B(
        Red_K1[61]), .Z(Red_AddRoundKeyOutput2[61]) );
  XOR2_X1 \Red_AddKeyXOR12_XORInst_3_2_U1  ( .A(Red_MCOutput2[62]), .B(
        Red_K1[62]), .Z(Red_AddRoundKeyOutput2[62]) );
  XOR2_X1 \Red_AddKeyXOR12_XORInst_3_3_U1  ( .A(Red_MCOutput2[63]), .B(
        Red_K1[63]), .Z(Red_AddRoundKeyOutput2[63]) );
  XOR2_X1 \Red_AddKeyConstXOR2_XORInst_0_0_U1  ( .A(Red_K1[40]), .B(
        Red_MCOutput2[40]), .Z(Red_AddRoundKeyOutput2[40]) );
  XOR2_X1 \Red_AddKeyConstXOR2_XORInst_0_1_U1  ( .A(Red_K1[41]), .B(
        Red_MCOutput2[41]), .Z(Red_AddRoundKeyOutput2[41]) );
  XOR2_X1 \Red_AddKeyConstXOR2_XORInst_0_2_U1  ( .A(Red_K1[42]), .B(
        Red_MCOutput2[42]), .Z(Red_AddRoundKeyOutput2[42]) );
  XOR2_X1 \Red_AddKeyConstXOR2_XORInst_0_3_U1  ( .A(Red_K1[43]), .B(
        Red_MCOutput2[43]), .Z(Red_AddRoundKeyOutput2[43]) );
  XOR2_X1 \Red_AddKeyConstXOR2_XORInst_1_0_U1  ( .A(Red_K1[44]), .B(
        Red_MCOutput2[44]), .Z(Red_AddRoundKeyOutput2[44]) );
  XOR2_X1 \Red_AddKeyConstXOR2_XORInst_1_1_U1  ( .A(Red_K1[45]), .B(
        Red_MCOutput2[45]), .Z(Red_AddRoundKeyOutput2[45]) );
  XOR2_X1 \Red_AddKeyConstXOR2_XORInst_1_2_U1  ( .A(Red_K1[46]), .B(
        Red_MCOutput2[46]), .Z(Red_AddRoundKeyOutput2[46]) );
  XOR2_X1 \Red_AddKeyConstXOR2_XORInst_1_3_U1  ( .A(Red_K1[47]), .B(
        Red_MCOutput2[47]), .Z(Red_AddRoundKeyOutput2[47]) );
  XOR2_X1 \Red_AddKeyXOR22_XORInst_0_0_U1  ( .A(Red_MCOutput2[0]), .B(
        Red_K1[0]), .Z(Red_AddRoundKeyOutput2[0]) );
  XOR2_X1 \Red_AddKeyXOR22_XORInst_0_1_U1  ( .A(Red_MCOutput2[1]), .B(
        Red_K1[1]), .Z(Red_AddRoundKeyOutput2[1]) );
  XOR2_X1 \Red_AddKeyXOR22_XORInst_0_2_U1  ( .A(Red_MCOutput2[2]), .B(
        Red_K1[2]), .Z(Red_AddRoundKeyOutput2[2]) );
  XOR2_X1 \Red_AddKeyXOR22_XORInst_0_3_U1  ( .A(Red_MCOutput2[3]), .B(
        Red_K1[3]), .Z(Red_AddRoundKeyOutput2[3]) );
  XOR2_X1 \Red_AddKeyXOR22_XORInst_1_0_U1  ( .A(Red_MCOutput2[4]), .B(
        Red_K1[4]), .Z(Red_AddRoundKeyOutput2[4]) );
  XOR2_X1 \Red_AddKeyXOR22_XORInst_1_1_U1  ( .A(Red_MCOutput2[5]), .B(
        Red_K1[5]), .Z(Red_AddRoundKeyOutput2[5]) );
  XOR2_X1 \Red_AddKeyXOR22_XORInst_1_2_U1  ( .A(Red_MCOutput2[6]), .B(
        Red_K1[6]), .Z(Red_AddRoundKeyOutput2[6]) );
  XOR2_X1 \Red_AddKeyXOR22_XORInst_1_3_U1  ( .A(Red_MCOutput2[7]), .B(
        Red_K1[7]), .Z(Red_AddRoundKeyOutput2[7]) );
  XOR2_X1 \Red_AddKeyXOR22_XORInst_2_0_U1  ( .A(Red_MCOutput2[8]), .B(
        Red_K1[8]), .Z(Red_AddRoundKeyOutput2[8]) );
  XOR2_X1 \Red_AddKeyXOR22_XORInst_2_1_U1  ( .A(Red_MCOutput2[9]), .B(
        Red_K1[9]), .Z(Red_AddRoundKeyOutput2[9]) );
  XOR2_X1 \Red_AddKeyXOR22_XORInst_2_2_U1  ( .A(Red_MCOutput2[10]), .B(
        Red_K1[10]), .Z(Red_AddRoundKeyOutput2[10]) );
  XOR2_X1 \Red_AddKeyXOR22_XORInst_2_3_U1  ( .A(Red_MCOutput2[11]), .B(
        Red_K1[11]), .Z(Red_AddRoundKeyOutput2[11]) );
  XOR2_X1 \Red_AddKeyXOR22_XORInst_3_0_U1  ( .A(Red_MCOutput2[12]), .B(
        Red_K1[12]), .Z(Red_AddRoundKeyOutput2[12]) );
  XOR2_X1 \Red_AddKeyXOR22_XORInst_3_1_U1  ( .A(Red_MCOutput2[13]), .B(
        Red_K1[13]), .Z(Red_AddRoundKeyOutput2[13]) );
  XOR2_X1 \Red_AddKeyXOR22_XORInst_3_2_U1  ( .A(Red_MCOutput2[14]), .B(
        Red_K1[14]), .Z(Red_AddRoundKeyOutput2[14]) );
  XOR2_X1 \Red_AddKeyXOR22_XORInst_3_3_U1  ( .A(Red_MCOutput2[15]), .B(
        Red_K1[15]), .Z(Red_AddRoundKeyOutput2[15]) );
  XOR2_X1 \Red_AddKeyXOR22_XORInst_4_0_U1  ( .A(Red_MCOutput2[16]), .B(
        Red_K1[16]), .Z(Red_AddRoundKeyOutput2[16]) );
  XOR2_X1 \Red_AddKeyXOR22_XORInst_4_1_U1  ( .A(Red_MCOutput2[17]), .B(
        Red_K1[17]), .Z(Red_AddRoundKeyOutput2[17]) );
  XOR2_X1 \Red_AddKeyXOR22_XORInst_4_2_U1  ( .A(Red_MCOutput2[18]), .B(
        Red_K1[18]), .Z(Red_AddRoundKeyOutput2[18]) );
  XOR2_X1 \Red_AddKeyXOR22_XORInst_4_3_U1  ( .A(Red_MCOutput2[19]), .B(
        Red_K1[19]), .Z(Red_AddRoundKeyOutput2[19]) );
  XOR2_X1 \Red_AddKeyXOR22_XORInst_5_0_U1  ( .A(Red_MCOutput2[20]), .B(
        Red_K1[20]), .Z(Red_AddRoundKeyOutput2[20]) );
  XOR2_X1 \Red_AddKeyXOR22_XORInst_5_1_U1  ( .A(Red_MCOutput2[21]), .B(
        Red_K1[21]), .Z(Red_AddRoundKeyOutput2[21]) );
  XOR2_X1 \Red_AddKeyXOR22_XORInst_5_2_U1  ( .A(Red_MCOutput2[22]), .B(
        Red_K1[22]), .Z(Red_AddRoundKeyOutput2[22]) );
  XOR2_X1 \Red_AddKeyXOR22_XORInst_5_3_U1  ( .A(Red_MCOutput2[23]), .B(
        Red_K1[23]), .Z(Red_AddRoundKeyOutput2[23]) );
  XOR2_X1 \Red_AddKeyXOR22_XORInst_6_0_U1  ( .A(Red_MCOutput2[24]), .B(
        Red_K1[24]), .Z(Red_AddRoundKeyOutput2[24]) );
  XOR2_X1 \Red_AddKeyXOR22_XORInst_6_1_U1  ( .A(Red_MCOutput2[25]), .B(
        Red_K1[25]), .Z(Red_AddRoundKeyOutput2[25]) );
  XOR2_X1 \Red_AddKeyXOR22_XORInst_6_2_U1  ( .A(Red_MCOutput2[26]), .B(
        Red_K1[26]), .Z(Red_AddRoundKeyOutput2[26]) );
  XOR2_X1 \Red_AddKeyXOR22_XORInst_6_3_U1  ( .A(Red_MCOutput2[27]), .B(
        Red_K1[27]), .Z(Red_AddRoundKeyOutput2[27]) );
  XOR2_X1 \Red_AddKeyXOR22_XORInst_7_0_U1  ( .A(Red_MCOutput2[28]), .B(
        Red_K1[28]), .Z(Red_AddRoundKeyOutput2[28]) );
  XOR2_X1 \Red_AddKeyXOR22_XORInst_7_1_U1  ( .A(Red_MCOutput2[29]), .B(
        Red_K1[29]), .Z(Red_AddRoundKeyOutput2[29]) );
  XOR2_X1 \Red_AddKeyXOR22_XORInst_7_2_U1  ( .A(Red_MCOutput2[30]), .B(
        Red_K1[30]), .Z(Red_AddRoundKeyOutput2[30]) );
  XOR2_X1 \Red_AddKeyXOR22_XORInst_7_3_U1  ( .A(Red_MCOutput2[31]), .B(
        Red_K1[31]), .Z(Red_AddRoundKeyOutput2[31]) );
  XOR2_X1 \Red_AddKeyXOR22_XORInst_8_0_U1  ( .A(Red_MCOutput2[32]), .B(
        Red_K1[32]), .Z(Red_AddRoundKeyOutput2[32]) );
  XOR2_X1 \Red_AddKeyXOR22_XORInst_8_1_U1  ( .A(Red_MCOutput2[33]), .B(
        Red_K1[33]), .Z(Red_AddRoundKeyOutput2[33]) );
  XOR2_X1 \Red_AddKeyXOR22_XORInst_8_2_U1  ( .A(Red_MCOutput2[34]), .B(
        Red_K1[34]), .Z(Red_AddRoundKeyOutput2[34]) );
  XOR2_X1 \Red_AddKeyXOR22_XORInst_8_3_U1  ( .A(Red_MCOutput2[35]), .B(
        Red_K1[35]), .Z(Red_AddRoundKeyOutput2[35]) );
  XOR2_X1 \Red_AddKeyXOR22_XORInst_9_0_U1  ( .A(Red_MCOutput2[36]), .B(
        Red_K1[36]), .Z(Red_AddRoundKeyOutput2[36]) );
  XOR2_X1 \Red_AddKeyXOR22_XORInst_9_1_U1  ( .A(Red_MCOutput2[37]), .B(
        Red_K1[37]), .Z(Red_AddRoundKeyOutput2[37]) );
  XOR2_X1 \Red_AddKeyXOR22_XORInst_9_2_U1  ( .A(Red_MCOutput2[38]), .B(
        Red_K1[38]), .Z(Red_AddRoundKeyOutput2[38]) );
  XOR2_X1 \Red_AddKeyXOR22_XORInst_9_3_U1  ( .A(Red_MCOutput2[39]), .B(
        Red_K1[39]), .Z(Red_AddRoundKeyOutput2[39]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[0]  ( .D(Red_AddRoundKeyOutput2[0]), .CK(clk), .Q(Red_StateRegOutput2[0]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[1]  ( .D(Red_AddRoundKeyOutput2[1]), .CK(clk), .Q(Red_StateRegOutput2[1]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[2]  ( .D(Red_AddRoundKeyOutput2[2]), .CK(clk), .Q(Red_StateRegOutput2[2]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[3]  ( .D(Red_AddRoundKeyOutput2[3]), .CK(clk), .Q(Red_StateRegOutput2[3]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[4]  ( .D(Red_AddRoundKeyOutput2[4]), .CK(clk), .Q(Red_StateRegOutput2[4]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[5]  ( .D(Red_AddRoundKeyOutput2[5]), .CK(clk), .Q(Red_StateRegOutput2[5]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[6]  ( .D(Red_AddRoundKeyOutput2[6]), .CK(clk), .Q(Red_StateRegOutput2[6]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[7]  ( .D(Red_AddRoundKeyOutput2[7]), .CK(clk), .Q(Red_StateRegOutput2[7]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[8]  ( .D(Red_AddRoundKeyOutput2[8]), .CK(clk), .Q(Red_StateRegOutput2[8]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[9]  ( .D(Red_AddRoundKeyOutput2[9]), .CK(clk), .Q(Red_StateRegOutput2[9]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[10]  ( .D(
        Red_AddRoundKeyOutput2[10]), .CK(clk), .Q(Red_StateRegOutput2[10]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[11]  ( .D(
        Red_AddRoundKeyOutput2[11]), .CK(clk), .Q(Red_StateRegOutput2[11]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[12]  ( .D(
        Red_AddRoundKeyOutput2[12]), .CK(clk), .Q(Red_StateRegOutput2[12]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[13]  ( .D(
        Red_AddRoundKeyOutput2[13]), .CK(clk), .Q(Red_StateRegOutput2[13]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[14]  ( .D(
        Red_AddRoundKeyOutput2[14]), .CK(clk), .Q(Red_StateRegOutput2[14]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[15]  ( .D(
        Red_AddRoundKeyOutput2[15]), .CK(clk), .Q(Red_StateRegOutput2[15]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[16]  ( .D(
        Red_AddRoundKeyOutput2[16]), .CK(clk), .Q(Red_StateRegOutput2[16]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[17]  ( .D(
        Red_AddRoundKeyOutput2[17]), .CK(clk), .Q(Red_StateRegOutput2[17]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[18]  ( .D(
        Red_AddRoundKeyOutput2[18]), .CK(clk), .Q(Red_StateRegOutput2[18]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[19]  ( .D(
        Red_AddRoundKeyOutput2[19]), .CK(clk), .Q(Red_StateRegOutput2[19]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[20]  ( .D(
        Red_AddRoundKeyOutput2[20]), .CK(clk), .Q(Red_StateRegOutput2[20]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[21]  ( .D(
        Red_AddRoundKeyOutput2[21]), .CK(clk), .Q(Red_StateRegOutput2[21]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[22]  ( .D(
        Red_AddRoundKeyOutput2[22]), .CK(clk), .Q(Red_StateRegOutput2[22]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[23]  ( .D(
        Red_AddRoundKeyOutput2[23]), .CK(clk), .Q(Red_StateRegOutput2[23]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[24]  ( .D(
        Red_AddRoundKeyOutput2[24]), .CK(clk), .Q(Red_StateRegOutput2[24]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[25]  ( .D(
        Red_AddRoundKeyOutput2[25]), .CK(clk), .Q(Red_StateRegOutput2[25]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[26]  ( .D(
        Red_AddRoundKeyOutput2[26]), .CK(clk), .Q(Red_StateRegOutput2[26]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[27]  ( .D(
        Red_AddRoundKeyOutput2[27]), .CK(clk), .Q(Red_StateRegOutput2[27]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[28]  ( .D(
        Red_AddRoundKeyOutput2[28]), .CK(clk), .Q(Red_StateRegOutput2[28]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[29]  ( .D(
        Red_AddRoundKeyOutput2[29]), .CK(clk), .Q(Red_StateRegOutput2[29]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[30]  ( .D(
        Red_AddRoundKeyOutput2[30]), .CK(clk), .Q(Red_StateRegOutput2[30]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[31]  ( .D(
        Red_AddRoundKeyOutput2[31]), .CK(clk), .Q(Red_StateRegOutput2[31]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[32]  ( .D(
        Red_AddRoundKeyOutput2[32]), .CK(clk), .Q(Red_StateRegOutput2[32]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[33]  ( .D(
        Red_AddRoundKeyOutput2[33]), .CK(clk), .Q(Red_StateRegOutput2[33]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[34]  ( .D(
        Red_AddRoundKeyOutput2[34]), .CK(clk), .Q(Red_StateRegOutput2[34]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[35]  ( .D(
        Red_AddRoundKeyOutput2[35]), .CK(clk), .Q(Red_StateRegOutput2[35]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[36]  ( .D(
        Red_AddRoundKeyOutput2[36]), .CK(clk), .Q(Red_StateRegOutput2[36]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[37]  ( .D(
        Red_AddRoundKeyOutput2[37]), .CK(clk), .Q(Red_StateRegOutput2[37]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[38]  ( .D(
        Red_AddRoundKeyOutput2[38]), .CK(clk), .Q(Red_StateRegOutput2[38]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[39]  ( .D(
        Red_AddRoundKeyOutput2[39]), .CK(clk), .Q(Red_StateRegOutput2[39]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[40]  ( .D(
        Red_AddRoundKeyOutput2[40]), .CK(clk), .Q(Red_StateRegOutput2[40]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[41]  ( .D(
        Red_AddRoundKeyOutput2[41]), .CK(clk), .Q(Red_StateRegOutput2[41]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[42]  ( .D(
        Red_AddRoundKeyOutput2[42]), .CK(clk), .Q(Red_StateRegOutput2[42]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[43]  ( .D(
        Red_AddRoundKeyOutput2[43]), .CK(clk), .Q(Red_StateRegOutput2[43]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[44]  ( .D(
        Red_AddRoundKeyOutput2[44]), .CK(clk), .Q(Red_StateRegOutput2[44]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[45]  ( .D(
        Red_AddRoundKeyOutput2[45]), .CK(clk), .Q(Red_StateRegOutput2[45]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[46]  ( .D(
        Red_AddRoundKeyOutput2[46]), .CK(clk), .Q(Red_StateRegOutput2[46]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[47]  ( .D(
        Red_AddRoundKeyOutput2[47]), .CK(clk), .Q(Red_StateRegOutput2[47]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[48]  ( .D(
        Red_AddRoundKeyOutput2[48]), .CK(clk), .Q(Red_StateRegOutput2[48]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[49]  ( .D(
        Red_AddRoundKeyOutput2[49]), .CK(clk), .Q(Red_StateRegOutput2[49]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[50]  ( .D(
        Red_AddRoundKeyOutput2[50]), .CK(clk), .Q(Red_StateRegOutput2[50]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[51]  ( .D(
        Red_AddRoundKeyOutput2[51]), .CK(clk), .Q(Red_StateRegOutput2[51]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[52]  ( .D(
        Red_AddRoundKeyOutput2[52]), .CK(clk), .Q(Red_StateRegOutput2[52]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[53]  ( .D(
        Red_AddRoundKeyOutput2[53]), .CK(clk), .Q(Red_StateRegOutput2[53]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[54]  ( .D(
        Red_AddRoundKeyOutput2[54]), .CK(clk), .Q(Red_StateRegOutput2[54]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[55]  ( .D(
        Red_AddRoundKeyOutput2[55]), .CK(clk), .Q(Red_StateRegOutput2[55]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[56]  ( .D(
        Red_AddRoundKeyOutput2[56]), .CK(clk), .Q(Red_StateRegOutput2[56]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[57]  ( .D(
        Red_AddRoundKeyOutput2[57]), .CK(clk), .Q(Red_StateRegOutput2[57]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[58]  ( .D(
        Red_AddRoundKeyOutput2[58]), .CK(clk), .Q(Red_StateRegOutput2[58]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[59]  ( .D(
        Red_AddRoundKeyOutput2[59]), .CK(clk), .Q(Red_StateRegOutput2[59]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[60]  ( .D(
        Red_AddRoundKeyOutput2[60]), .CK(clk), .Q(Red_StateRegOutput2[60]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[61]  ( .D(
        Red_AddRoundKeyOutput2[61]), .CK(clk), .Q(Red_StateRegOutput2[61]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[62]  ( .D(
        Red_AddRoundKeyOutput2[62]), .CK(clk), .Q(Red_StateRegOutput2[62]) );
  DFF_X1 \Red_StateReg2_s_current_state_reg[63]  ( .D(
        Red_AddRoundKeyOutput2[63]), .CK(clk), .Q(Red_StateRegOutput2[63]) );
  NAND2_X1 \Red_SubCellInst2_LFInst_0_LFInst_0_U10  ( .A1(
        \Red_SubCellInst2_LFInst_0_LFInst_0_n14 ), .A2(
        \Red_SubCellInst2_LFInst_0_LFInst_0_n13 ), .ZN(Red_MCOutput3[0]) );
  NAND2_X1 \Red_SubCellInst2_LFInst_0_LFInst_0_U9  ( .A1(PermutationOutput2[0]), .A2(\Red_SubCellInst2_LFInst_0_LFInst_0_n12 ), .ZN(
        \Red_SubCellInst2_LFInst_0_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_0_LFInst_0_U8  ( .A1(
        \Red_SubCellInst2_LFInst_0_LFInst_0_n11 ), .A2(PermutationOutput2[2]), 
        .ZN(\Red_SubCellInst2_LFInst_0_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_0_LFInst_0_U7  ( .A(
        \Red_SubCellInst2_LFInst_0_LFInst_0_n10 ), .B(
        \Red_SubCellInst2_LFInst_0_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst2_LFInst_0_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_0_LFInst_0_U6  ( .A1(PermutationOutput2[3]), .A2(\Red_SubCellInst2_LFInst_0_LFInst_0_n11 ), .ZN(
        \Red_SubCellInst2_LFInst_0_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst2_LFInst_0_LFInst_0_U5  ( .A(PermutationOutput2[1]), 
        .ZN(\Red_SubCellInst2_LFInst_0_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_0_LFInst_0_U4  ( .A1(PermutationOutput2[2]), .A2(\Red_SubCellInst2_LFInst_0_LFInst_0_n8 ), .ZN(
        \Red_SubCellInst2_LFInst_0_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst2_LFInst_0_LFInst_0_U3  ( .A(PermutationOutput2[0]), 
        .ZN(\Red_SubCellInst2_LFInst_0_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_0_LFInst_1_U8  ( .A1(
        \Red_SubCellInst2_LFInst_0_LFInst_1_n15 ), .A2(
        \Red_SubCellInst2_LFInst_0_LFInst_1_n14 ), .ZN(Red_MCOutput3[1]) );
  NAND2_X1 \Red_SubCellInst2_LFInst_0_LFInst_1_U7  ( .A1(
        \Red_SubCellInst2_LFInst_0_LFInst_1_n13 ), .A2(PermutationOutput2[1]), 
        .ZN(\Red_SubCellInst2_LFInst_0_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_0_LFInst_1_U6  ( .A1(
        \Red_SubCellInst2_LFInst_0_LFInst_1_n12 ), .A2(PermutationOutput2[0]), 
        .ZN(\Red_SubCellInst2_LFInst_0_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_0_LFInst_1_U5  ( .A1(PermutationOutput2[3]), .A2(PermutationOutput2[2]), .ZN(\Red_SubCellInst2_LFInst_0_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst2_LFInst_0_LFInst_1_U4  ( .A1(PermutationOutput2[2]), 
        .A2(\Red_SubCellInst2_LFInst_0_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst2_LFInst_0_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_0_LFInst_1_U3  ( .A(PermutationOutput2[0]), 
        .B(PermutationOutput2[3]), .ZN(
        \Red_SubCellInst2_LFInst_0_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_0_LFInst_2_U10  ( .A1(
        \Red_SubCellInst2_LFInst_0_LFInst_2_n19 ), .A2(
        \Red_SubCellInst2_LFInst_0_LFInst_2_n18 ), .ZN(Red_MCOutput3[2]) );
  AND2_X1 \Red_SubCellInst2_LFInst_0_LFInst_2_U9  ( .A1(
        \Red_SubCellInst2_LFInst_0_LFInst_2_n17 ), .A2(PermutationOutput2[0]), 
        .ZN(\Red_SubCellInst2_LFInst_0_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_0_LFInst_2_U8  ( .A1(PermutationOutput2[2]), 
        .A2(PermutationOutput2[1]), .ZN(
        \Red_SubCellInst2_LFInst_0_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_0_LFInst_2_U7  ( .A(
        \Red_SubCellInst2_LFInst_0_LFInst_2_n16 ), .B(
        \Red_SubCellInst2_LFInst_0_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst2_LFInst_0_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_0_LFInst_2_U6  ( .A1(PermutationOutput2[3]), 
        .A2(\Red_SubCellInst2_LFInst_0_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst2_LFInst_0_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst2_LFInst_0_LFInst_2_U5  ( .A(PermutationOutput2[1]), 
        .ZN(\Red_SubCellInst2_LFInst_0_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_0_LFInst_2_U4  ( .A1(PermutationOutput2[2]), .A2(\Red_SubCellInst2_LFInst_0_LFInst_2_n13 ), .ZN(
        \Red_SubCellInst2_LFInst_0_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst2_LFInst_0_LFInst_2_U3  ( .A(PermutationOutput2[0]), 
        .ZN(\Red_SubCellInst2_LFInst_0_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_0_LFInst_3_U6  ( .A(PermutationOutput2[1]), 
        .B(\Red_SubCellInst2_LFInst_0_LFInst_3_n8 ), .ZN(Red_MCOutput3[3]) );
  NOR2_X1 \Red_SubCellInst2_LFInst_0_LFInst_3_U5  ( .A1(
        \Red_SubCellInst2_LFInst_0_LFInst_3_n7 ), .A2(
        \Red_SubCellInst2_LFInst_0_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst2_LFInst_0_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_0_LFInst_3_U4  ( .A1(PermutationOutput2[2]), 
        .A2(PermutationOutput2[3]), .ZN(
        \Red_SubCellInst2_LFInst_0_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst2_LFInst_0_LFInst_3_U3  ( .A1(PermutationOutput2[3]), 
        .A2(PermutationOutput2[0]), .ZN(
        \Red_SubCellInst2_LFInst_0_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_1_LFInst_0_U10  ( .A1(
        \Red_SubCellInst2_LFInst_1_LFInst_0_n14 ), .A2(
        \Red_SubCellInst2_LFInst_1_LFInst_0_n13 ), .ZN(Red_MCOutput3[4]) );
  NAND2_X1 \Red_SubCellInst2_LFInst_1_LFInst_0_U9  ( .A1(PermutationOutput2[4]), .A2(\Red_SubCellInst2_LFInst_1_LFInst_0_n12 ), .ZN(
        \Red_SubCellInst2_LFInst_1_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_1_LFInst_0_U8  ( .A1(
        \Red_SubCellInst2_LFInst_1_LFInst_0_n11 ), .A2(PermutationOutput2[6]), 
        .ZN(\Red_SubCellInst2_LFInst_1_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_1_LFInst_0_U7  ( .A(
        \Red_SubCellInst2_LFInst_1_LFInst_0_n10 ), .B(
        \Red_SubCellInst2_LFInst_1_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst2_LFInst_1_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_1_LFInst_0_U6  ( .A1(PermutationOutput2[7]), .A2(\Red_SubCellInst2_LFInst_1_LFInst_0_n11 ), .ZN(
        \Red_SubCellInst2_LFInst_1_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst2_LFInst_1_LFInst_0_U5  ( .A(PermutationOutput2[5]), 
        .ZN(\Red_SubCellInst2_LFInst_1_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_1_LFInst_0_U4  ( .A1(PermutationOutput2[6]), .A2(\Red_SubCellInst2_LFInst_1_LFInst_0_n8 ), .ZN(
        \Red_SubCellInst2_LFInst_1_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst2_LFInst_1_LFInst_0_U3  ( .A(PermutationOutput2[4]), 
        .ZN(\Red_SubCellInst2_LFInst_1_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_1_LFInst_1_U8  ( .A1(
        \Red_SubCellInst2_LFInst_1_LFInst_1_n15 ), .A2(
        \Red_SubCellInst2_LFInst_1_LFInst_1_n14 ), .ZN(Red_MCOutput3[5]) );
  NAND2_X1 \Red_SubCellInst2_LFInst_1_LFInst_1_U7  ( .A1(
        \Red_SubCellInst2_LFInst_1_LFInst_1_n13 ), .A2(PermutationOutput2[5]), 
        .ZN(\Red_SubCellInst2_LFInst_1_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_1_LFInst_1_U6  ( .A1(
        \Red_SubCellInst2_LFInst_1_LFInst_1_n12 ), .A2(PermutationOutput2[4]), 
        .ZN(\Red_SubCellInst2_LFInst_1_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_1_LFInst_1_U5  ( .A1(PermutationOutput2[7]), .A2(PermutationOutput2[6]), .ZN(\Red_SubCellInst2_LFInst_1_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst2_LFInst_1_LFInst_1_U4  ( .A1(PermutationOutput2[6]), 
        .A2(\Red_SubCellInst2_LFInst_1_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst2_LFInst_1_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_1_LFInst_1_U3  ( .A(PermutationOutput2[4]), 
        .B(PermutationOutput2[7]), .ZN(
        \Red_SubCellInst2_LFInst_1_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_1_LFInst_2_U10  ( .A1(
        \Red_SubCellInst2_LFInst_1_LFInst_2_n19 ), .A2(
        \Red_SubCellInst2_LFInst_1_LFInst_2_n18 ), .ZN(Red_MCOutput3[6]) );
  AND2_X1 \Red_SubCellInst2_LFInst_1_LFInst_2_U9  ( .A1(
        \Red_SubCellInst2_LFInst_1_LFInst_2_n17 ), .A2(PermutationOutput2[4]), 
        .ZN(\Red_SubCellInst2_LFInst_1_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_1_LFInst_2_U8  ( .A1(PermutationOutput2[6]), 
        .A2(PermutationOutput2[5]), .ZN(
        \Red_SubCellInst2_LFInst_1_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_1_LFInst_2_U7  ( .A(
        \Red_SubCellInst2_LFInst_1_LFInst_2_n16 ), .B(
        \Red_SubCellInst2_LFInst_1_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst2_LFInst_1_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_1_LFInst_2_U6  ( .A1(PermutationOutput2[7]), 
        .A2(\Red_SubCellInst2_LFInst_1_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst2_LFInst_1_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst2_LFInst_1_LFInst_2_U5  ( .A(PermutationOutput2[5]), 
        .ZN(\Red_SubCellInst2_LFInst_1_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_1_LFInst_2_U4  ( .A1(PermutationOutput2[6]), .A2(\Red_SubCellInst2_LFInst_1_LFInst_2_n13 ), .ZN(
        \Red_SubCellInst2_LFInst_1_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst2_LFInst_1_LFInst_2_U3  ( .A(PermutationOutput2[4]), 
        .ZN(\Red_SubCellInst2_LFInst_1_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_1_LFInst_3_U6  ( .A(PermutationOutput2[5]), 
        .B(\Red_SubCellInst2_LFInst_1_LFInst_3_n8 ), .ZN(Red_MCOutput3[7]) );
  NOR2_X1 \Red_SubCellInst2_LFInst_1_LFInst_3_U5  ( .A1(
        \Red_SubCellInst2_LFInst_1_LFInst_3_n7 ), .A2(
        \Red_SubCellInst2_LFInst_1_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst2_LFInst_1_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_1_LFInst_3_U4  ( .A1(PermutationOutput2[6]), 
        .A2(PermutationOutput2[7]), .ZN(
        \Red_SubCellInst2_LFInst_1_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst2_LFInst_1_LFInst_3_U3  ( .A1(PermutationOutput2[7]), 
        .A2(PermutationOutput2[4]), .ZN(
        \Red_SubCellInst2_LFInst_1_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_2_LFInst_0_U10  ( .A1(
        \Red_SubCellInst2_LFInst_2_LFInst_0_n14 ), .A2(
        \Red_SubCellInst2_LFInst_2_LFInst_0_n13 ), .ZN(Red_MCOutput3[8]) );
  NAND2_X1 \Red_SubCellInst2_LFInst_2_LFInst_0_U9  ( .A1(PermutationOutput2[8]), .A2(\Red_SubCellInst2_LFInst_2_LFInst_0_n12 ), .ZN(
        \Red_SubCellInst2_LFInst_2_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_2_LFInst_0_U8  ( .A1(
        \Red_SubCellInst2_LFInst_2_LFInst_0_n11 ), .A2(PermutationOutput2[10]), 
        .ZN(\Red_SubCellInst2_LFInst_2_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_2_LFInst_0_U7  ( .A(
        \Red_SubCellInst2_LFInst_2_LFInst_0_n10 ), .B(
        \Red_SubCellInst2_LFInst_2_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst2_LFInst_2_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_2_LFInst_0_U6  ( .A1(
        PermutationOutput2[11]), .A2(\Red_SubCellInst2_LFInst_2_LFInst_0_n11 ), 
        .ZN(\Red_SubCellInst2_LFInst_2_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst2_LFInst_2_LFInst_0_U5  ( .A(PermutationOutput2[9]), 
        .ZN(\Red_SubCellInst2_LFInst_2_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_2_LFInst_0_U4  ( .A1(
        PermutationOutput2[10]), .A2(\Red_SubCellInst2_LFInst_2_LFInst_0_n8 ), 
        .ZN(\Red_SubCellInst2_LFInst_2_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst2_LFInst_2_LFInst_0_U3  ( .A(PermutationOutput2[8]), 
        .ZN(\Red_SubCellInst2_LFInst_2_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_2_LFInst_1_U8  ( .A1(
        \Red_SubCellInst2_LFInst_2_LFInst_1_n15 ), .A2(
        \Red_SubCellInst2_LFInst_2_LFInst_1_n14 ), .ZN(Red_MCOutput3[9]) );
  NAND2_X1 \Red_SubCellInst2_LFInst_2_LFInst_1_U7  ( .A1(
        \Red_SubCellInst2_LFInst_2_LFInst_1_n13 ), .A2(PermutationOutput2[9]), 
        .ZN(\Red_SubCellInst2_LFInst_2_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_2_LFInst_1_U6  ( .A1(
        \Red_SubCellInst2_LFInst_2_LFInst_1_n12 ), .A2(PermutationOutput2[8]), 
        .ZN(\Red_SubCellInst2_LFInst_2_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_2_LFInst_1_U5  ( .A1(
        PermutationOutput2[11]), .A2(PermutationOutput2[10]), .ZN(
        \Red_SubCellInst2_LFInst_2_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst2_LFInst_2_LFInst_1_U4  ( .A1(PermutationOutput2[10]), 
        .A2(\Red_SubCellInst2_LFInst_2_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst2_LFInst_2_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_2_LFInst_1_U3  ( .A(PermutationOutput2[8]), 
        .B(PermutationOutput2[11]), .ZN(
        \Red_SubCellInst2_LFInst_2_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_2_LFInst_2_U10  ( .A1(
        \Red_SubCellInst2_LFInst_2_LFInst_2_n19 ), .A2(
        \Red_SubCellInst2_LFInst_2_LFInst_2_n18 ), .ZN(Red_MCOutput3[10]) );
  AND2_X1 \Red_SubCellInst2_LFInst_2_LFInst_2_U9  ( .A1(
        \Red_SubCellInst2_LFInst_2_LFInst_2_n17 ), .A2(PermutationOutput2[8]), 
        .ZN(\Red_SubCellInst2_LFInst_2_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_2_LFInst_2_U8  ( .A1(PermutationOutput2[10]), .A2(PermutationOutput2[9]), .ZN(\Red_SubCellInst2_LFInst_2_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_2_LFInst_2_U7  ( .A(
        \Red_SubCellInst2_LFInst_2_LFInst_2_n16 ), .B(
        \Red_SubCellInst2_LFInst_2_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst2_LFInst_2_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_2_LFInst_2_U6  ( .A1(PermutationOutput2[11]), .A2(\Red_SubCellInst2_LFInst_2_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst2_LFInst_2_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst2_LFInst_2_LFInst_2_U5  ( .A(PermutationOutput2[9]), 
        .ZN(\Red_SubCellInst2_LFInst_2_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_2_LFInst_2_U4  ( .A1(
        PermutationOutput2[10]), .A2(\Red_SubCellInst2_LFInst_2_LFInst_2_n13 ), 
        .ZN(\Red_SubCellInst2_LFInst_2_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst2_LFInst_2_LFInst_2_U3  ( .A(PermutationOutput2[8]), 
        .ZN(\Red_SubCellInst2_LFInst_2_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_2_LFInst_3_U6  ( .A(PermutationOutput2[9]), 
        .B(\Red_SubCellInst2_LFInst_2_LFInst_3_n8 ), .ZN(Red_MCOutput3[11]) );
  NOR2_X1 \Red_SubCellInst2_LFInst_2_LFInst_3_U5  ( .A1(
        \Red_SubCellInst2_LFInst_2_LFInst_3_n7 ), .A2(
        \Red_SubCellInst2_LFInst_2_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst2_LFInst_2_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_2_LFInst_3_U4  ( .A1(PermutationOutput2[10]), .A2(PermutationOutput2[11]), .ZN(\Red_SubCellInst2_LFInst_2_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst2_LFInst_2_LFInst_3_U3  ( .A1(PermutationOutput2[11]), .A2(PermutationOutput2[8]), .ZN(\Red_SubCellInst2_LFInst_2_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_3_LFInst_0_U10  ( .A1(
        \Red_SubCellInst2_LFInst_3_LFInst_0_n14 ), .A2(
        \Red_SubCellInst2_LFInst_3_LFInst_0_n13 ), .ZN(Red_MCOutput3[12]) );
  NAND2_X1 \Red_SubCellInst2_LFInst_3_LFInst_0_U9  ( .A1(
        PermutationOutput2[12]), .A2(\Red_SubCellInst2_LFInst_3_LFInst_0_n12 ), 
        .ZN(\Red_SubCellInst2_LFInst_3_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_3_LFInst_0_U8  ( .A1(
        \Red_SubCellInst2_LFInst_3_LFInst_0_n11 ), .A2(PermutationOutput2[14]), 
        .ZN(\Red_SubCellInst2_LFInst_3_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_3_LFInst_0_U7  ( .A(
        \Red_SubCellInst2_LFInst_3_LFInst_0_n10 ), .B(
        \Red_SubCellInst2_LFInst_3_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst2_LFInst_3_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_3_LFInst_0_U6  ( .A1(
        PermutationOutput2[15]), .A2(\Red_SubCellInst2_LFInst_3_LFInst_0_n11 ), 
        .ZN(\Red_SubCellInst2_LFInst_3_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst2_LFInst_3_LFInst_0_U5  ( .A(PermutationOutput2[13]), 
        .ZN(\Red_SubCellInst2_LFInst_3_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_3_LFInst_0_U4  ( .A1(
        PermutationOutput2[14]), .A2(\Red_SubCellInst2_LFInst_3_LFInst_0_n8 ), 
        .ZN(\Red_SubCellInst2_LFInst_3_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst2_LFInst_3_LFInst_0_U3  ( .A(PermutationOutput2[12]), 
        .ZN(\Red_SubCellInst2_LFInst_3_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_3_LFInst_1_U8  ( .A1(
        \Red_SubCellInst2_LFInst_3_LFInst_1_n15 ), .A2(
        \Red_SubCellInst2_LFInst_3_LFInst_1_n14 ), .ZN(Red_MCOutput3[13]) );
  NAND2_X1 \Red_SubCellInst2_LFInst_3_LFInst_1_U7  ( .A1(
        \Red_SubCellInst2_LFInst_3_LFInst_1_n13 ), .A2(PermutationOutput2[13]), 
        .ZN(\Red_SubCellInst2_LFInst_3_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_3_LFInst_1_U6  ( .A1(
        \Red_SubCellInst2_LFInst_3_LFInst_1_n12 ), .A2(PermutationOutput2[12]), 
        .ZN(\Red_SubCellInst2_LFInst_3_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_3_LFInst_1_U5  ( .A1(
        PermutationOutput2[15]), .A2(PermutationOutput2[14]), .ZN(
        \Red_SubCellInst2_LFInst_3_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst2_LFInst_3_LFInst_1_U4  ( .A1(PermutationOutput2[14]), 
        .A2(\Red_SubCellInst2_LFInst_3_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst2_LFInst_3_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_3_LFInst_1_U3  ( .A(PermutationOutput2[12]), .B(PermutationOutput2[15]), .ZN(\Red_SubCellInst2_LFInst_3_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_3_LFInst_2_U10  ( .A1(
        \Red_SubCellInst2_LFInst_3_LFInst_2_n19 ), .A2(
        \Red_SubCellInst2_LFInst_3_LFInst_2_n18 ), .ZN(Red_MCOutput3[14]) );
  AND2_X1 \Red_SubCellInst2_LFInst_3_LFInst_2_U9  ( .A1(
        \Red_SubCellInst2_LFInst_3_LFInst_2_n17 ), .A2(PermutationOutput2[12]), 
        .ZN(\Red_SubCellInst2_LFInst_3_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_3_LFInst_2_U8  ( .A1(PermutationOutput2[14]), .A2(PermutationOutput2[13]), .ZN(\Red_SubCellInst2_LFInst_3_LFInst_2_n17 )
         );
  XNOR2_X1 \Red_SubCellInst2_LFInst_3_LFInst_2_U7  ( .A(
        \Red_SubCellInst2_LFInst_3_LFInst_2_n16 ), .B(
        \Red_SubCellInst2_LFInst_3_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst2_LFInst_3_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_3_LFInst_2_U6  ( .A1(PermutationOutput2[15]), .A2(\Red_SubCellInst2_LFInst_3_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst2_LFInst_3_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst2_LFInst_3_LFInst_2_U5  ( .A(PermutationOutput2[13]), 
        .ZN(\Red_SubCellInst2_LFInst_3_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_3_LFInst_2_U4  ( .A1(
        PermutationOutput2[14]), .A2(\Red_SubCellInst2_LFInst_3_LFInst_2_n13 ), 
        .ZN(\Red_SubCellInst2_LFInst_3_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst2_LFInst_3_LFInst_2_U3  ( .A(PermutationOutput2[12]), 
        .ZN(\Red_SubCellInst2_LFInst_3_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_3_LFInst_3_U6  ( .A(PermutationOutput2[13]), .B(\Red_SubCellInst2_LFInst_3_LFInst_3_n8 ), .ZN(Red_MCOutput3[15]) );
  NOR2_X1 \Red_SubCellInst2_LFInst_3_LFInst_3_U5  ( .A1(
        \Red_SubCellInst2_LFInst_3_LFInst_3_n7 ), .A2(
        \Red_SubCellInst2_LFInst_3_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst2_LFInst_3_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_3_LFInst_3_U4  ( .A1(PermutationOutput2[14]), .A2(PermutationOutput2[15]), .ZN(\Red_SubCellInst2_LFInst_3_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst2_LFInst_3_LFInst_3_U3  ( .A1(PermutationOutput2[15]), .A2(PermutationOutput2[12]), .ZN(\Red_SubCellInst2_LFInst_3_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_4_LFInst_0_U10  ( .A1(
        \Red_SubCellInst2_LFInst_4_LFInst_0_n14 ), .A2(
        \Red_SubCellInst2_LFInst_4_LFInst_0_n13 ), .ZN(Red_MCOutput3[16]) );
  NAND2_X1 \Red_SubCellInst2_LFInst_4_LFInst_0_U9  ( .A1(
        PermutationOutput2[16]), .A2(\Red_SubCellInst2_LFInst_4_LFInst_0_n12 ), 
        .ZN(\Red_SubCellInst2_LFInst_4_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_4_LFInst_0_U8  ( .A1(
        \Red_SubCellInst2_LFInst_4_LFInst_0_n11 ), .A2(PermutationOutput2[18]), 
        .ZN(\Red_SubCellInst2_LFInst_4_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_4_LFInst_0_U7  ( .A(
        \Red_SubCellInst2_LFInst_4_LFInst_0_n10 ), .B(
        \Red_SubCellInst2_LFInst_4_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst2_LFInst_4_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_4_LFInst_0_U6  ( .A1(
        PermutationOutput2[19]), .A2(\Red_SubCellInst2_LFInst_4_LFInst_0_n11 ), 
        .ZN(\Red_SubCellInst2_LFInst_4_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst2_LFInst_4_LFInst_0_U5  ( .A(PermutationOutput2[17]), 
        .ZN(\Red_SubCellInst2_LFInst_4_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_4_LFInst_0_U4  ( .A1(
        PermutationOutput2[18]), .A2(\Red_SubCellInst2_LFInst_4_LFInst_0_n8 ), 
        .ZN(\Red_SubCellInst2_LFInst_4_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst2_LFInst_4_LFInst_0_U3  ( .A(PermutationOutput2[16]), 
        .ZN(\Red_SubCellInst2_LFInst_4_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_4_LFInst_1_U8  ( .A1(
        \Red_SubCellInst2_LFInst_4_LFInst_1_n15 ), .A2(
        \Red_SubCellInst2_LFInst_4_LFInst_1_n14 ), .ZN(Red_MCOutput3[17]) );
  NAND2_X1 \Red_SubCellInst2_LFInst_4_LFInst_1_U7  ( .A1(
        \Red_SubCellInst2_LFInst_4_LFInst_1_n13 ), .A2(PermutationOutput2[17]), 
        .ZN(\Red_SubCellInst2_LFInst_4_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_4_LFInst_1_U6  ( .A1(
        \Red_SubCellInst2_LFInst_4_LFInst_1_n12 ), .A2(PermutationOutput2[16]), 
        .ZN(\Red_SubCellInst2_LFInst_4_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_4_LFInst_1_U5  ( .A1(
        PermutationOutput2[19]), .A2(PermutationOutput2[18]), .ZN(
        \Red_SubCellInst2_LFInst_4_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst2_LFInst_4_LFInst_1_U4  ( .A1(PermutationOutput2[18]), 
        .A2(\Red_SubCellInst2_LFInst_4_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst2_LFInst_4_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_4_LFInst_1_U3  ( .A(PermutationOutput2[16]), .B(PermutationOutput2[19]), .ZN(\Red_SubCellInst2_LFInst_4_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_4_LFInst_2_U10  ( .A1(
        \Red_SubCellInst2_LFInst_4_LFInst_2_n19 ), .A2(
        \Red_SubCellInst2_LFInst_4_LFInst_2_n18 ), .ZN(Red_MCOutput3[18]) );
  AND2_X1 \Red_SubCellInst2_LFInst_4_LFInst_2_U9  ( .A1(
        \Red_SubCellInst2_LFInst_4_LFInst_2_n17 ), .A2(PermutationOutput2[16]), 
        .ZN(\Red_SubCellInst2_LFInst_4_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_4_LFInst_2_U8  ( .A1(PermutationOutput2[18]), .A2(PermutationOutput2[17]), .ZN(\Red_SubCellInst2_LFInst_4_LFInst_2_n17 )
         );
  XNOR2_X1 \Red_SubCellInst2_LFInst_4_LFInst_2_U7  ( .A(
        \Red_SubCellInst2_LFInst_4_LFInst_2_n16 ), .B(
        \Red_SubCellInst2_LFInst_4_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst2_LFInst_4_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_4_LFInst_2_U6  ( .A1(PermutationOutput2[19]), .A2(\Red_SubCellInst2_LFInst_4_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst2_LFInst_4_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst2_LFInst_4_LFInst_2_U5  ( .A(PermutationOutput2[17]), 
        .ZN(\Red_SubCellInst2_LFInst_4_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_4_LFInst_2_U4  ( .A1(
        PermutationOutput2[18]), .A2(\Red_SubCellInst2_LFInst_4_LFInst_2_n13 ), 
        .ZN(\Red_SubCellInst2_LFInst_4_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst2_LFInst_4_LFInst_2_U3  ( .A(PermutationOutput2[16]), 
        .ZN(\Red_SubCellInst2_LFInst_4_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_4_LFInst_3_U6  ( .A(PermutationOutput2[17]), .B(\Red_SubCellInst2_LFInst_4_LFInst_3_n8 ), .ZN(Red_MCOutput3[19]) );
  NOR2_X1 \Red_SubCellInst2_LFInst_4_LFInst_3_U5  ( .A1(
        \Red_SubCellInst2_LFInst_4_LFInst_3_n7 ), .A2(
        \Red_SubCellInst2_LFInst_4_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst2_LFInst_4_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_4_LFInst_3_U4  ( .A1(PermutationOutput2[18]), .A2(PermutationOutput2[19]), .ZN(\Red_SubCellInst2_LFInst_4_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst2_LFInst_4_LFInst_3_U3  ( .A1(PermutationOutput2[19]), .A2(PermutationOutput2[16]), .ZN(\Red_SubCellInst2_LFInst_4_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_5_LFInst_0_U10  ( .A1(
        \Red_SubCellInst2_LFInst_5_LFInst_0_n14 ), .A2(
        \Red_SubCellInst2_LFInst_5_LFInst_0_n13 ), .ZN(Red_MCOutput3[20]) );
  NAND2_X1 \Red_SubCellInst2_LFInst_5_LFInst_0_U9  ( .A1(
        PermutationOutput2[20]), .A2(\Red_SubCellInst2_LFInst_5_LFInst_0_n12 ), 
        .ZN(\Red_SubCellInst2_LFInst_5_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_5_LFInst_0_U8  ( .A1(
        \Red_SubCellInst2_LFInst_5_LFInst_0_n11 ), .A2(PermutationOutput2[22]), 
        .ZN(\Red_SubCellInst2_LFInst_5_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_5_LFInst_0_U7  ( .A(
        \Red_SubCellInst2_LFInst_5_LFInst_0_n10 ), .B(
        \Red_SubCellInst2_LFInst_5_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst2_LFInst_5_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_5_LFInst_0_U6  ( .A1(
        PermutationOutput2[23]), .A2(\Red_SubCellInst2_LFInst_5_LFInst_0_n11 ), 
        .ZN(\Red_SubCellInst2_LFInst_5_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst2_LFInst_5_LFInst_0_U5  ( .A(PermutationOutput2[21]), 
        .ZN(\Red_SubCellInst2_LFInst_5_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_5_LFInst_0_U4  ( .A1(
        PermutationOutput2[22]), .A2(\Red_SubCellInst2_LFInst_5_LFInst_0_n8 ), 
        .ZN(\Red_SubCellInst2_LFInst_5_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst2_LFInst_5_LFInst_0_U3  ( .A(PermutationOutput2[20]), 
        .ZN(\Red_SubCellInst2_LFInst_5_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_5_LFInst_1_U8  ( .A1(
        \Red_SubCellInst2_LFInst_5_LFInst_1_n15 ), .A2(
        \Red_SubCellInst2_LFInst_5_LFInst_1_n14 ), .ZN(Red_MCOutput3[21]) );
  NAND2_X1 \Red_SubCellInst2_LFInst_5_LFInst_1_U7  ( .A1(
        \Red_SubCellInst2_LFInst_5_LFInst_1_n13 ), .A2(PermutationOutput2[21]), 
        .ZN(\Red_SubCellInst2_LFInst_5_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_5_LFInst_1_U6  ( .A1(
        \Red_SubCellInst2_LFInst_5_LFInst_1_n12 ), .A2(PermutationOutput2[20]), 
        .ZN(\Red_SubCellInst2_LFInst_5_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_5_LFInst_1_U5  ( .A1(
        PermutationOutput2[23]), .A2(PermutationOutput2[22]), .ZN(
        \Red_SubCellInst2_LFInst_5_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst2_LFInst_5_LFInst_1_U4  ( .A1(PermutationOutput2[22]), 
        .A2(\Red_SubCellInst2_LFInst_5_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst2_LFInst_5_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_5_LFInst_1_U3  ( .A(PermutationOutput2[20]), .B(PermutationOutput2[23]), .ZN(\Red_SubCellInst2_LFInst_5_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_5_LFInst_2_U10  ( .A1(
        \Red_SubCellInst2_LFInst_5_LFInst_2_n19 ), .A2(
        \Red_SubCellInst2_LFInst_5_LFInst_2_n18 ), .ZN(Red_MCOutput3[22]) );
  AND2_X1 \Red_SubCellInst2_LFInst_5_LFInst_2_U9  ( .A1(
        \Red_SubCellInst2_LFInst_5_LFInst_2_n17 ), .A2(PermutationOutput2[20]), 
        .ZN(\Red_SubCellInst2_LFInst_5_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_5_LFInst_2_U8  ( .A1(PermutationOutput2[22]), .A2(PermutationOutput2[21]), .ZN(\Red_SubCellInst2_LFInst_5_LFInst_2_n17 )
         );
  XNOR2_X1 \Red_SubCellInst2_LFInst_5_LFInst_2_U7  ( .A(
        \Red_SubCellInst2_LFInst_5_LFInst_2_n16 ), .B(
        \Red_SubCellInst2_LFInst_5_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst2_LFInst_5_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_5_LFInst_2_U6  ( .A1(PermutationOutput2[23]), .A2(\Red_SubCellInst2_LFInst_5_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst2_LFInst_5_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst2_LFInst_5_LFInst_2_U5  ( .A(PermutationOutput2[21]), 
        .ZN(\Red_SubCellInst2_LFInst_5_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_5_LFInst_2_U4  ( .A1(
        PermutationOutput2[22]), .A2(\Red_SubCellInst2_LFInst_5_LFInst_2_n13 ), 
        .ZN(\Red_SubCellInst2_LFInst_5_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst2_LFInst_5_LFInst_2_U3  ( .A(PermutationOutput2[20]), 
        .ZN(\Red_SubCellInst2_LFInst_5_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_5_LFInst_3_U6  ( .A(PermutationOutput2[21]), .B(\Red_SubCellInst2_LFInst_5_LFInst_3_n8 ), .ZN(Red_MCOutput3[23]) );
  NOR2_X1 \Red_SubCellInst2_LFInst_5_LFInst_3_U5  ( .A1(
        \Red_SubCellInst2_LFInst_5_LFInst_3_n7 ), .A2(
        \Red_SubCellInst2_LFInst_5_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst2_LFInst_5_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_5_LFInst_3_U4  ( .A1(PermutationOutput2[22]), .A2(PermutationOutput2[23]), .ZN(\Red_SubCellInst2_LFInst_5_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst2_LFInst_5_LFInst_3_U3  ( .A1(PermutationOutput2[23]), .A2(PermutationOutput2[20]), .ZN(\Red_SubCellInst2_LFInst_5_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_6_LFInst_0_U10  ( .A1(
        \Red_SubCellInst2_LFInst_6_LFInst_0_n14 ), .A2(
        \Red_SubCellInst2_LFInst_6_LFInst_0_n13 ), .ZN(Red_MCOutput3[24]) );
  NAND2_X1 \Red_SubCellInst2_LFInst_6_LFInst_0_U9  ( .A1(
        PermutationOutput2[24]), .A2(\Red_SubCellInst2_LFInst_6_LFInst_0_n12 ), 
        .ZN(\Red_SubCellInst2_LFInst_6_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_6_LFInst_0_U8  ( .A1(
        \Red_SubCellInst2_LFInst_6_LFInst_0_n11 ), .A2(PermutationOutput2[26]), 
        .ZN(\Red_SubCellInst2_LFInst_6_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_6_LFInst_0_U7  ( .A(
        \Red_SubCellInst2_LFInst_6_LFInst_0_n10 ), .B(
        \Red_SubCellInst2_LFInst_6_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst2_LFInst_6_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_6_LFInst_0_U6  ( .A1(
        PermutationOutput2[27]), .A2(\Red_SubCellInst2_LFInst_6_LFInst_0_n11 ), 
        .ZN(\Red_SubCellInst2_LFInst_6_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst2_LFInst_6_LFInst_0_U5  ( .A(PermutationOutput2[25]), 
        .ZN(\Red_SubCellInst2_LFInst_6_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_6_LFInst_0_U4  ( .A1(
        PermutationOutput2[26]), .A2(\Red_SubCellInst2_LFInst_6_LFInst_0_n8 ), 
        .ZN(\Red_SubCellInst2_LFInst_6_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst2_LFInst_6_LFInst_0_U3  ( .A(PermutationOutput2[24]), 
        .ZN(\Red_SubCellInst2_LFInst_6_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_6_LFInst_1_U8  ( .A1(
        \Red_SubCellInst2_LFInst_6_LFInst_1_n15 ), .A2(
        \Red_SubCellInst2_LFInst_6_LFInst_1_n14 ), .ZN(Red_MCOutput3[25]) );
  NAND2_X1 \Red_SubCellInst2_LFInst_6_LFInst_1_U7  ( .A1(
        \Red_SubCellInst2_LFInst_6_LFInst_1_n13 ), .A2(PermutationOutput2[25]), 
        .ZN(\Red_SubCellInst2_LFInst_6_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_6_LFInst_1_U6  ( .A1(
        \Red_SubCellInst2_LFInst_6_LFInst_1_n12 ), .A2(PermutationOutput2[24]), 
        .ZN(\Red_SubCellInst2_LFInst_6_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_6_LFInst_1_U5  ( .A1(
        PermutationOutput2[27]), .A2(PermutationOutput2[26]), .ZN(
        \Red_SubCellInst2_LFInst_6_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst2_LFInst_6_LFInst_1_U4  ( .A1(PermutationOutput2[26]), 
        .A2(\Red_SubCellInst2_LFInst_6_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst2_LFInst_6_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_6_LFInst_1_U3  ( .A(PermutationOutput2[24]), .B(PermutationOutput2[27]), .ZN(\Red_SubCellInst2_LFInst_6_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_6_LFInst_2_U10  ( .A1(
        \Red_SubCellInst2_LFInst_6_LFInst_2_n19 ), .A2(
        \Red_SubCellInst2_LFInst_6_LFInst_2_n18 ), .ZN(Red_MCOutput3[26]) );
  AND2_X1 \Red_SubCellInst2_LFInst_6_LFInst_2_U9  ( .A1(
        \Red_SubCellInst2_LFInst_6_LFInst_2_n17 ), .A2(PermutationOutput2[24]), 
        .ZN(\Red_SubCellInst2_LFInst_6_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_6_LFInst_2_U8  ( .A1(PermutationOutput2[26]), .A2(PermutationOutput2[25]), .ZN(\Red_SubCellInst2_LFInst_6_LFInst_2_n17 )
         );
  XNOR2_X1 \Red_SubCellInst2_LFInst_6_LFInst_2_U7  ( .A(
        \Red_SubCellInst2_LFInst_6_LFInst_2_n16 ), .B(
        \Red_SubCellInst2_LFInst_6_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst2_LFInst_6_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_6_LFInst_2_U6  ( .A1(PermutationOutput2[27]), .A2(\Red_SubCellInst2_LFInst_6_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst2_LFInst_6_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst2_LFInst_6_LFInst_2_U5  ( .A(PermutationOutput2[25]), 
        .ZN(\Red_SubCellInst2_LFInst_6_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_6_LFInst_2_U4  ( .A1(
        PermutationOutput2[26]), .A2(\Red_SubCellInst2_LFInst_6_LFInst_2_n13 ), 
        .ZN(\Red_SubCellInst2_LFInst_6_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst2_LFInst_6_LFInst_2_U3  ( .A(PermutationOutput2[24]), 
        .ZN(\Red_SubCellInst2_LFInst_6_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_6_LFInst_3_U6  ( .A(PermutationOutput2[25]), .B(\Red_SubCellInst2_LFInst_6_LFInst_3_n8 ), .ZN(Red_MCOutput3[27]) );
  NOR2_X1 \Red_SubCellInst2_LFInst_6_LFInst_3_U5  ( .A1(
        \Red_SubCellInst2_LFInst_6_LFInst_3_n7 ), .A2(
        \Red_SubCellInst2_LFInst_6_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst2_LFInst_6_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_6_LFInst_3_U4  ( .A1(PermutationOutput2[26]), .A2(PermutationOutput2[27]), .ZN(\Red_SubCellInst2_LFInst_6_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst2_LFInst_6_LFInst_3_U3  ( .A1(PermutationOutput2[27]), .A2(PermutationOutput2[24]), .ZN(\Red_SubCellInst2_LFInst_6_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_7_LFInst_0_U10  ( .A1(
        \Red_SubCellInst2_LFInst_7_LFInst_0_n14 ), .A2(
        \Red_SubCellInst2_LFInst_7_LFInst_0_n13 ), .ZN(Red_MCOutput3[28]) );
  NAND2_X1 \Red_SubCellInst2_LFInst_7_LFInst_0_U9  ( .A1(
        PermutationOutput2[28]), .A2(\Red_SubCellInst2_LFInst_7_LFInst_0_n12 ), 
        .ZN(\Red_SubCellInst2_LFInst_7_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_7_LFInst_0_U8  ( .A1(
        \Red_SubCellInst2_LFInst_7_LFInst_0_n11 ), .A2(PermutationOutput2[30]), 
        .ZN(\Red_SubCellInst2_LFInst_7_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_7_LFInst_0_U7  ( .A(
        \Red_SubCellInst2_LFInst_7_LFInst_0_n10 ), .B(
        \Red_SubCellInst2_LFInst_7_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst2_LFInst_7_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_7_LFInst_0_U6  ( .A1(
        PermutationOutput2[31]), .A2(\Red_SubCellInst2_LFInst_7_LFInst_0_n11 ), 
        .ZN(\Red_SubCellInst2_LFInst_7_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst2_LFInst_7_LFInst_0_U5  ( .A(PermutationOutput2[29]), 
        .ZN(\Red_SubCellInst2_LFInst_7_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_7_LFInst_0_U4  ( .A1(
        PermutationOutput2[30]), .A2(\Red_SubCellInst2_LFInst_7_LFInst_0_n8 ), 
        .ZN(\Red_SubCellInst2_LFInst_7_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst2_LFInst_7_LFInst_0_U3  ( .A(PermutationOutput2[28]), 
        .ZN(\Red_SubCellInst2_LFInst_7_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_7_LFInst_1_U8  ( .A1(
        \Red_SubCellInst2_LFInst_7_LFInst_1_n15 ), .A2(
        \Red_SubCellInst2_LFInst_7_LFInst_1_n14 ), .ZN(Red_MCOutput3[29]) );
  NAND2_X1 \Red_SubCellInst2_LFInst_7_LFInst_1_U7  ( .A1(
        \Red_SubCellInst2_LFInst_7_LFInst_1_n13 ), .A2(PermutationOutput2[29]), 
        .ZN(\Red_SubCellInst2_LFInst_7_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_7_LFInst_1_U6  ( .A1(
        \Red_SubCellInst2_LFInst_7_LFInst_1_n12 ), .A2(PermutationOutput2[28]), 
        .ZN(\Red_SubCellInst2_LFInst_7_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_7_LFInst_1_U5  ( .A1(
        PermutationOutput2[31]), .A2(PermutationOutput2[30]), .ZN(
        \Red_SubCellInst2_LFInst_7_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst2_LFInst_7_LFInst_1_U4  ( .A1(PermutationOutput2[30]), 
        .A2(\Red_SubCellInst2_LFInst_7_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst2_LFInst_7_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_7_LFInst_1_U3  ( .A(PermutationOutput2[28]), .B(PermutationOutput2[31]), .ZN(\Red_SubCellInst2_LFInst_7_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_7_LFInst_2_U10  ( .A1(
        \Red_SubCellInst2_LFInst_7_LFInst_2_n19 ), .A2(
        \Red_SubCellInst2_LFInst_7_LFInst_2_n18 ), .ZN(Red_MCOutput3[30]) );
  AND2_X1 \Red_SubCellInst2_LFInst_7_LFInst_2_U9  ( .A1(
        \Red_SubCellInst2_LFInst_7_LFInst_2_n17 ), .A2(PermutationOutput2[28]), 
        .ZN(\Red_SubCellInst2_LFInst_7_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_7_LFInst_2_U8  ( .A1(PermutationOutput2[30]), .A2(PermutationOutput2[29]), .ZN(\Red_SubCellInst2_LFInst_7_LFInst_2_n17 )
         );
  XNOR2_X1 \Red_SubCellInst2_LFInst_7_LFInst_2_U7  ( .A(
        \Red_SubCellInst2_LFInst_7_LFInst_2_n16 ), .B(
        \Red_SubCellInst2_LFInst_7_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst2_LFInst_7_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_7_LFInst_2_U6  ( .A1(PermutationOutput2[31]), .A2(\Red_SubCellInst2_LFInst_7_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst2_LFInst_7_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst2_LFInst_7_LFInst_2_U5  ( .A(PermutationOutput2[29]), 
        .ZN(\Red_SubCellInst2_LFInst_7_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_7_LFInst_2_U4  ( .A1(
        PermutationOutput2[30]), .A2(\Red_SubCellInst2_LFInst_7_LFInst_2_n13 ), 
        .ZN(\Red_SubCellInst2_LFInst_7_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst2_LFInst_7_LFInst_2_U3  ( .A(PermutationOutput2[28]), 
        .ZN(\Red_SubCellInst2_LFInst_7_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_7_LFInst_3_U6  ( .A(PermutationOutput2[29]), .B(\Red_SubCellInst2_LFInst_7_LFInst_3_n8 ), .ZN(Red_MCOutput3[31]) );
  NOR2_X1 \Red_SubCellInst2_LFInst_7_LFInst_3_U5  ( .A1(
        \Red_SubCellInst2_LFInst_7_LFInst_3_n7 ), .A2(
        \Red_SubCellInst2_LFInst_7_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst2_LFInst_7_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_7_LFInst_3_U4  ( .A1(PermutationOutput2[30]), .A2(PermutationOutput2[31]), .ZN(\Red_SubCellInst2_LFInst_7_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst2_LFInst_7_LFInst_3_U3  ( .A1(PermutationOutput2[31]), .A2(PermutationOutput2[28]), .ZN(\Red_SubCellInst2_LFInst_7_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_8_LFInst_0_U10  ( .A1(
        \Red_SubCellInst2_LFInst_8_LFInst_0_n14 ), .A2(
        \Red_SubCellInst2_LFInst_8_LFInst_0_n13 ), .ZN(Red_Feedback2[32]) );
  NAND2_X1 \Red_SubCellInst2_LFInst_8_LFInst_0_U9  ( .A1(
        PermutationOutput2[32]), .A2(\Red_SubCellInst2_LFInst_8_LFInst_0_n12 ), 
        .ZN(\Red_SubCellInst2_LFInst_8_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_8_LFInst_0_U8  ( .A1(
        \Red_SubCellInst2_LFInst_8_LFInst_0_n11 ), .A2(PermutationOutput2[34]), 
        .ZN(\Red_SubCellInst2_LFInst_8_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_8_LFInst_0_U7  ( .A(
        \Red_SubCellInst2_LFInst_8_LFInst_0_n10 ), .B(
        \Red_SubCellInst2_LFInst_8_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst2_LFInst_8_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_8_LFInst_0_U6  ( .A1(
        PermutationOutput2[35]), .A2(\Red_SubCellInst2_LFInst_8_LFInst_0_n11 ), 
        .ZN(\Red_SubCellInst2_LFInst_8_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst2_LFInst_8_LFInst_0_U5  ( .A(PermutationOutput2[33]), 
        .ZN(\Red_SubCellInst2_LFInst_8_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_8_LFInst_0_U4  ( .A1(
        PermutationOutput2[34]), .A2(\Red_SubCellInst2_LFInst_8_LFInst_0_n8 ), 
        .ZN(\Red_SubCellInst2_LFInst_8_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst2_LFInst_8_LFInst_0_U3  ( .A(PermutationOutput2[32]), 
        .ZN(\Red_SubCellInst2_LFInst_8_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_8_LFInst_1_U8  ( .A1(
        \Red_SubCellInst2_LFInst_8_LFInst_1_n15 ), .A2(
        \Red_SubCellInst2_LFInst_8_LFInst_1_n14 ), .ZN(Red_Feedback2[33]) );
  NAND2_X1 \Red_SubCellInst2_LFInst_8_LFInst_1_U7  ( .A1(
        \Red_SubCellInst2_LFInst_8_LFInst_1_n13 ), .A2(PermutationOutput2[33]), 
        .ZN(\Red_SubCellInst2_LFInst_8_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_8_LFInst_1_U6  ( .A1(
        \Red_SubCellInst2_LFInst_8_LFInst_1_n12 ), .A2(PermutationOutput2[32]), 
        .ZN(\Red_SubCellInst2_LFInst_8_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_8_LFInst_1_U5  ( .A1(
        PermutationOutput2[35]), .A2(PermutationOutput2[34]), .ZN(
        \Red_SubCellInst2_LFInst_8_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst2_LFInst_8_LFInst_1_U4  ( .A1(PermutationOutput2[34]), 
        .A2(\Red_SubCellInst2_LFInst_8_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst2_LFInst_8_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_8_LFInst_1_U3  ( .A(PermutationOutput2[32]), .B(PermutationOutput2[35]), .ZN(\Red_SubCellInst2_LFInst_8_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_8_LFInst_2_U10  ( .A1(
        \Red_SubCellInst2_LFInst_8_LFInst_2_n19 ), .A2(
        \Red_SubCellInst2_LFInst_8_LFInst_2_n18 ), .ZN(Red_Feedback2[34]) );
  AND2_X1 \Red_SubCellInst2_LFInst_8_LFInst_2_U9  ( .A1(
        \Red_SubCellInst2_LFInst_8_LFInst_2_n17 ), .A2(PermutationOutput2[32]), 
        .ZN(\Red_SubCellInst2_LFInst_8_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_8_LFInst_2_U8  ( .A1(PermutationOutput2[34]), .A2(PermutationOutput2[33]), .ZN(\Red_SubCellInst2_LFInst_8_LFInst_2_n17 )
         );
  XNOR2_X1 \Red_SubCellInst2_LFInst_8_LFInst_2_U7  ( .A(
        \Red_SubCellInst2_LFInst_8_LFInst_2_n16 ), .B(
        \Red_SubCellInst2_LFInst_8_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst2_LFInst_8_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_8_LFInst_2_U6  ( .A1(PermutationOutput2[35]), .A2(\Red_SubCellInst2_LFInst_8_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst2_LFInst_8_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst2_LFInst_8_LFInst_2_U5  ( .A(PermutationOutput2[33]), 
        .ZN(\Red_SubCellInst2_LFInst_8_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_8_LFInst_2_U4  ( .A1(
        PermutationOutput2[34]), .A2(\Red_SubCellInst2_LFInst_8_LFInst_2_n13 ), 
        .ZN(\Red_SubCellInst2_LFInst_8_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst2_LFInst_8_LFInst_2_U3  ( .A(PermutationOutput2[32]), 
        .ZN(\Red_SubCellInst2_LFInst_8_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_8_LFInst_3_U6  ( .A(PermutationOutput2[33]), .B(\Red_SubCellInst2_LFInst_8_LFInst_3_n8 ), .ZN(Red_Feedback2[35]) );
  NOR2_X1 \Red_SubCellInst2_LFInst_8_LFInst_3_U5  ( .A1(
        \Red_SubCellInst2_LFInst_8_LFInst_3_n7 ), .A2(
        \Red_SubCellInst2_LFInst_8_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst2_LFInst_8_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_8_LFInst_3_U4  ( .A1(PermutationOutput2[34]), .A2(PermutationOutput2[35]), .ZN(\Red_SubCellInst2_LFInst_8_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst2_LFInst_8_LFInst_3_U3  ( .A1(PermutationOutput2[35]), .A2(PermutationOutput2[32]), .ZN(\Red_SubCellInst2_LFInst_8_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_9_LFInst_0_U10  ( .A1(
        \Red_SubCellInst2_LFInst_9_LFInst_0_n14 ), .A2(
        \Red_SubCellInst2_LFInst_9_LFInst_0_n13 ), .ZN(Red_Feedback2[36]) );
  NAND2_X1 \Red_SubCellInst2_LFInst_9_LFInst_0_U9  ( .A1(
        PermutationOutput2[36]), .A2(\Red_SubCellInst2_LFInst_9_LFInst_0_n12 ), 
        .ZN(\Red_SubCellInst2_LFInst_9_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_9_LFInst_0_U8  ( .A1(
        \Red_SubCellInst2_LFInst_9_LFInst_0_n11 ), .A2(PermutationOutput2[38]), 
        .ZN(\Red_SubCellInst2_LFInst_9_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_9_LFInst_0_U7  ( .A(
        \Red_SubCellInst2_LFInst_9_LFInst_0_n10 ), .B(
        \Red_SubCellInst2_LFInst_9_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst2_LFInst_9_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_9_LFInst_0_U6  ( .A1(
        PermutationOutput2[39]), .A2(\Red_SubCellInst2_LFInst_9_LFInst_0_n11 ), 
        .ZN(\Red_SubCellInst2_LFInst_9_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst2_LFInst_9_LFInst_0_U5  ( .A(PermutationOutput2[37]), 
        .ZN(\Red_SubCellInst2_LFInst_9_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_9_LFInst_0_U4  ( .A1(
        PermutationOutput2[38]), .A2(\Red_SubCellInst2_LFInst_9_LFInst_0_n8 ), 
        .ZN(\Red_SubCellInst2_LFInst_9_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst2_LFInst_9_LFInst_0_U3  ( .A(PermutationOutput2[36]), 
        .ZN(\Red_SubCellInst2_LFInst_9_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_9_LFInst_1_U8  ( .A1(
        \Red_SubCellInst2_LFInst_9_LFInst_1_n15 ), .A2(
        \Red_SubCellInst2_LFInst_9_LFInst_1_n14 ), .ZN(Red_Feedback2[37]) );
  NAND2_X1 \Red_SubCellInst2_LFInst_9_LFInst_1_U7  ( .A1(
        \Red_SubCellInst2_LFInst_9_LFInst_1_n13 ), .A2(PermutationOutput2[37]), 
        .ZN(\Red_SubCellInst2_LFInst_9_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_9_LFInst_1_U6  ( .A1(
        \Red_SubCellInst2_LFInst_9_LFInst_1_n12 ), .A2(PermutationOutput2[36]), 
        .ZN(\Red_SubCellInst2_LFInst_9_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_9_LFInst_1_U5  ( .A1(
        PermutationOutput2[39]), .A2(PermutationOutput2[38]), .ZN(
        \Red_SubCellInst2_LFInst_9_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst2_LFInst_9_LFInst_1_U4  ( .A1(PermutationOutput2[38]), 
        .A2(\Red_SubCellInst2_LFInst_9_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst2_LFInst_9_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_9_LFInst_1_U3  ( .A(PermutationOutput2[36]), .B(PermutationOutput2[39]), .ZN(\Red_SubCellInst2_LFInst_9_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_9_LFInst_2_U10  ( .A1(
        \Red_SubCellInst2_LFInst_9_LFInst_2_n19 ), .A2(
        \Red_SubCellInst2_LFInst_9_LFInst_2_n18 ), .ZN(Red_Feedback2[38]) );
  AND2_X1 \Red_SubCellInst2_LFInst_9_LFInst_2_U9  ( .A1(
        \Red_SubCellInst2_LFInst_9_LFInst_2_n17 ), .A2(PermutationOutput2[36]), 
        .ZN(\Red_SubCellInst2_LFInst_9_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_9_LFInst_2_U8  ( .A1(PermutationOutput2[38]), .A2(PermutationOutput2[37]), .ZN(\Red_SubCellInst2_LFInst_9_LFInst_2_n17 )
         );
  XNOR2_X1 \Red_SubCellInst2_LFInst_9_LFInst_2_U7  ( .A(
        \Red_SubCellInst2_LFInst_9_LFInst_2_n16 ), .B(
        \Red_SubCellInst2_LFInst_9_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst2_LFInst_9_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_9_LFInst_2_U6  ( .A1(PermutationOutput2[39]), .A2(\Red_SubCellInst2_LFInst_9_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst2_LFInst_9_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst2_LFInst_9_LFInst_2_U5  ( .A(PermutationOutput2[37]), 
        .ZN(\Red_SubCellInst2_LFInst_9_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_9_LFInst_2_U4  ( .A1(
        PermutationOutput2[38]), .A2(\Red_SubCellInst2_LFInst_9_LFInst_2_n13 ), 
        .ZN(\Red_SubCellInst2_LFInst_9_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst2_LFInst_9_LFInst_2_U3  ( .A(PermutationOutput2[36]), 
        .ZN(\Red_SubCellInst2_LFInst_9_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_9_LFInst_3_U6  ( .A(PermutationOutput2[37]), .B(\Red_SubCellInst2_LFInst_9_LFInst_3_n8 ), .ZN(Red_Feedback2[39]) );
  NOR2_X1 \Red_SubCellInst2_LFInst_9_LFInst_3_U5  ( .A1(
        \Red_SubCellInst2_LFInst_9_LFInst_3_n7 ), .A2(
        \Red_SubCellInst2_LFInst_9_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst2_LFInst_9_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_9_LFInst_3_U4  ( .A1(PermutationOutput2[38]), .A2(PermutationOutput2[39]), .ZN(\Red_SubCellInst2_LFInst_9_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst2_LFInst_9_LFInst_3_U3  ( .A1(PermutationOutput2[39]), .A2(PermutationOutput2[36]), .ZN(\Red_SubCellInst2_LFInst_9_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_10_LFInst_0_U10  ( .A1(
        \Red_SubCellInst2_LFInst_10_LFInst_0_n14 ), .A2(
        \Red_SubCellInst2_LFInst_10_LFInst_0_n13 ), .ZN(Red_Feedback2[40]) );
  NAND2_X1 \Red_SubCellInst2_LFInst_10_LFInst_0_U9  ( .A1(
        PermutationOutput2[40]), .A2(\Red_SubCellInst2_LFInst_10_LFInst_0_n12 ), .ZN(\Red_SubCellInst2_LFInst_10_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_10_LFInst_0_U8  ( .A1(
        \Red_SubCellInst2_LFInst_10_LFInst_0_n11 ), .A2(PermutationOutput2[42]), .ZN(\Red_SubCellInst2_LFInst_10_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_10_LFInst_0_U7  ( .A(
        \Red_SubCellInst2_LFInst_10_LFInst_0_n10 ), .B(
        \Red_SubCellInst2_LFInst_10_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst2_LFInst_10_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_10_LFInst_0_U6  ( .A1(
        PermutationOutput2[43]), .A2(\Red_SubCellInst2_LFInst_10_LFInst_0_n11 ), .ZN(\Red_SubCellInst2_LFInst_10_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst2_LFInst_10_LFInst_0_U5  ( .A(PermutationOutput2[41]), 
        .ZN(\Red_SubCellInst2_LFInst_10_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_10_LFInst_0_U4  ( .A1(
        PermutationOutput2[42]), .A2(\Red_SubCellInst2_LFInst_10_LFInst_0_n8 ), 
        .ZN(\Red_SubCellInst2_LFInst_10_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst2_LFInst_10_LFInst_0_U3  ( .A(PermutationOutput2[40]), 
        .ZN(\Red_SubCellInst2_LFInst_10_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_10_LFInst_1_U8  ( .A1(
        \Red_SubCellInst2_LFInst_10_LFInst_1_n15 ), .A2(
        \Red_SubCellInst2_LFInst_10_LFInst_1_n14 ), .ZN(Red_Feedback2[41]) );
  NAND2_X1 \Red_SubCellInst2_LFInst_10_LFInst_1_U7  ( .A1(
        \Red_SubCellInst2_LFInst_10_LFInst_1_n13 ), .A2(PermutationOutput2[41]), .ZN(\Red_SubCellInst2_LFInst_10_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_10_LFInst_1_U6  ( .A1(
        \Red_SubCellInst2_LFInst_10_LFInst_1_n12 ), .A2(PermutationOutput2[40]), .ZN(\Red_SubCellInst2_LFInst_10_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_10_LFInst_1_U5  ( .A1(
        PermutationOutput2[43]), .A2(PermutationOutput2[42]), .ZN(
        \Red_SubCellInst2_LFInst_10_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst2_LFInst_10_LFInst_1_U4  ( .A1(PermutationOutput2[42]), .A2(\Red_SubCellInst2_LFInst_10_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst2_LFInst_10_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_10_LFInst_1_U3  ( .A(
        PermutationOutput2[40]), .B(PermutationOutput2[43]), .ZN(
        \Red_SubCellInst2_LFInst_10_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_10_LFInst_2_U10  ( .A1(
        \Red_SubCellInst2_LFInst_10_LFInst_2_n19 ), .A2(
        \Red_SubCellInst2_LFInst_10_LFInst_2_n18 ), .ZN(Red_Feedback2[42]) );
  AND2_X1 \Red_SubCellInst2_LFInst_10_LFInst_2_U9  ( .A1(
        \Red_SubCellInst2_LFInst_10_LFInst_2_n17 ), .A2(PermutationOutput2[40]), .ZN(\Red_SubCellInst2_LFInst_10_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_10_LFInst_2_U8  ( .A1(
        PermutationOutput2[42]), .A2(PermutationOutput2[41]), .ZN(
        \Red_SubCellInst2_LFInst_10_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_10_LFInst_2_U7  ( .A(
        \Red_SubCellInst2_LFInst_10_LFInst_2_n16 ), .B(
        \Red_SubCellInst2_LFInst_10_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst2_LFInst_10_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_10_LFInst_2_U6  ( .A1(
        PermutationOutput2[43]), .A2(\Red_SubCellInst2_LFInst_10_LFInst_2_n14 ), .ZN(\Red_SubCellInst2_LFInst_10_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst2_LFInst_10_LFInst_2_U5  ( .A(PermutationOutput2[41]), 
        .ZN(\Red_SubCellInst2_LFInst_10_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_10_LFInst_2_U4  ( .A1(
        PermutationOutput2[42]), .A2(\Red_SubCellInst2_LFInst_10_LFInst_2_n13 ), .ZN(\Red_SubCellInst2_LFInst_10_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst2_LFInst_10_LFInst_2_U3  ( .A(PermutationOutput2[40]), 
        .ZN(\Red_SubCellInst2_LFInst_10_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_10_LFInst_3_U6  ( .A(
        PermutationOutput2[41]), .B(\Red_SubCellInst2_LFInst_10_LFInst_3_n8 ), 
        .ZN(Red_Feedback2[43]) );
  NOR2_X1 \Red_SubCellInst2_LFInst_10_LFInst_3_U5  ( .A1(
        \Red_SubCellInst2_LFInst_10_LFInst_3_n7 ), .A2(
        \Red_SubCellInst2_LFInst_10_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst2_LFInst_10_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_10_LFInst_3_U4  ( .A1(
        PermutationOutput2[42]), .A2(PermutationOutput2[43]), .ZN(
        \Red_SubCellInst2_LFInst_10_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst2_LFInst_10_LFInst_3_U3  ( .A1(
        PermutationOutput2[43]), .A2(PermutationOutput2[40]), .ZN(
        \Red_SubCellInst2_LFInst_10_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_11_LFInst_0_U10  ( .A1(
        \Red_SubCellInst2_LFInst_11_LFInst_0_n14 ), .A2(
        \Red_SubCellInst2_LFInst_11_LFInst_0_n13 ), .ZN(Red_Feedback2[44]) );
  NAND2_X1 \Red_SubCellInst2_LFInst_11_LFInst_0_U9  ( .A1(
        PermutationOutput2[44]), .A2(\Red_SubCellInst2_LFInst_11_LFInst_0_n12 ), .ZN(\Red_SubCellInst2_LFInst_11_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_11_LFInst_0_U8  ( .A1(
        \Red_SubCellInst2_LFInst_11_LFInst_0_n11 ), .A2(PermutationOutput2[46]), .ZN(\Red_SubCellInst2_LFInst_11_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_11_LFInst_0_U7  ( .A(
        \Red_SubCellInst2_LFInst_11_LFInst_0_n10 ), .B(
        \Red_SubCellInst2_LFInst_11_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst2_LFInst_11_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_11_LFInst_0_U6  ( .A1(
        PermutationOutput2[47]), .A2(\Red_SubCellInst2_LFInst_11_LFInst_0_n11 ), .ZN(\Red_SubCellInst2_LFInst_11_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst2_LFInst_11_LFInst_0_U5  ( .A(PermutationOutput2[45]), 
        .ZN(\Red_SubCellInst2_LFInst_11_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_11_LFInst_0_U4  ( .A1(
        PermutationOutput2[46]), .A2(\Red_SubCellInst2_LFInst_11_LFInst_0_n8 ), 
        .ZN(\Red_SubCellInst2_LFInst_11_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst2_LFInst_11_LFInst_0_U3  ( .A(PermutationOutput2[44]), 
        .ZN(\Red_SubCellInst2_LFInst_11_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_11_LFInst_1_U8  ( .A1(
        \Red_SubCellInst2_LFInst_11_LFInst_1_n15 ), .A2(
        \Red_SubCellInst2_LFInst_11_LFInst_1_n14 ), .ZN(Red_Feedback2[45]) );
  NAND2_X1 \Red_SubCellInst2_LFInst_11_LFInst_1_U7  ( .A1(
        \Red_SubCellInst2_LFInst_11_LFInst_1_n13 ), .A2(PermutationOutput2[45]), .ZN(\Red_SubCellInst2_LFInst_11_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_11_LFInst_1_U6  ( .A1(
        \Red_SubCellInst2_LFInst_11_LFInst_1_n12 ), .A2(PermutationOutput2[44]), .ZN(\Red_SubCellInst2_LFInst_11_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_11_LFInst_1_U5  ( .A1(
        PermutationOutput2[47]), .A2(PermutationOutput2[46]), .ZN(
        \Red_SubCellInst2_LFInst_11_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst2_LFInst_11_LFInst_1_U4  ( .A1(PermutationOutput2[46]), .A2(\Red_SubCellInst2_LFInst_11_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst2_LFInst_11_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_11_LFInst_1_U3  ( .A(
        PermutationOutput2[44]), .B(PermutationOutput2[47]), .ZN(
        \Red_SubCellInst2_LFInst_11_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_11_LFInst_2_U10  ( .A1(
        \Red_SubCellInst2_LFInst_11_LFInst_2_n19 ), .A2(
        \Red_SubCellInst2_LFInst_11_LFInst_2_n18 ), .ZN(Red_Feedback2[46]) );
  AND2_X1 \Red_SubCellInst2_LFInst_11_LFInst_2_U9  ( .A1(
        \Red_SubCellInst2_LFInst_11_LFInst_2_n17 ), .A2(PermutationOutput2[44]), .ZN(\Red_SubCellInst2_LFInst_11_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_11_LFInst_2_U8  ( .A1(
        PermutationOutput2[46]), .A2(PermutationOutput2[45]), .ZN(
        \Red_SubCellInst2_LFInst_11_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_11_LFInst_2_U7  ( .A(
        \Red_SubCellInst2_LFInst_11_LFInst_2_n16 ), .B(
        \Red_SubCellInst2_LFInst_11_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst2_LFInst_11_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_11_LFInst_2_U6  ( .A1(
        PermutationOutput2[47]), .A2(\Red_SubCellInst2_LFInst_11_LFInst_2_n14 ), .ZN(\Red_SubCellInst2_LFInst_11_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst2_LFInst_11_LFInst_2_U5  ( .A(PermutationOutput2[45]), 
        .ZN(\Red_SubCellInst2_LFInst_11_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_11_LFInst_2_U4  ( .A1(
        PermutationOutput2[46]), .A2(\Red_SubCellInst2_LFInst_11_LFInst_2_n13 ), .ZN(\Red_SubCellInst2_LFInst_11_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst2_LFInst_11_LFInst_2_U3  ( .A(PermutationOutput2[44]), 
        .ZN(\Red_SubCellInst2_LFInst_11_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_11_LFInst_3_U6  ( .A(
        PermutationOutput2[45]), .B(\Red_SubCellInst2_LFInst_11_LFInst_3_n8 ), 
        .ZN(Red_Feedback2[47]) );
  NOR2_X1 \Red_SubCellInst2_LFInst_11_LFInst_3_U5  ( .A1(
        \Red_SubCellInst2_LFInst_11_LFInst_3_n7 ), .A2(
        \Red_SubCellInst2_LFInst_11_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst2_LFInst_11_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_11_LFInst_3_U4  ( .A1(
        PermutationOutput2[46]), .A2(PermutationOutput2[47]), .ZN(
        \Red_SubCellInst2_LFInst_11_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst2_LFInst_11_LFInst_3_U3  ( .A1(
        PermutationOutput2[47]), .A2(PermutationOutput2[44]), .ZN(
        \Red_SubCellInst2_LFInst_11_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_12_LFInst_0_U10  ( .A1(
        \Red_SubCellInst2_LFInst_12_LFInst_0_n14 ), .A2(
        \Red_SubCellInst2_LFInst_12_LFInst_0_n13 ), .ZN(Red_Feedback2[48]) );
  NAND2_X1 \Red_SubCellInst2_LFInst_12_LFInst_0_U9  ( .A1(
        PermutationOutput2[48]), .A2(\Red_SubCellInst2_LFInst_12_LFInst_0_n12 ), .ZN(\Red_SubCellInst2_LFInst_12_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_12_LFInst_0_U8  ( .A1(
        \Red_SubCellInst2_LFInst_12_LFInst_0_n11 ), .A2(PermutationOutput2[50]), .ZN(\Red_SubCellInst2_LFInst_12_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_12_LFInst_0_U7  ( .A(
        \Red_SubCellInst2_LFInst_12_LFInst_0_n10 ), .B(
        \Red_SubCellInst2_LFInst_12_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst2_LFInst_12_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_12_LFInst_0_U6  ( .A1(
        PermutationOutput2[51]), .A2(\Red_SubCellInst2_LFInst_12_LFInst_0_n11 ), .ZN(\Red_SubCellInst2_LFInst_12_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst2_LFInst_12_LFInst_0_U5  ( .A(PermutationOutput2[49]), 
        .ZN(\Red_SubCellInst2_LFInst_12_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_12_LFInst_0_U4  ( .A1(
        PermutationOutput2[50]), .A2(\Red_SubCellInst2_LFInst_12_LFInst_0_n8 ), 
        .ZN(\Red_SubCellInst2_LFInst_12_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst2_LFInst_12_LFInst_0_U3  ( .A(PermutationOutput2[48]), 
        .ZN(\Red_SubCellInst2_LFInst_12_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_12_LFInst_1_U8  ( .A1(
        \Red_SubCellInst2_LFInst_12_LFInst_1_n15 ), .A2(
        \Red_SubCellInst2_LFInst_12_LFInst_1_n14 ), .ZN(Red_Feedback2[49]) );
  NAND2_X1 \Red_SubCellInst2_LFInst_12_LFInst_1_U7  ( .A1(
        \Red_SubCellInst2_LFInst_12_LFInst_1_n13 ), .A2(PermutationOutput2[49]), .ZN(\Red_SubCellInst2_LFInst_12_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_12_LFInst_1_U6  ( .A1(
        \Red_SubCellInst2_LFInst_12_LFInst_1_n12 ), .A2(PermutationOutput2[48]), .ZN(\Red_SubCellInst2_LFInst_12_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_12_LFInst_1_U5  ( .A1(
        PermutationOutput2[51]), .A2(PermutationOutput2[50]), .ZN(
        \Red_SubCellInst2_LFInst_12_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst2_LFInst_12_LFInst_1_U4  ( .A1(PermutationOutput2[50]), .A2(\Red_SubCellInst2_LFInst_12_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst2_LFInst_12_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_12_LFInst_1_U3  ( .A(
        PermutationOutput2[48]), .B(PermutationOutput2[51]), .ZN(
        \Red_SubCellInst2_LFInst_12_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_12_LFInst_2_U10  ( .A1(
        \Red_SubCellInst2_LFInst_12_LFInst_2_n19 ), .A2(
        \Red_SubCellInst2_LFInst_12_LFInst_2_n18 ), .ZN(Red_Feedback2[50]) );
  AND2_X1 \Red_SubCellInst2_LFInst_12_LFInst_2_U9  ( .A1(
        \Red_SubCellInst2_LFInst_12_LFInst_2_n17 ), .A2(PermutationOutput2[48]), .ZN(\Red_SubCellInst2_LFInst_12_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_12_LFInst_2_U8  ( .A1(
        PermutationOutput2[50]), .A2(PermutationOutput2[49]), .ZN(
        \Red_SubCellInst2_LFInst_12_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_12_LFInst_2_U7  ( .A(
        \Red_SubCellInst2_LFInst_12_LFInst_2_n16 ), .B(
        \Red_SubCellInst2_LFInst_12_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst2_LFInst_12_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_12_LFInst_2_U6  ( .A1(
        PermutationOutput2[51]), .A2(\Red_SubCellInst2_LFInst_12_LFInst_2_n14 ), .ZN(\Red_SubCellInst2_LFInst_12_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst2_LFInst_12_LFInst_2_U5  ( .A(PermutationOutput2[49]), 
        .ZN(\Red_SubCellInst2_LFInst_12_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_12_LFInst_2_U4  ( .A1(
        PermutationOutput2[50]), .A2(\Red_SubCellInst2_LFInst_12_LFInst_2_n13 ), .ZN(\Red_SubCellInst2_LFInst_12_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst2_LFInst_12_LFInst_2_U3  ( .A(PermutationOutput2[48]), 
        .ZN(\Red_SubCellInst2_LFInst_12_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_12_LFInst_3_U6  ( .A(
        PermutationOutput2[49]), .B(\Red_SubCellInst2_LFInst_12_LFInst_3_n8 ), 
        .ZN(Red_Feedback2[51]) );
  NOR2_X1 \Red_SubCellInst2_LFInst_12_LFInst_3_U5  ( .A1(
        \Red_SubCellInst2_LFInst_12_LFInst_3_n7 ), .A2(
        \Red_SubCellInst2_LFInst_12_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst2_LFInst_12_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_12_LFInst_3_U4  ( .A1(
        PermutationOutput2[50]), .A2(PermutationOutput2[51]), .ZN(
        \Red_SubCellInst2_LFInst_12_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst2_LFInst_12_LFInst_3_U3  ( .A1(
        PermutationOutput2[51]), .A2(PermutationOutput2[48]), .ZN(
        \Red_SubCellInst2_LFInst_12_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_13_LFInst_0_U10  ( .A1(
        \Red_SubCellInst2_LFInst_13_LFInst_0_n14 ), .A2(
        \Red_SubCellInst2_LFInst_13_LFInst_0_n13 ), .ZN(Red_Feedback2[52]) );
  NAND2_X1 \Red_SubCellInst2_LFInst_13_LFInst_0_U9  ( .A1(
        PermutationOutput2[52]), .A2(\Red_SubCellInst2_LFInst_13_LFInst_0_n12 ), .ZN(\Red_SubCellInst2_LFInst_13_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_13_LFInst_0_U8  ( .A1(
        \Red_SubCellInst2_LFInst_13_LFInst_0_n11 ), .A2(PermutationOutput2[54]), .ZN(\Red_SubCellInst2_LFInst_13_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_13_LFInst_0_U7  ( .A(
        \Red_SubCellInst2_LFInst_13_LFInst_0_n10 ), .B(
        \Red_SubCellInst2_LFInst_13_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst2_LFInst_13_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_13_LFInst_0_U6  ( .A1(
        PermutationOutput2[55]), .A2(\Red_SubCellInst2_LFInst_13_LFInst_0_n11 ), .ZN(\Red_SubCellInst2_LFInst_13_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst2_LFInst_13_LFInst_0_U5  ( .A(PermutationOutput2[53]), 
        .ZN(\Red_SubCellInst2_LFInst_13_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_13_LFInst_0_U4  ( .A1(
        PermutationOutput2[54]), .A2(\Red_SubCellInst2_LFInst_13_LFInst_0_n8 ), 
        .ZN(\Red_SubCellInst2_LFInst_13_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst2_LFInst_13_LFInst_0_U3  ( .A(PermutationOutput2[52]), 
        .ZN(\Red_SubCellInst2_LFInst_13_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_13_LFInst_1_U8  ( .A1(
        \Red_SubCellInst2_LFInst_13_LFInst_1_n15 ), .A2(
        \Red_SubCellInst2_LFInst_13_LFInst_1_n14 ), .ZN(Red_Feedback2[53]) );
  NAND2_X1 \Red_SubCellInst2_LFInst_13_LFInst_1_U7  ( .A1(
        \Red_SubCellInst2_LFInst_13_LFInst_1_n13 ), .A2(PermutationOutput2[53]), .ZN(\Red_SubCellInst2_LFInst_13_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_13_LFInst_1_U6  ( .A1(
        \Red_SubCellInst2_LFInst_13_LFInst_1_n12 ), .A2(PermutationOutput2[52]), .ZN(\Red_SubCellInst2_LFInst_13_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_13_LFInst_1_U5  ( .A1(
        PermutationOutput2[55]), .A2(PermutationOutput2[54]), .ZN(
        \Red_SubCellInst2_LFInst_13_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst2_LFInst_13_LFInst_1_U4  ( .A1(PermutationOutput2[54]), .A2(\Red_SubCellInst2_LFInst_13_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst2_LFInst_13_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_13_LFInst_1_U3  ( .A(
        PermutationOutput2[52]), .B(PermutationOutput2[55]), .ZN(
        \Red_SubCellInst2_LFInst_13_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_13_LFInst_2_U10  ( .A1(
        \Red_SubCellInst2_LFInst_13_LFInst_2_n19 ), .A2(
        \Red_SubCellInst2_LFInst_13_LFInst_2_n18 ), .ZN(Red_Feedback2[54]) );
  AND2_X1 \Red_SubCellInst2_LFInst_13_LFInst_2_U9  ( .A1(
        \Red_SubCellInst2_LFInst_13_LFInst_2_n17 ), .A2(PermutationOutput2[52]), .ZN(\Red_SubCellInst2_LFInst_13_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_13_LFInst_2_U8  ( .A1(
        PermutationOutput2[54]), .A2(PermutationOutput2[53]), .ZN(
        \Red_SubCellInst2_LFInst_13_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_13_LFInst_2_U7  ( .A(
        \Red_SubCellInst2_LFInst_13_LFInst_2_n16 ), .B(
        \Red_SubCellInst2_LFInst_13_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst2_LFInst_13_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_13_LFInst_2_U6  ( .A1(
        PermutationOutput2[55]), .A2(\Red_SubCellInst2_LFInst_13_LFInst_2_n14 ), .ZN(\Red_SubCellInst2_LFInst_13_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst2_LFInst_13_LFInst_2_U5  ( .A(PermutationOutput2[53]), 
        .ZN(\Red_SubCellInst2_LFInst_13_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_13_LFInst_2_U4  ( .A1(
        PermutationOutput2[54]), .A2(\Red_SubCellInst2_LFInst_13_LFInst_2_n13 ), .ZN(\Red_SubCellInst2_LFInst_13_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst2_LFInst_13_LFInst_2_U3  ( .A(PermutationOutput2[52]), 
        .ZN(\Red_SubCellInst2_LFInst_13_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_13_LFInst_3_U6  ( .A(
        PermutationOutput2[53]), .B(\Red_SubCellInst2_LFInst_13_LFInst_3_n8 ), 
        .ZN(Red_Feedback2[55]) );
  NOR2_X1 \Red_SubCellInst2_LFInst_13_LFInst_3_U5  ( .A1(
        \Red_SubCellInst2_LFInst_13_LFInst_3_n7 ), .A2(
        \Red_SubCellInst2_LFInst_13_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst2_LFInst_13_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_13_LFInst_3_U4  ( .A1(
        PermutationOutput2[54]), .A2(PermutationOutput2[55]), .ZN(
        \Red_SubCellInst2_LFInst_13_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst2_LFInst_13_LFInst_3_U3  ( .A1(
        PermutationOutput2[55]), .A2(PermutationOutput2[52]), .ZN(
        \Red_SubCellInst2_LFInst_13_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_14_LFInst_0_U10  ( .A1(
        \Red_SubCellInst2_LFInst_14_LFInst_0_n14 ), .A2(
        \Red_SubCellInst2_LFInst_14_LFInst_0_n13 ), .ZN(Red_Feedback2[56]) );
  NAND2_X1 \Red_SubCellInst2_LFInst_14_LFInst_0_U9  ( .A1(
        PermutationOutput2[56]), .A2(\Red_SubCellInst2_LFInst_14_LFInst_0_n12 ), .ZN(\Red_SubCellInst2_LFInst_14_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_14_LFInst_0_U8  ( .A1(
        \Red_SubCellInst2_LFInst_14_LFInst_0_n11 ), .A2(PermutationOutput2[58]), .ZN(\Red_SubCellInst2_LFInst_14_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_14_LFInst_0_U7  ( .A(
        \Red_SubCellInst2_LFInst_14_LFInst_0_n10 ), .B(
        \Red_SubCellInst2_LFInst_14_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst2_LFInst_14_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_14_LFInst_0_U6  ( .A1(
        PermutationOutput2[59]), .A2(\Red_SubCellInst2_LFInst_14_LFInst_0_n11 ), .ZN(\Red_SubCellInst2_LFInst_14_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst2_LFInst_14_LFInst_0_U5  ( .A(PermutationOutput2[57]), 
        .ZN(\Red_SubCellInst2_LFInst_14_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_14_LFInst_0_U4  ( .A1(
        PermutationOutput2[58]), .A2(\Red_SubCellInst2_LFInst_14_LFInst_0_n8 ), 
        .ZN(\Red_SubCellInst2_LFInst_14_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst2_LFInst_14_LFInst_0_U3  ( .A(PermutationOutput2[56]), 
        .ZN(\Red_SubCellInst2_LFInst_14_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_14_LFInst_1_U8  ( .A1(
        \Red_SubCellInst2_LFInst_14_LFInst_1_n15 ), .A2(
        \Red_SubCellInst2_LFInst_14_LFInst_1_n14 ), .ZN(Red_Feedback2[57]) );
  NAND2_X1 \Red_SubCellInst2_LFInst_14_LFInst_1_U7  ( .A1(
        \Red_SubCellInst2_LFInst_14_LFInst_1_n13 ), .A2(PermutationOutput2[57]), .ZN(\Red_SubCellInst2_LFInst_14_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_14_LFInst_1_U6  ( .A1(
        \Red_SubCellInst2_LFInst_14_LFInst_1_n12 ), .A2(PermutationOutput2[56]), .ZN(\Red_SubCellInst2_LFInst_14_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_14_LFInst_1_U5  ( .A1(
        PermutationOutput2[59]), .A2(PermutationOutput2[58]), .ZN(
        \Red_SubCellInst2_LFInst_14_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst2_LFInst_14_LFInst_1_U4  ( .A1(PermutationOutput2[58]), .A2(\Red_SubCellInst2_LFInst_14_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst2_LFInst_14_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_14_LFInst_1_U3  ( .A(
        PermutationOutput2[56]), .B(PermutationOutput2[59]), .ZN(
        \Red_SubCellInst2_LFInst_14_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_14_LFInst_2_U10  ( .A1(
        \Red_SubCellInst2_LFInst_14_LFInst_2_n19 ), .A2(
        \Red_SubCellInst2_LFInst_14_LFInst_2_n18 ), .ZN(Red_Feedback2[58]) );
  AND2_X1 \Red_SubCellInst2_LFInst_14_LFInst_2_U9  ( .A1(
        \Red_SubCellInst2_LFInst_14_LFInst_2_n17 ), .A2(PermutationOutput2[56]), .ZN(\Red_SubCellInst2_LFInst_14_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_14_LFInst_2_U8  ( .A1(
        PermutationOutput2[58]), .A2(PermutationOutput2[57]), .ZN(
        \Red_SubCellInst2_LFInst_14_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_14_LFInst_2_U7  ( .A(
        \Red_SubCellInst2_LFInst_14_LFInst_2_n16 ), .B(
        \Red_SubCellInst2_LFInst_14_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst2_LFInst_14_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_14_LFInst_2_U6  ( .A1(
        PermutationOutput2[59]), .A2(\Red_SubCellInst2_LFInst_14_LFInst_2_n14 ), .ZN(\Red_SubCellInst2_LFInst_14_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst2_LFInst_14_LFInst_2_U5  ( .A(PermutationOutput2[57]), 
        .ZN(\Red_SubCellInst2_LFInst_14_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_14_LFInst_2_U4  ( .A1(
        PermutationOutput2[58]), .A2(\Red_SubCellInst2_LFInst_14_LFInst_2_n13 ), .ZN(\Red_SubCellInst2_LFInst_14_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst2_LFInst_14_LFInst_2_U3  ( .A(PermutationOutput2[56]), 
        .ZN(\Red_SubCellInst2_LFInst_14_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_14_LFInst_3_U6  ( .A(
        PermutationOutput2[57]), .B(\Red_SubCellInst2_LFInst_14_LFInst_3_n8 ), 
        .ZN(Red_Feedback2[59]) );
  NOR2_X1 \Red_SubCellInst2_LFInst_14_LFInst_3_U5  ( .A1(
        \Red_SubCellInst2_LFInst_14_LFInst_3_n7 ), .A2(
        \Red_SubCellInst2_LFInst_14_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst2_LFInst_14_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_14_LFInst_3_U4  ( .A1(
        PermutationOutput2[58]), .A2(PermutationOutput2[59]), .ZN(
        \Red_SubCellInst2_LFInst_14_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst2_LFInst_14_LFInst_3_U3  ( .A1(
        PermutationOutput2[59]), .A2(PermutationOutput2[56]), .ZN(
        \Red_SubCellInst2_LFInst_14_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_15_LFInst_0_U10  ( .A1(
        \Red_SubCellInst2_LFInst_15_LFInst_0_n14 ), .A2(
        \Red_SubCellInst2_LFInst_15_LFInst_0_n13 ), .ZN(Red_Feedback2[60]) );
  NAND2_X1 \Red_SubCellInst2_LFInst_15_LFInst_0_U9  ( .A1(
        PermutationOutput2[60]), .A2(\Red_SubCellInst2_LFInst_15_LFInst_0_n12 ), .ZN(\Red_SubCellInst2_LFInst_15_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_15_LFInst_0_U8  ( .A1(
        \Red_SubCellInst2_LFInst_15_LFInst_0_n11 ), .A2(PermutationOutput2[62]), .ZN(\Red_SubCellInst2_LFInst_15_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_15_LFInst_0_U7  ( .A(
        \Red_SubCellInst2_LFInst_15_LFInst_0_n10 ), .B(
        \Red_SubCellInst2_LFInst_15_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst2_LFInst_15_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_15_LFInst_0_U6  ( .A1(
        PermutationOutput2[63]), .A2(\Red_SubCellInst2_LFInst_15_LFInst_0_n11 ), .ZN(\Red_SubCellInst2_LFInst_15_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst2_LFInst_15_LFInst_0_U5  ( .A(PermutationOutput2[61]), 
        .ZN(\Red_SubCellInst2_LFInst_15_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_15_LFInst_0_U4  ( .A1(
        PermutationOutput2[62]), .A2(\Red_SubCellInst2_LFInst_15_LFInst_0_n8 ), 
        .ZN(\Red_SubCellInst2_LFInst_15_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst2_LFInst_15_LFInst_0_U3  ( .A(PermutationOutput2[60]), 
        .ZN(\Red_SubCellInst2_LFInst_15_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_15_LFInst_1_U8  ( .A1(
        \Red_SubCellInst2_LFInst_15_LFInst_1_n15 ), .A2(
        \Red_SubCellInst2_LFInst_15_LFInst_1_n14 ), .ZN(Red_Feedback2[61]) );
  NAND2_X1 \Red_SubCellInst2_LFInst_15_LFInst_1_U7  ( .A1(
        \Red_SubCellInst2_LFInst_15_LFInst_1_n13 ), .A2(PermutationOutput2[61]), .ZN(\Red_SubCellInst2_LFInst_15_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_15_LFInst_1_U6  ( .A1(
        \Red_SubCellInst2_LFInst_15_LFInst_1_n12 ), .A2(PermutationOutput2[60]), .ZN(\Red_SubCellInst2_LFInst_15_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_15_LFInst_1_U5  ( .A1(
        PermutationOutput2[63]), .A2(PermutationOutput2[62]), .ZN(
        \Red_SubCellInst2_LFInst_15_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst2_LFInst_15_LFInst_1_U4  ( .A1(PermutationOutput2[62]), .A2(\Red_SubCellInst2_LFInst_15_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst2_LFInst_15_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_15_LFInst_1_U3  ( .A(
        PermutationOutput2[60]), .B(PermutationOutput2[63]), .ZN(
        \Red_SubCellInst2_LFInst_15_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_15_LFInst_2_U10  ( .A1(
        \Red_SubCellInst2_LFInst_15_LFInst_2_n19 ), .A2(
        \Red_SubCellInst2_LFInst_15_LFInst_2_n18 ), .ZN(Red_Feedback2[62]) );
  AND2_X1 \Red_SubCellInst2_LFInst_15_LFInst_2_U9  ( .A1(
        \Red_SubCellInst2_LFInst_15_LFInst_2_n17 ), .A2(PermutationOutput2[60]), .ZN(\Red_SubCellInst2_LFInst_15_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_15_LFInst_2_U8  ( .A1(
        PermutationOutput2[62]), .A2(PermutationOutput2[61]), .ZN(
        \Red_SubCellInst2_LFInst_15_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_15_LFInst_2_U7  ( .A(
        \Red_SubCellInst2_LFInst_15_LFInst_2_n16 ), .B(
        \Red_SubCellInst2_LFInst_15_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst2_LFInst_15_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_15_LFInst_2_U6  ( .A1(
        PermutationOutput2[63]), .A2(\Red_SubCellInst2_LFInst_15_LFInst_2_n14 ), .ZN(\Red_SubCellInst2_LFInst_15_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst2_LFInst_15_LFInst_2_U5  ( .A(PermutationOutput2[61]), 
        .ZN(\Red_SubCellInst2_LFInst_15_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst2_LFInst_15_LFInst_2_U4  ( .A1(
        PermutationOutput2[62]), .A2(\Red_SubCellInst2_LFInst_15_LFInst_2_n13 ), .ZN(\Red_SubCellInst2_LFInst_15_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst2_LFInst_15_LFInst_2_U3  ( .A(PermutationOutput2[60]), 
        .ZN(\Red_SubCellInst2_LFInst_15_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst2_LFInst_15_LFInst_3_U6  ( .A(
        PermutationOutput2[61]), .B(\Red_SubCellInst2_LFInst_15_LFInst_3_n8 ), 
        .ZN(Red_Feedback2[63]) );
  NOR2_X1 \Red_SubCellInst2_LFInst_15_LFInst_3_U5  ( .A1(
        \Red_SubCellInst2_LFInst_15_LFInst_3_n7 ), .A2(
        \Red_SubCellInst2_LFInst_15_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst2_LFInst_15_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst2_LFInst_15_LFInst_3_U4  ( .A1(
        PermutationOutput2[62]), .A2(PermutationOutput2[63]), .ZN(
        \Red_SubCellInst2_LFInst_15_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst2_LFInst_15_LFInst_3_U3  ( .A1(
        PermutationOutput2[63]), .A2(PermutationOutput2[60]), .ZN(
        \Red_SubCellInst2_LFInst_15_LFInst_3_n7 ) );
  XNOR2_X1 \Red_MCInst3_XOR_r0_Inst_0_U2  ( .A(\Red_MCInst3_XOR_r0_Inst_0_n3 ), 
        .B(Red_MCOutput3[0]), .ZN(Red_MCOutput3[48]) );
  XNOR2_X1 \Red_MCInst3_XOR_r0_Inst_0_U1  ( .A(Red_Feedback2[48]), .B(
        Red_MCOutput3[16]), .ZN(\Red_MCInst3_XOR_r0_Inst_0_n3 ) );
  XOR2_X1 \Red_MCInst3_XOR_r1_Inst_0_U1  ( .A(Red_Feedback2[32]), .B(
        Red_MCOutput3[0]), .Z(Red_MCOutput3[32]) );
  XNOR2_X1 \Red_MCInst3_XOR_r0_Inst_1_U2  ( .A(\Red_MCInst3_XOR_r0_Inst_1_n3 ), 
        .B(Red_MCOutput3[1]), .ZN(Red_MCOutput3[49]) );
  XNOR2_X1 \Red_MCInst3_XOR_r0_Inst_1_U1  ( .A(Red_Feedback2[49]), .B(
        Red_MCOutput3[17]), .ZN(\Red_MCInst3_XOR_r0_Inst_1_n3 ) );
  XOR2_X1 \Red_MCInst3_XOR_r1_Inst_1_U1  ( .A(Red_Feedback2[33]), .B(
        Red_MCOutput3[1]), .Z(Red_MCOutput3[33]) );
  XNOR2_X1 \Red_MCInst3_XOR_r0_Inst_2_U2  ( .A(\Red_MCInst3_XOR_r0_Inst_2_n3 ), 
        .B(Red_MCOutput3[2]), .ZN(Red_MCOutput3[50]) );
  XNOR2_X1 \Red_MCInst3_XOR_r0_Inst_2_U1  ( .A(Red_Feedback2[50]), .B(
        Red_MCOutput3[18]), .ZN(\Red_MCInst3_XOR_r0_Inst_2_n3 ) );
  XOR2_X1 \Red_MCInst3_XOR_r1_Inst_2_U1  ( .A(Red_Feedback2[34]), .B(
        Red_MCOutput3[2]), .Z(Red_MCOutput3[34]) );
  XNOR2_X1 \Red_MCInst3_XOR_r0_Inst_3_U2  ( .A(\Red_MCInst3_XOR_r0_Inst_3_n3 ), 
        .B(Red_MCOutput3[3]), .ZN(Red_MCOutput3[51]) );
  XNOR2_X1 \Red_MCInst3_XOR_r0_Inst_3_U1  ( .A(Red_Feedback2[51]), .B(
        Red_MCOutput3[19]), .ZN(\Red_MCInst3_XOR_r0_Inst_3_n3 ) );
  XOR2_X1 \Red_MCInst3_XOR_r1_Inst_3_U1  ( .A(Red_Feedback2[35]), .B(
        Red_MCOutput3[3]), .Z(Red_MCOutput3[35]) );
  XNOR2_X1 \Red_MCInst3_XOR_r0_Inst_4_U2  ( .A(\Red_MCInst3_XOR_r0_Inst_4_n3 ), 
        .B(Red_MCOutput3[4]), .ZN(Red_MCOutput3[52]) );
  XNOR2_X1 \Red_MCInst3_XOR_r0_Inst_4_U1  ( .A(Red_Feedback2[52]), .B(
        Red_MCOutput3[20]), .ZN(\Red_MCInst3_XOR_r0_Inst_4_n3 ) );
  XOR2_X1 \Red_MCInst3_XOR_r1_Inst_4_U1  ( .A(Red_Feedback2[36]), .B(
        Red_MCOutput3[4]), .Z(Red_MCOutput3[36]) );
  XNOR2_X1 \Red_MCInst3_XOR_r0_Inst_5_U2  ( .A(\Red_MCInst3_XOR_r0_Inst_5_n3 ), 
        .B(Red_MCOutput3[5]), .ZN(Red_MCOutput3[53]) );
  XNOR2_X1 \Red_MCInst3_XOR_r0_Inst_5_U1  ( .A(Red_Feedback2[53]), .B(
        Red_MCOutput3[21]), .ZN(\Red_MCInst3_XOR_r0_Inst_5_n3 ) );
  XOR2_X1 \Red_MCInst3_XOR_r1_Inst_5_U1  ( .A(Red_Feedback2[37]), .B(
        Red_MCOutput3[5]), .Z(Red_MCOutput3[37]) );
  XNOR2_X1 \Red_MCInst3_XOR_r0_Inst_6_U2  ( .A(\Red_MCInst3_XOR_r0_Inst_6_n3 ), 
        .B(Red_MCOutput3[6]), .ZN(Red_MCOutput3[54]) );
  XNOR2_X1 \Red_MCInst3_XOR_r0_Inst_6_U1  ( .A(Red_Feedback2[54]), .B(
        Red_MCOutput3[22]), .ZN(\Red_MCInst3_XOR_r0_Inst_6_n3 ) );
  XOR2_X1 \Red_MCInst3_XOR_r1_Inst_6_U1  ( .A(Red_Feedback2[38]), .B(
        Red_MCOutput3[6]), .Z(Red_MCOutput3[38]) );
  XNOR2_X1 \Red_MCInst3_XOR_r0_Inst_7_U2  ( .A(\Red_MCInst3_XOR_r0_Inst_7_n3 ), 
        .B(Red_MCOutput3[7]), .ZN(Red_MCOutput3[55]) );
  XNOR2_X1 \Red_MCInst3_XOR_r0_Inst_7_U1  ( .A(Red_Feedback2[55]), .B(
        Red_MCOutput3[23]), .ZN(\Red_MCInst3_XOR_r0_Inst_7_n3 ) );
  XOR2_X1 \Red_MCInst3_XOR_r1_Inst_7_U1  ( .A(Red_Feedback2[39]), .B(
        Red_MCOutput3[7]), .Z(Red_MCOutput3[39]) );
  XNOR2_X1 \Red_MCInst3_XOR_r0_Inst_8_U2  ( .A(\Red_MCInst3_XOR_r0_Inst_8_n3 ), 
        .B(Red_MCOutput3[8]), .ZN(Red_MCOutput3[56]) );
  XNOR2_X1 \Red_MCInst3_XOR_r0_Inst_8_U1  ( .A(Red_Feedback2[56]), .B(
        Red_MCOutput3[24]), .ZN(\Red_MCInst3_XOR_r0_Inst_8_n3 ) );
  XOR2_X1 \Red_MCInst3_XOR_r1_Inst_8_U1  ( .A(Red_Feedback2[40]), .B(
        Red_MCOutput3[8]), .Z(Red_MCOutput3[40]) );
  XNOR2_X1 \Red_MCInst3_XOR_r0_Inst_9_U2  ( .A(\Red_MCInst3_XOR_r0_Inst_9_n3 ), 
        .B(Red_MCOutput3[9]), .ZN(Red_MCOutput3[57]) );
  XNOR2_X1 \Red_MCInst3_XOR_r0_Inst_9_U1  ( .A(Red_Feedback2[57]), .B(
        Red_MCOutput3[25]), .ZN(\Red_MCInst3_XOR_r0_Inst_9_n3 ) );
  XOR2_X1 \Red_MCInst3_XOR_r1_Inst_9_U1  ( .A(Red_Feedback2[41]), .B(
        Red_MCOutput3[9]), .Z(Red_MCOutput3[41]) );
  XNOR2_X1 \Red_MCInst3_XOR_r0_Inst_10_U2  ( .A(
        \Red_MCInst3_XOR_r0_Inst_10_n3 ), .B(Red_MCOutput3[10]), .ZN(
        Red_MCOutput3[58]) );
  XNOR2_X1 \Red_MCInst3_XOR_r0_Inst_10_U1  ( .A(Red_Feedback2[58]), .B(
        Red_MCOutput3[26]), .ZN(\Red_MCInst3_XOR_r0_Inst_10_n3 ) );
  XOR2_X1 \Red_MCInst3_XOR_r1_Inst_10_U1  ( .A(Red_Feedback2[42]), .B(
        Red_MCOutput3[10]), .Z(Red_MCOutput3[42]) );
  XNOR2_X1 \Red_MCInst3_XOR_r0_Inst_11_U2  ( .A(
        \Red_MCInst3_XOR_r0_Inst_11_n3 ), .B(Red_MCOutput3[11]), .ZN(
        Red_MCOutput3[59]) );
  XNOR2_X1 \Red_MCInst3_XOR_r0_Inst_11_U1  ( .A(Red_Feedback2[59]), .B(
        Red_MCOutput3[27]), .ZN(\Red_MCInst3_XOR_r0_Inst_11_n3 ) );
  XOR2_X1 \Red_MCInst3_XOR_r1_Inst_11_U1  ( .A(Red_Feedback2[43]), .B(
        Red_MCOutput3[11]), .Z(Red_MCOutput3[43]) );
  XNOR2_X1 \Red_MCInst3_XOR_r0_Inst_12_U2  ( .A(
        \Red_MCInst3_XOR_r0_Inst_12_n3 ), .B(Red_MCOutput3[12]), .ZN(
        Red_MCOutput3[60]) );
  XNOR2_X1 \Red_MCInst3_XOR_r0_Inst_12_U1  ( .A(Red_Feedback2[60]), .B(
        Red_MCOutput3[28]), .ZN(\Red_MCInst3_XOR_r0_Inst_12_n3 ) );
  XOR2_X1 \Red_MCInst3_XOR_r1_Inst_12_U1  ( .A(Red_Feedback2[44]), .B(
        Red_MCOutput3[12]), .Z(Red_MCOutput3[44]) );
  XNOR2_X1 \Red_MCInst3_XOR_r0_Inst_13_U2  ( .A(
        \Red_MCInst3_XOR_r0_Inst_13_n3 ), .B(Red_MCOutput3[13]), .ZN(
        Red_MCOutput3[61]) );
  XNOR2_X1 \Red_MCInst3_XOR_r0_Inst_13_U1  ( .A(Red_Feedback2[61]), .B(
        Red_MCOutput3[29]), .ZN(\Red_MCInst3_XOR_r0_Inst_13_n3 ) );
  XOR2_X1 \Red_MCInst3_XOR_r1_Inst_13_U1  ( .A(Red_Feedback2[45]), .B(
        Red_MCOutput3[13]), .Z(Red_MCOutput3[45]) );
  XNOR2_X1 \Red_MCInst3_XOR_r0_Inst_14_U2  ( .A(
        \Red_MCInst3_XOR_r0_Inst_14_n3 ), .B(Red_MCOutput3[14]), .ZN(
        Red_MCOutput3[62]) );
  XNOR2_X1 \Red_MCInst3_XOR_r0_Inst_14_U1  ( .A(Red_Feedback2[62]), .B(
        Red_MCOutput3[30]), .ZN(\Red_MCInst3_XOR_r0_Inst_14_n3 ) );
  XOR2_X1 \Red_MCInst3_XOR_r1_Inst_14_U1  ( .A(Red_Feedback2[46]), .B(
        Red_MCOutput3[14]), .Z(Red_MCOutput3[46]) );
  XNOR2_X1 \Red_MCInst3_XOR_r0_Inst_15_U2  ( .A(
        \Red_MCInst3_XOR_r0_Inst_15_n3 ), .B(Red_MCOutput3[15]), .ZN(
        Red_MCOutput3[63]) );
  XNOR2_X1 \Red_MCInst3_XOR_r0_Inst_15_U1  ( .A(Red_Feedback2[63]), .B(
        Red_MCOutput3[31]), .ZN(\Red_MCInst3_XOR_r0_Inst_15_n3 ) );
  XOR2_X1 \Red_MCInst3_XOR_r1_Inst_15_U1  ( .A(Red_Feedback2[47]), .B(
        Red_MCOutput3[15]), .Z(Red_MCOutput3[47]) );
  XOR2_X1 \Red_AddKeyXOR13_XORInst_0_0_U1  ( .A(Red_MCOutput3[48]), .B(
        Red_K2[48]), .Z(Red_AddRoundKeyOutput3[48]) );
  XOR2_X1 \Red_AddKeyXOR13_XORInst_0_1_U1  ( .A(Red_MCOutput3[49]), .B(
        Red_K2[49]), .Z(Red_AddRoundKeyOutput3[49]) );
  XOR2_X1 \Red_AddKeyXOR13_XORInst_0_2_U1  ( .A(Red_MCOutput3[50]), .B(
        Red_K2[50]), .Z(Red_AddRoundKeyOutput3[50]) );
  XOR2_X1 \Red_AddKeyXOR13_XORInst_0_3_U1  ( .A(Red_MCOutput3[51]), .B(
        Red_K2[51]), .Z(Red_AddRoundKeyOutput3[51]) );
  XOR2_X1 \Red_AddKeyXOR13_XORInst_1_0_U1  ( .A(Red_MCOutput3[52]), .B(
        Red_K2[52]), .Z(Red_AddRoundKeyOutput3[52]) );
  XOR2_X1 \Red_AddKeyXOR13_XORInst_1_1_U1  ( .A(Red_MCOutput3[53]), .B(
        Red_K2[53]), .Z(Red_AddRoundKeyOutput3[53]) );
  XOR2_X1 \Red_AddKeyXOR13_XORInst_1_2_U1  ( .A(Red_MCOutput3[54]), .B(
        Red_K2[54]), .Z(Red_AddRoundKeyOutput3[54]) );
  XOR2_X1 \Red_AddKeyXOR13_XORInst_1_3_U1  ( .A(Red_MCOutput3[55]), .B(
        Red_K2[55]), .Z(Red_AddRoundKeyOutput3[55]) );
  XOR2_X1 \Red_AddKeyXOR13_XORInst_2_0_U1  ( .A(Red_MCOutput3[56]), .B(
        Red_K2[56]), .Z(Red_AddRoundKeyOutput3[56]) );
  XOR2_X1 \Red_AddKeyXOR13_XORInst_2_1_U1  ( .A(Red_MCOutput3[57]), .B(
        Red_K2[57]), .Z(Red_AddRoundKeyOutput3[57]) );
  XOR2_X1 \Red_AddKeyXOR13_XORInst_2_2_U1  ( .A(Red_MCOutput3[58]), .B(
        Red_K2[58]), .Z(Red_AddRoundKeyOutput3[58]) );
  XOR2_X1 \Red_AddKeyXOR13_XORInst_2_3_U1  ( .A(Red_MCOutput3[59]), .B(
        Red_K2[59]), .Z(Red_AddRoundKeyOutput3[59]) );
  XOR2_X1 \Red_AddKeyXOR13_XORInst_3_0_U1  ( .A(Red_MCOutput3[60]), .B(
        Red_K2[60]), .Z(Red_AddRoundKeyOutput3[60]) );
  XOR2_X1 \Red_AddKeyXOR13_XORInst_3_1_U1  ( .A(Red_MCOutput3[61]), .B(
        Red_K2[61]), .Z(Red_AddRoundKeyOutput3[61]) );
  XOR2_X1 \Red_AddKeyXOR13_XORInst_3_2_U1  ( .A(Red_MCOutput3[62]), .B(
        Red_K2[62]), .Z(Red_AddRoundKeyOutput3[62]) );
  XOR2_X1 \Red_AddKeyXOR13_XORInst_3_3_U1  ( .A(Red_MCOutput3[63]), .B(
        Red_K2[63]), .Z(Red_AddRoundKeyOutput3[63]) );
  XOR2_X1 \Red_AddKeyConstXOR3_XORInst_0_0_U1  ( .A(Red_K2[40]), .B(
        Red_MCOutput3[40]), .Z(Red_AddRoundKeyOutput3[40]) );
  XOR2_X1 \Red_AddKeyConstXOR3_XORInst_0_1_U1  ( .A(Red_K2[41]), .B(
        Red_MCOutput3[41]), .Z(Red_AddRoundKeyOutput3[41]) );
  XOR2_X1 \Red_AddKeyConstXOR3_XORInst_0_2_U1  ( .A(Red_K2[42]), .B(
        Red_MCOutput3[42]), .Z(Red_AddRoundKeyOutput3[42]) );
  XOR2_X1 \Red_AddKeyConstXOR3_XORInst_0_3_U1  ( .A(Red_K2[43]), .B(
        Red_MCOutput3[43]), .Z(Red_AddRoundKeyOutput3[43]) );
  XOR2_X1 \Red_AddKeyConstXOR3_XORInst_1_0_U1  ( .A(Red_K2[44]), .B(
        Red_MCOutput3[44]), .Z(Red_AddRoundKeyOutput3[44]) );
  XOR2_X1 \Red_AddKeyConstXOR3_XORInst_1_1_U1  ( .A(Red_K2[45]), .B(
        Red_MCOutput3[45]), .Z(Red_AddRoundKeyOutput3[45]) );
  XOR2_X1 \Red_AddKeyConstXOR3_XORInst_1_2_U1  ( .A(Red_K2[46]), .B(
        Red_MCOutput3[46]), .Z(Red_AddRoundKeyOutput3[46]) );
  XOR2_X1 \Red_AddKeyConstXOR3_XORInst_1_3_U1  ( .A(Red_K2[47]), .B(
        Red_MCOutput3[47]), .Z(Red_AddRoundKeyOutput3[47]) );
  XOR2_X1 \Red_AddKeyXOR23_XORInst_0_0_U1  ( .A(Red_MCOutput3[0]), .B(
        Red_K2[0]), .Z(Red_AddRoundKeyOutput3[0]) );
  XOR2_X1 \Red_AddKeyXOR23_XORInst_0_1_U1  ( .A(Red_MCOutput3[1]), .B(
        Red_K2[1]), .Z(Red_AddRoundKeyOutput3[1]) );
  XOR2_X1 \Red_AddKeyXOR23_XORInst_0_2_U1  ( .A(Red_MCOutput3[2]), .B(
        Red_K2[2]), .Z(Red_AddRoundKeyOutput3[2]) );
  XOR2_X1 \Red_AddKeyXOR23_XORInst_0_3_U1  ( .A(Red_MCOutput3[3]), .B(
        Red_K2[3]), .Z(Red_AddRoundKeyOutput3[3]) );
  XOR2_X1 \Red_AddKeyXOR23_XORInst_1_0_U1  ( .A(Red_MCOutput3[4]), .B(
        Red_K2[4]), .Z(Red_AddRoundKeyOutput3[4]) );
  XOR2_X1 \Red_AddKeyXOR23_XORInst_1_1_U1  ( .A(Red_MCOutput3[5]), .B(
        Red_K2[5]), .Z(Red_AddRoundKeyOutput3[5]) );
  XOR2_X1 \Red_AddKeyXOR23_XORInst_1_2_U1  ( .A(Red_MCOutput3[6]), .B(
        Red_K2[6]), .Z(Red_AddRoundKeyOutput3[6]) );
  XOR2_X1 \Red_AddKeyXOR23_XORInst_1_3_U1  ( .A(Red_MCOutput3[7]), .B(
        Red_K2[7]), .Z(Red_AddRoundKeyOutput3[7]) );
  XOR2_X1 \Red_AddKeyXOR23_XORInst_2_0_U1  ( .A(Red_MCOutput3[8]), .B(
        Red_K2[8]), .Z(Red_AddRoundKeyOutput3[8]) );
  XOR2_X1 \Red_AddKeyXOR23_XORInst_2_1_U1  ( .A(Red_MCOutput3[9]), .B(
        Red_K2[9]), .Z(Red_AddRoundKeyOutput3[9]) );
  XOR2_X1 \Red_AddKeyXOR23_XORInst_2_2_U1  ( .A(Red_MCOutput3[10]), .B(
        Red_K2[10]), .Z(Red_AddRoundKeyOutput3[10]) );
  XOR2_X1 \Red_AddKeyXOR23_XORInst_2_3_U1  ( .A(Red_MCOutput3[11]), .B(
        Red_K2[11]), .Z(Red_AddRoundKeyOutput3[11]) );
  XOR2_X1 \Red_AddKeyXOR23_XORInst_3_0_U1  ( .A(Red_MCOutput3[12]), .B(
        Red_K2[12]), .Z(Red_AddRoundKeyOutput3[12]) );
  XOR2_X1 \Red_AddKeyXOR23_XORInst_3_1_U1  ( .A(Red_MCOutput3[13]), .B(
        Red_K2[13]), .Z(Red_AddRoundKeyOutput3[13]) );
  XOR2_X1 \Red_AddKeyXOR23_XORInst_3_2_U1  ( .A(Red_MCOutput3[14]), .B(
        Red_K2[14]), .Z(Red_AddRoundKeyOutput3[14]) );
  XOR2_X1 \Red_AddKeyXOR23_XORInst_3_3_U1  ( .A(Red_MCOutput3[15]), .B(
        Red_K2[15]), .Z(Red_AddRoundKeyOutput3[15]) );
  XOR2_X1 \Red_AddKeyXOR23_XORInst_4_0_U1  ( .A(Red_MCOutput3[16]), .B(
        Red_K2[16]), .Z(Red_AddRoundKeyOutput3[16]) );
  XOR2_X1 \Red_AddKeyXOR23_XORInst_4_1_U1  ( .A(Red_MCOutput3[17]), .B(
        Red_K2[17]), .Z(Red_AddRoundKeyOutput3[17]) );
  XOR2_X1 \Red_AddKeyXOR23_XORInst_4_2_U1  ( .A(Red_MCOutput3[18]), .B(
        Red_K2[18]), .Z(Red_AddRoundKeyOutput3[18]) );
  XOR2_X1 \Red_AddKeyXOR23_XORInst_4_3_U1  ( .A(Red_MCOutput3[19]), .B(
        Red_K2[19]), .Z(Red_AddRoundKeyOutput3[19]) );
  XOR2_X1 \Red_AddKeyXOR23_XORInst_5_0_U1  ( .A(Red_MCOutput3[20]), .B(
        Red_K2[20]), .Z(Red_AddRoundKeyOutput3[20]) );
  XOR2_X1 \Red_AddKeyXOR23_XORInst_5_1_U1  ( .A(Red_MCOutput3[21]), .B(
        Red_K2[21]), .Z(Red_AddRoundKeyOutput3[21]) );
  XOR2_X1 \Red_AddKeyXOR23_XORInst_5_2_U1  ( .A(Red_MCOutput3[22]), .B(
        Red_K2[22]), .Z(Red_AddRoundKeyOutput3[22]) );
  XOR2_X1 \Red_AddKeyXOR23_XORInst_5_3_U1  ( .A(Red_MCOutput3[23]), .B(
        Red_K2[23]), .Z(Red_AddRoundKeyOutput3[23]) );
  XOR2_X1 \Red_AddKeyXOR23_XORInst_6_0_U1  ( .A(Red_MCOutput3[24]), .B(
        Red_K2[24]), .Z(Red_AddRoundKeyOutput3[24]) );
  XOR2_X1 \Red_AddKeyXOR23_XORInst_6_1_U1  ( .A(Red_MCOutput3[25]), .B(
        Red_K2[25]), .Z(Red_AddRoundKeyOutput3[25]) );
  XOR2_X1 \Red_AddKeyXOR23_XORInst_6_2_U1  ( .A(Red_MCOutput3[26]), .B(
        Red_K2[26]), .Z(Red_AddRoundKeyOutput3[26]) );
  XOR2_X1 \Red_AddKeyXOR23_XORInst_6_3_U1  ( .A(Red_MCOutput3[27]), .B(
        Red_K2[27]), .Z(Red_AddRoundKeyOutput3[27]) );
  XOR2_X1 \Red_AddKeyXOR23_XORInst_7_0_U1  ( .A(Red_MCOutput3[28]), .B(
        Red_K2[28]), .Z(Red_AddRoundKeyOutput3[28]) );
  XOR2_X1 \Red_AddKeyXOR23_XORInst_7_1_U1  ( .A(Red_MCOutput3[29]), .B(
        Red_K2[29]), .Z(Red_AddRoundKeyOutput3[29]) );
  XOR2_X1 \Red_AddKeyXOR23_XORInst_7_2_U1  ( .A(Red_MCOutput3[30]), .B(
        Red_K2[30]), .Z(Red_AddRoundKeyOutput3[30]) );
  XOR2_X1 \Red_AddKeyXOR23_XORInst_7_3_U1  ( .A(Red_MCOutput3[31]), .B(
        Red_K2[31]), .Z(Red_AddRoundKeyOutput3[31]) );
  XOR2_X1 \Red_AddKeyXOR23_XORInst_8_0_U1  ( .A(Red_MCOutput3[32]), .B(
        Red_K2[32]), .Z(Red_AddRoundKeyOutput3[32]) );
  XOR2_X1 \Red_AddKeyXOR23_XORInst_8_1_U1  ( .A(Red_MCOutput3[33]), .B(
        Red_K2[33]), .Z(Red_AddRoundKeyOutput3[33]) );
  XOR2_X1 \Red_AddKeyXOR23_XORInst_8_2_U1  ( .A(Red_MCOutput3[34]), .B(
        Red_K2[34]), .Z(Red_AddRoundKeyOutput3[34]) );
  XOR2_X1 \Red_AddKeyXOR23_XORInst_8_3_U1  ( .A(Red_MCOutput3[35]), .B(
        Red_K2[35]), .Z(Red_AddRoundKeyOutput3[35]) );
  XOR2_X1 \Red_AddKeyXOR23_XORInst_9_0_U1  ( .A(Red_MCOutput3[36]), .B(
        Red_K2[36]), .Z(Red_AddRoundKeyOutput3[36]) );
  XOR2_X1 \Red_AddKeyXOR23_XORInst_9_1_U1  ( .A(Red_MCOutput3[37]), .B(
        Red_K2[37]), .Z(Red_AddRoundKeyOutput3[37]) );
  XOR2_X1 \Red_AddKeyXOR23_XORInst_9_2_U1  ( .A(Red_MCOutput3[38]), .B(
        Red_K2[38]), .Z(Red_AddRoundKeyOutput3[38]) );
  XOR2_X1 \Red_AddKeyXOR23_XORInst_9_3_U1  ( .A(Red_MCOutput3[39]), .B(
        Red_K2[39]), .Z(Red_AddRoundKeyOutput3[39]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[0]  ( .D(Red_AddRoundKeyOutput3[0]), .CK(clk), .Q(Red_StateRegOutput3[0]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[1]  ( .D(Red_AddRoundKeyOutput3[1]), .CK(clk), .Q(Red_StateRegOutput3[1]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[2]  ( .D(Red_AddRoundKeyOutput3[2]), .CK(clk), .Q(Red_StateRegOutput3[2]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[3]  ( .D(Red_AddRoundKeyOutput3[3]), .CK(clk), .Q(Red_StateRegOutput3[3]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[4]  ( .D(Red_AddRoundKeyOutput3[4]), .CK(clk), .Q(Red_StateRegOutput3[4]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[5]  ( .D(Red_AddRoundKeyOutput3[5]), .CK(clk), .Q(Red_StateRegOutput3[5]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[6]  ( .D(Red_AddRoundKeyOutput3[6]), .CK(clk), .Q(Red_StateRegOutput3[6]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[7]  ( .D(Red_AddRoundKeyOutput3[7]), .CK(clk), .Q(Red_StateRegOutput3[7]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[8]  ( .D(Red_AddRoundKeyOutput3[8]), .CK(clk), .Q(Red_StateRegOutput3[8]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[9]  ( .D(Red_AddRoundKeyOutput3[9]), .CK(clk), .Q(Red_StateRegOutput3[9]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[10]  ( .D(
        Red_AddRoundKeyOutput3[10]), .CK(clk), .Q(Red_StateRegOutput3[10]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[11]  ( .D(
        Red_AddRoundKeyOutput3[11]), .CK(clk), .Q(Red_StateRegOutput3[11]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[12]  ( .D(
        Red_AddRoundKeyOutput3[12]), .CK(clk), .Q(Red_StateRegOutput3[12]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[13]  ( .D(
        Red_AddRoundKeyOutput3[13]), .CK(clk), .Q(Red_StateRegOutput3[13]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[14]  ( .D(
        Red_AddRoundKeyOutput3[14]), .CK(clk), .Q(Red_StateRegOutput3[14]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[15]  ( .D(
        Red_AddRoundKeyOutput3[15]), .CK(clk), .Q(Red_StateRegOutput3[15]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[16]  ( .D(
        Red_AddRoundKeyOutput3[16]), .CK(clk), .Q(Red_StateRegOutput3[16]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[17]  ( .D(
        Red_AddRoundKeyOutput3[17]), .CK(clk), .Q(Red_StateRegOutput3[17]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[18]  ( .D(
        Red_AddRoundKeyOutput3[18]), .CK(clk), .Q(Red_StateRegOutput3[18]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[19]  ( .D(
        Red_AddRoundKeyOutput3[19]), .CK(clk), .Q(Red_StateRegOutput3[19]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[20]  ( .D(
        Red_AddRoundKeyOutput3[20]), .CK(clk), .Q(Red_StateRegOutput3[20]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[21]  ( .D(
        Red_AddRoundKeyOutput3[21]), .CK(clk), .Q(Red_StateRegOutput3[21]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[22]  ( .D(
        Red_AddRoundKeyOutput3[22]), .CK(clk), .Q(Red_StateRegOutput3[22]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[23]  ( .D(
        Red_AddRoundKeyOutput3[23]), .CK(clk), .Q(Red_StateRegOutput3[23]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[24]  ( .D(
        Red_AddRoundKeyOutput3[24]), .CK(clk), .Q(Red_StateRegOutput3[24]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[25]  ( .D(
        Red_AddRoundKeyOutput3[25]), .CK(clk), .Q(Red_StateRegOutput3[25]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[26]  ( .D(
        Red_AddRoundKeyOutput3[26]), .CK(clk), .Q(Red_StateRegOutput3[26]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[27]  ( .D(
        Red_AddRoundKeyOutput3[27]), .CK(clk), .Q(Red_StateRegOutput3[27]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[28]  ( .D(
        Red_AddRoundKeyOutput3[28]), .CK(clk), .Q(Red_StateRegOutput3[28]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[29]  ( .D(
        Red_AddRoundKeyOutput3[29]), .CK(clk), .Q(Red_StateRegOutput3[29]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[30]  ( .D(
        Red_AddRoundKeyOutput3[30]), .CK(clk), .Q(Red_StateRegOutput3[30]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[31]  ( .D(
        Red_AddRoundKeyOutput3[31]), .CK(clk), .Q(Red_StateRegOutput3[31]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[32]  ( .D(
        Red_AddRoundKeyOutput3[32]), .CK(clk), .Q(Red_StateRegOutput3[32]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[33]  ( .D(
        Red_AddRoundKeyOutput3[33]), .CK(clk), .Q(Red_StateRegOutput3[33]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[34]  ( .D(
        Red_AddRoundKeyOutput3[34]), .CK(clk), .Q(Red_StateRegOutput3[34]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[35]  ( .D(
        Red_AddRoundKeyOutput3[35]), .CK(clk), .Q(Red_StateRegOutput3[35]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[36]  ( .D(
        Red_AddRoundKeyOutput3[36]), .CK(clk), .Q(Red_StateRegOutput3[36]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[37]  ( .D(
        Red_AddRoundKeyOutput3[37]), .CK(clk), .Q(Red_StateRegOutput3[37]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[38]  ( .D(
        Red_AddRoundKeyOutput3[38]), .CK(clk), .Q(Red_StateRegOutput3[38]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[39]  ( .D(
        Red_AddRoundKeyOutput3[39]), .CK(clk), .Q(Red_StateRegOutput3[39]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[40]  ( .D(
        Red_AddRoundKeyOutput3[40]), .CK(clk), .Q(Red_StateRegOutput3[40]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[41]  ( .D(
        Red_AddRoundKeyOutput3[41]), .CK(clk), .Q(Red_StateRegOutput3[41]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[42]  ( .D(
        Red_AddRoundKeyOutput3[42]), .CK(clk), .Q(Red_StateRegOutput3[42]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[43]  ( .D(
        Red_AddRoundKeyOutput3[43]), .CK(clk), .Q(Red_StateRegOutput3[43]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[44]  ( .D(
        Red_AddRoundKeyOutput3[44]), .CK(clk), .Q(Red_StateRegOutput3[44]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[45]  ( .D(
        Red_AddRoundKeyOutput3[45]), .CK(clk), .Q(Red_StateRegOutput3[45]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[46]  ( .D(
        Red_AddRoundKeyOutput3[46]), .CK(clk), .Q(Red_StateRegOutput3[46]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[47]  ( .D(
        Red_AddRoundKeyOutput3[47]), .CK(clk), .Q(Red_StateRegOutput3[47]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[48]  ( .D(
        Red_AddRoundKeyOutput3[48]), .CK(clk), .Q(Red_StateRegOutput3[48]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[49]  ( .D(
        Red_AddRoundKeyOutput3[49]), .CK(clk), .Q(Red_StateRegOutput3[49]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[50]  ( .D(
        Red_AddRoundKeyOutput3[50]), .CK(clk), .Q(Red_StateRegOutput3[50]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[51]  ( .D(
        Red_AddRoundKeyOutput3[51]), .CK(clk), .Q(Red_StateRegOutput3[51]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[52]  ( .D(
        Red_AddRoundKeyOutput3[52]), .CK(clk), .Q(Red_StateRegOutput3[52]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[53]  ( .D(
        Red_AddRoundKeyOutput3[53]), .CK(clk), .Q(Red_StateRegOutput3[53]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[54]  ( .D(
        Red_AddRoundKeyOutput3[54]), .CK(clk), .Q(Red_StateRegOutput3[54]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[55]  ( .D(
        Red_AddRoundKeyOutput3[55]), .CK(clk), .Q(Red_StateRegOutput3[55]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[56]  ( .D(
        Red_AddRoundKeyOutput3[56]), .CK(clk), .Q(Red_StateRegOutput3[56]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[57]  ( .D(
        Red_AddRoundKeyOutput3[57]), .CK(clk), .Q(Red_StateRegOutput3[57]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[58]  ( .D(
        Red_AddRoundKeyOutput3[58]), .CK(clk), .Q(Red_StateRegOutput3[58]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[59]  ( .D(
        Red_AddRoundKeyOutput3[59]), .CK(clk), .Q(Red_StateRegOutput3[59]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[60]  ( .D(
        Red_AddRoundKeyOutput3[60]), .CK(clk), .Q(Red_StateRegOutput3[60]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[61]  ( .D(
        Red_AddRoundKeyOutput3[61]), .CK(clk), .Q(Red_StateRegOutput3[61]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[62]  ( .D(
        Red_AddRoundKeyOutput3[62]), .CK(clk), .Q(Red_StateRegOutput3[62]) );
  DFF_X1 \Red_StateReg3_s_current_state_reg[63]  ( .D(
        Red_AddRoundKeyOutput3[63]), .CK(clk), .Q(Red_StateRegOutput3[63]) );
  NAND2_X1 \Red_SubCellInst3_LFInst_0_LFInst_0_U10  ( .A1(
        \Red_SubCellInst3_LFInst_0_LFInst_0_n14 ), .A2(
        \Red_SubCellInst3_LFInst_0_LFInst_0_n13 ), .ZN(Red_Feedback3[0]) );
  NAND2_X1 \Red_SubCellInst3_LFInst_0_LFInst_0_U9  ( .A1(PermutationOutput3[0]), .A2(\Red_SubCellInst3_LFInst_0_LFInst_0_n12 ), .ZN(
        \Red_SubCellInst3_LFInst_0_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_0_LFInst_0_U8  ( .A1(
        \Red_SubCellInst3_LFInst_0_LFInst_0_n11 ), .A2(PermutationOutput3[2]), 
        .ZN(\Red_SubCellInst3_LFInst_0_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_0_LFInst_0_U7  ( .A(
        \Red_SubCellInst3_LFInst_0_LFInst_0_n10 ), .B(
        \Red_SubCellInst3_LFInst_0_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst3_LFInst_0_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_0_LFInst_0_U6  ( .A1(PermutationOutput3[3]), .A2(\Red_SubCellInst3_LFInst_0_LFInst_0_n11 ), .ZN(
        \Red_SubCellInst3_LFInst_0_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst3_LFInst_0_LFInst_0_U5  ( .A(PermutationOutput3[1]), 
        .ZN(\Red_SubCellInst3_LFInst_0_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_0_LFInst_0_U4  ( .A1(PermutationOutput3[2]), .A2(\Red_SubCellInst3_LFInst_0_LFInst_0_n8 ), .ZN(
        \Red_SubCellInst3_LFInst_0_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst3_LFInst_0_LFInst_0_U3  ( .A(PermutationOutput3[0]), 
        .ZN(\Red_SubCellInst3_LFInst_0_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_0_LFInst_1_U8  ( .A1(
        \Red_SubCellInst3_LFInst_0_LFInst_1_n15 ), .A2(
        \Red_SubCellInst3_LFInst_0_LFInst_1_n14 ), .ZN(Red_Feedback3[1]) );
  NAND2_X1 \Red_SubCellInst3_LFInst_0_LFInst_1_U7  ( .A1(
        \Red_SubCellInst3_LFInst_0_LFInst_1_n13 ), .A2(PermutationOutput3[1]), 
        .ZN(\Red_SubCellInst3_LFInst_0_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_0_LFInst_1_U6  ( .A1(
        \Red_SubCellInst3_LFInst_0_LFInst_1_n12 ), .A2(PermutationOutput3[0]), 
        .ZN(\Red_SubCellInst3_LFInst_0_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_0_LFInst_1_U5  ( .A1(PermutationOutput3[3]), .A2(PermutationOutput3[2]), .ZN(\Red_SubCellInst3_LFInst_0_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst3_LFInst_0_LFInst_1_U4  ( .A1(PermutationOutput3[2]), 
        .A2(\Red_SubCellInst3_LFInst_0_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst3_LFInst_0_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_0_LFInst_1_U3  ( .A(PermutationOutput3[0]), 
        .B(PermutationOutput3[3]), .ZN(
        \Red_SubCellInst3_LFInst_0_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_0_LFInst_2_U10  ( .A1(
        \Red_SubCellInst3_LFInst_0_LFInst_2_n19 ), .A2(
        \Red_SubCellInst3_LFInst_0_LFInst_2_n18 ), .ZN(Red_Feedback3[2]) );
  AND2_X1 \Red_SubCellInst3_LFInst_0_LFInst_2_U9  ( .A1(
        \Red_SubCellInst3_LFInst_0_LFInst_2_n17 ), .A2(PermutationOutput3[0]), 
        .ZN(\Red_SubCellInst3_LFInst_0_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_0_LFInst_2_U8  ( .A1(PermutationOutput3[2]), 
        .A2(PermutationOutput3[1]), .ZN(
        \Red_SubCellInst3_LFInst_0_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_0_LFInst_2_U7  ( .A(
        \Red_SubCellInst3_LFInst_0_LFInst_2_n16 ), .B(
        \Red_SubCellInst3_LFInst_0_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst3_LFInst_0_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_0_LFInst_2_U6  ( .A1(PermutationOutput3[3]), 
        .A2(\Red_SubCellInst3_LFInst_0_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst3_LFInst_0_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst3_LFInst_0_LFInst_2_U5  ( .A(PermutationOutput3[1]), 
        .ZN(\Red_SubCellInst3_LFInst_0_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_0_LFInst_2_U4  ( .A1(PermutationOutput3[2]), .A2(\Red_SubCellInst3_LFInst_0_LFInst_2_n13 ), .ZN(
        \Red_SubCellInst3_LFInst_0_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst3_LFInst_0_LFInst_2_U3  ( .A(PermutationOutput3[0]), 
        .ZN(\Red_SubCellInst3_LFInst_0_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_0_LFInst_3_U6  ( .A(PermutationOutput3[1]), 
        .B(\Red_SubCellInst3_LFInst_0_LFInst_3_n8 ), .ZN(Red_Feedback3[3]) );
  NOR2_X1 \Red_SubCellInst3_LFInst_0_LFInst_3_U5  ( .A1(
        \Red_SubCellInst3_LFInst_0_LFInst_3_n7 ), .A2(
        \Red_SubCellInst3_LFInst_0_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst3_LFInst_0_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_0_LFInst_3_U4  ( .A1(PermutationOutput3[2]), 
        .A2(PermutationOutput3[3]), .ZN(
        \Red_SubCellInst3_LFInst_0_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst3_LFInst_0_LFInst_3_U3  ( .A1(PermutationOutput3[3]), 
        .A2(PermutationOutput3[0]), .ZN(
        \Red_SubCellInst3_LFInst_0_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_1_LFInst_0_U10  ( .A1(
        \Red_SubCellInst3_LFInst_1_LFInst_0_n14 ), .A2(
        \Red_SubCellInst3_LFInst_1_LFInst_0_n13 ), .ZN(Red_Feedback3[4]) );
  NAND2_X1 \Red_SubCellInst3_LFInst_1_LFInst_0_U9  ( .A1(PermutationOutput3[4]), .A2(\Red_SubCellInst3_LFInst_1_LFInst_0_n12 ), .ZN(
        \Red_SubCellInst3_LFInst_1_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_1_LFInst_0_U8  ( .A1(
        \Red_SubCellInst3_LFInst_1_LFInst_0_n11 ), .A2(PermutationOutput3[6]), 
        .ZN(\Red_SubCellInst3_LFInst_1_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_1_LFInst_0_U7  ( .A(
        \Red_SubCellInst3_LFInst_1_LFInst_0_n10 ), .B(
        \Red_SubCellInst3_LFInst_1_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst3_LFInst_1_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_1_LFInst_0_U6  ( .A1(PermutationOutput3[7]), .A2(\Red_SubCellInst3_LFInst_1_LFInst_0_n11 ), .ZN(
        \Red_SubCellInst3_LFInst_1_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst3_LFInst_1_LFInst_0_U5  ( .A(PermutationOutput3[5]), 
        .ZN(\Red_SubCellInst3_LFInst_1_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_1_LFInst_0_U4  ( .A1(PermutationOutput3[6]), .A2(\Red_SubCellInst3_LFInst_1_LFInst_0_n8 ), .ZN(
        \Red_SubCellInst3_LFInst_1_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst3_LFInst_1_LFInst_0_U3  ( .A(PermutationOutput3[4]), 
        .ZN(\Red_SubCellInst3_LFInst_1_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_1_LFInst_1_U8  ( .A1(
        \Red_SubCellInst3_LFInst_1_LFInst_1_n15 ), .A2(
        \Red_SubCellInst3_LFInst_1_LFInst_1_n14 ), .ZN(Red_Feedback3[5]) );
  NAND2_X1 \Red_SubCellInst3_LFInst_1_LFInst_1_U7  ( .A1(
        \Red_SubCellInst3_LFInst_1_LFInst_1_n13 ), .A2(PermutationOutput3[5]), 
        .ZN(\Red_SubCellInst3_LFInst_1_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_1_LFInst_1_U6  ( .A1(
        \Red_SubCellInst3_LFInst_1_LFInst_1_n12 ), .A2(PermutationOutput3[4]), 
        .ZN(\Red_SubCellInst3_LFInst_1_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_1_LFInst_1_U5  ( .A1(PermutationOutput3[7]), .A2(PermutationOutput3[6]), .ZN(\Red_SubCellInst3_LFInst_1_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst3_LFInst_1_LFInst_1_U4  ( .A1(PermutationOutput3[6]), 
        .A2(\Red_SubCellInst3_LFInst_1_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst3_LFInst_1_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_1_LFInst_1_U3  ( .A(PermutationOutput3[4]), 
        .B(PermutationOutput3[7]), .ZN(
        \Red_SubCellInst3_LFInst_1_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_1_LFInst_2_U10  ( .A1(
        \Red_SubCellInst3_LFInst_1_LFInst_2_n19 ), .A2(
        \Red_SubCellInst3_LFInst_1_LFInst_2_n18 ), .ZN(Red_Feedback3[6]) );
  AND2_X1 \Red_SubCellInst3_LFInst_1_LFInst_2_U9  ( .A1(
        \Red_SubCellInst3_LFInst_1_LFInst_2_n17 ), .A2(PermutationOutput3[4]), 
        .ZN(\Red_SubCellInst3_LFInst_1_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_1_LFInst_2_U8  ( .A1(PermutationOutput3[6]), 
        .A2(PermutationOutput3[5]), .ZN(
        \Red_SubCellInst3_LFInst_1_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_1_LFInst_2_U7  ( .A(
        \Red_SubCellInst3_LFInst_1_LFInst_2_n16 ), .B(
        \Red_SubCellInst3_LFInst_1_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst3_LFInst_1_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_1_LFInst_2_U6  ( .A1(PermutationOutput3[7]), 
        .A2(\Red_SubCellInst3_LFInst_1_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst3_LFInst_1_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst3_LFInst_1_LFInst_2_U5  ( .A(PermutationOutput3[5]), 
        .ZN(\Red_SubCellInst3_LFInst_1_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_1_LFInst_2_U4  ( .A1(PermutationOutput3[6]), .A2(\Red_SubCellInst3_LFInst_1_LFInst_2_n13 ), .ZN(
        \Red_SubCellInst3_LFInst_1_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst3_LFInst_1_LFInst_2_U3  ( .A(PermutationOutput3[4]), 
        .ZN(\Red_SubCellInst3_LFInst_1_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_1_LFInst_3_U6  ( .A(PermutationOutput3[5]), 
        .B(\Red_SubCellInst3_LFInst_1_LFInst_3_n8 ), .ZN(Red_Feedback3[7]) );
  NOR2_X1 \Red_SubCellInst3_LFInst_1_LFInst_3_U5  ( .A1(
        \Red_SubCellInst3_LFInst_1_LFInst_3_n7 ), .A2(
        \Red_SubCellInst3_LFInst_1_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst3_LFInst_1_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_1_LFInst_3_U4  ( .A1(PermutationOutput3[6]), 
        .A2(PermutationOutput3[7]), .ZN(
        \Red_SubCellInst3_LFInst_1_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst3_LFInst_1_LFInst_3_U3  ( .A1(PermutationOutput3[7]), 
        .A2(PermutationOutput3[4]), .ZN(
        \Red_SubCellInst3_LFInst_1_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_2_LFInst_0_U10  ( .A1(
        \Red_SubCellInst3_LFInst_2_LFInst_0_n14 ), .A2(
        \Red_SubCellInst3_LFInst_2_LFInst_0_n13 ), .ZN(Red_Feedback3[8]) );
  NAND2_X1 \Red_SubCellInst3_LFInst_2_LFInst_0_U9  ( .A1(PermutationOutput3[8]), .A2(\Red_SubCellInst3_LFInst_2_LFInst_0_n12 ), .ZN(
        \Red_SubCellInst3_LFInst_2_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_2_LFInst_0_U8  ( .A1(
        \Red_SubCellInst3_LFInst_2_LFInst_0_n11 ), .A2(PermutationOutput3[10]), 
        .ZN(\Red_SubCellInst3_LFInst_2_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_2_LFInst_0_U7  ( .A(
        \Red_SubCellInst3_LFInst_2_LFInst_0_n10 ), .B(
        \Red_SubCellInst3_LFInst_2_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst3_LFInst_2_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_2_LFInst_0_U6  ( .A1(
        PermutationOutput3[11]), .A2(\Red_SubCellInst3_LFInst_2_LFInst_0_n11 ), 
        .ZN(\Red_SubCellInst3_LFInst_2_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst3_LFInst_2_LFInst_0_U5  ( .A(PermutationOutput3[9]), 
        .ZN(\Red_SubCellInst3_LFInst_2_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_2_LFInst_0_U4  ( .A1(
        PermutationOutput3[10]), .A2(\Red_SubCellInst3_LFInst_2_LFInst_0_n8 ), 
        .ZN(\Red_SubCellInst3_LFInst_2_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst3_LFInst_2_LFInst_0_U3  ( .A(PermutationOutput3[8]), 
        .ZN(\Red_SubCellInst3_LFInst_2_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_2_LFInst_1_U8  ( .A1(
        \Red_SubCellInst3_LFInst_2_LFInst_1_n15 ), .A2(
        \Red_SubCellInst3_LFInst_2_LFInst_1_n14 ), .ZN(Red_Feedback3[9]) );
  NAND2_X1 \Red_SubCellInst3_LFInst_2_LFInst_1_U7  ( .A1(
        \Red_SubCellInst3_LFInst_2_LFInst_1_n13 ), .A2(PermutationOutput3[9]), 
        .ZN(\Red_SubCellInst3_LFInst_2_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_2_LFInst_1_U6  ( .A1(
        \Red_SubCellInst3_LFInst_2_LFInst_1_n12 ), .A2(PermutationOutput3[8]), 
        .ZN(\Red_SubCellInst3_LFInst_2_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_2_LFInst_1_U5  ( .A1(
        PermutationOutput3[11]), .A2(PermutationOutput3[10]), .ZN(
        \Red_SubCellInst3_LFInst_2_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst3_LFInst_2_LFInst_1_U4  ( .A1(PermutationOutput3[10]), 
        .A2(\Red_SubCellInst3_LFInst_2_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst3_LFInst_2_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_2_LFInst_1_U3  ( .A(PermutationOutput3[8]), 
        .B(PermutationOutput3[11]), .ZN(
        \Red_SubCellInst3_LFInst_2_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_2_LFInst_2_U10  ( .A1(
        \Red_SubCellInst3_LFInst_2_LFInst_2_n19 ), .A2(
        \Red_SubCellInst3_LFInst_2_LFInst_2_n18 ), .ZN(Red_Feedback3[10]) );
  AND2_X1 \Red_SubCellInst3_LFInst_2_LFInst_2_U9  ( .A1(
        \Red_SubCellInst3_LFInst_2_LFInst_2_n17 ), .A2(PermutationOutput3[8]), 
        .ZN(\Red_SubCellInst3_LFInst_2_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_2_LFInst_2_U8  ( .A1(PermutationOutput3[10]), .A2(PermutationOutput3[9]), .ZN(\Red_SubCellInst3_LFInst_2_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_2_LFInst_2_U7  ( .A(
        \Red_SubCellInst3_LFInst_2_LFInst_2_n16 ), .B(
        \Red_SubCellInst3_LFInst_2_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst3_LFInst_2_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_2_LFInst_2_U6  ( .A1(PermutationOutput3[11]), .A2(\Red_SubCellInst3_LFInst_2_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst3_LFInst_2_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst3_LFInst_2_LFInst_2_U5  ( .A(PermutationOutput3[9]), 
        .ZN(\Red_SubCellInst3_LFInst_2_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_2_LFInst_2_U4  ( .A1(
        PermutationOutput3[10]), .A2(\Red_SubCellInst3_LFInst_2_LFInst_2_n13 ), 
        .ZN(\Red_SubCellInst3_LFInst_2_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst3_LFInst_2_LFInst_2_U3  ( .A(PermutationOutput3[8]), 
        .ZN(\Red_SubCellInst3_LFInst_2_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_2_LFInst_3_U6  ( .A(PermutationOutput3[9]), 
        .B(\Red_SubCellInst3_LFInst_2_LFInst_3_n8 ), .ZN(Red_Feedback3[11]) );
  NOR2_X1 \Red_SubCellInst3_LFInst_2_LFInst_3_U5  ( .A1(
        \Red_SubCellInst3_LFInst_2_LFInst_3_n7 ), .A2(
        \Red_SubCellInst3_LFInst_2_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst3_LFInst_2_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_2_LFInst_3_U4  ( .A1(PermutationOutput3[10]), .A2(PermutationOutput3[11]), .ZN(\Red_SubCellInst3_LFInst_2_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst3_LFInst_2_LFInst_3_U3  ( .A1(PermutationOutput3[11]), .A2(PermutationOutput3[8]), .ZN(\Red_SubCellInst3_LFInst_2_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_3_LFInst_0_U10  ( .A1(
        \Red_SubCellInst3_LFInst_3_LFInst_0_n14 ), .A2(
        \Red_SubCellInst3_LFInst_3_LFInst_0_n13 ), .ZN(Red_Feedback3[12]) );
  NAND2_X1 \Red_SubCellInst3_LFInst_3_LFInst_0_U9  ( .A1(
        PermutationOutput3[12]), .A2(\Red_SubCellInst3_LFInst_3_LFInst_0_n12 ), 
        .ZN(\Red_SubCellInst3_LFInst_3_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_3_LFInst_0_U8  ( .A1(
        \Red_SubCellInst3_LFInst_3_LFInst_0_n11 ), .A2(PermutationOutput3[14]), 
        .ZN(\Red_SubCellInst3_LFInst_3_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_3_LFInst_0_U7  ( .A(
        \Red_SubCellInst3_LFInst_3_LFInst_0_n10 ), .B(
        \Red_SubCellInst3_LFInst_3_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst3_LFInst_3_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_3_LFInst_0_U6  ( .A1(
        PermutationOutput3[15]), .A2(\Red_SubCellInst3_LFInst_3_LFInst_0_n11 ), 
        .ZN(\Red_SubCellInst3_LFInst_3_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst3_LFInst_3_LFInst_0_U5  ( .A(PermutationOutput3[13]), 
        .ZN(\Red_SubCellInst3_LFInst_3_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_3_LFInst_0_U4  ( .A1(
        PermutationOutput3[14]), .A2(\Red_SubCellInst3_LFInst_3_LFInst_0_n8 ), 
        .ZN(\Red_SubCellInst3_LFInst_3_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst3_LFInst_3_LFInst_0_U3  ( .A(PermutationOutput3[12]), 
        .ZN(\Red_SubCellInst3_LFInst_3_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_3_LFInst_1_U8  ( .A1(
        \Red_SubCellInst3_LFInst_3_LFInst_1_n15 ), .A2(
        \Red_SubCellInst3_LFInst_3_LFInst_1_n14 ), .ZN(Red_Feedback3[13]) );
  NAND2_X1 \Red_SubCellInst3_LFInst_3_LFInst_1_U7  ( .A1(
        \Red_SubCellInst3_LFInst_3_LFInst_1_n13 ), .A2(PermutationOutput3[13]), 
        .ZN(\Red_SubCellInst3_LFInst_3_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_3_LFInst_1_U6  ( .A1(
        \Red_SubCellInst3_LFInst_3_LFInst_1_n12 ), .A2(PermutationOutput3[12]), 
        .ZN(\Red_SubCellInst3_LFInst_3_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_3_LFInst_1_U5  ( .A1(
        PermutationOutput3[15]), .A2(PermutationOutput3[14]), .ZN(
        \Red_SubCellInst3_LFInst_3_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst3_LFInst_3_LFInst_1_U4  ( .A1(PermutationOutput3[14]), 
        .A2(\Red_SubCellInst3_LFInst_3_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst3_LFInst_3_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_3_LFInst_1_U3  ( .A(PermutationOutput3[12]), .B(PermutationOutput3[15]), .ZN(\Red_SubCellInst3_LFInst_3_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_3_LFInst_2_U10  ( .A1(
        \Red_SubCellInst3_LFInst_3_LFInst_2_n19 ), .A2(
        \Red_SubCellInst3_LFInst_3_LFInst_2_n18 ), .ZN(Red_Feedback3[14]) );
  AND2_X1 \Red_SubCellInst3_LFInst_3_LFInst_2_U9  ( .A1(
        \Red_SubCellInst3_LFInst_3_LFInst_2_n17 ), .A2(PermutationOutput3[12]), 
        .ZN(\Red_SubCellInst3_LFInst_3_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_3_LFInst_2_U8  ( .A1(PermutationOutput3[14]), .A2(PermutationOutput3[13]), .ZN(\Red_SubCellInst3_LFInst_3_LFInst_2_n17 )
         );
  XNOR2_X1 \Red_SubCellInst3_LFInst_3_LFInst_2_U7  ( .A(
        \Red_SubCellInst3_LFInst_3_LFInst_2_n16 ), .B(
        \Red_SubCellInst3_LFInst_3_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst3_LFInst_3_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_3_LFInst_2_U6  ( .A1(PermutationOutput3[15]), .A2(\Red_SubCellInst3_LFInst_3_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst3_LFInst_3_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst3_LFInst_3_LFInst_2_U5  ( .A(PermutationOutput3[13]), 
        .ZN(\Red_SubCellInst3_LFInst_3_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_3_LFInst_2_U4  ( .A1(
        PermutationOutput3[14]), .A2(\Red_SubCellInst3_LFInst_3_LFInst_2_n13 ), 
        .ZN(\Red_SubCellInst3_LFInst_3_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst3_LFInst_3_LFInst_2_U3  ( .A(PermutationOutput3[12]), 
        .ZN(\Red_SubCellInst3_LFInst_3_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_3_LFInst_3_U6  ( .A(PermutationOutput3[13]), .B(\Red_SubCellInst3_LFInst_3_LFInst_3_n8 ), .ZN(Red_Feedback3[15]) );
  NOR2_X1 \Red_SubCellInst3_LFInst_3_LFInst_3_U5  ( .A1(
        \Red_SubCellInst3_LFInst_3_LFInst_3_n7 ), .A2(
        \Red_SubCellInst3_LFInst_3_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst3_LFInst_3_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_3_LFInst_3_U4  ( .A1(PermutationOutput3[14]), .A2(PermutationOutput3[15]), .ZN(\Red_SubCellInst3_LFInst_3_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst3_LFInst_3_LFInst_3_U3  ( .A1(PermutationOutput3[15]), .A2(PermutationOutput3[12]), .ZN(\Red_SubCellInst3_LFInst_3_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_4_LFInst_0_U10  ( .A1(
        \Red_SubCellInst3_LFInst_4_LFInst_0_n14 ), .A2(
        \Red_SubCellInst3_LFInst_4_LFInst_0_n13 ), .ZN(Red_Feedback3[16]) );
  NAND2_X1 \Red_SubCellInst3_LFInst_4_LFInst_0_U9  ( .A1(
        PermutationOutput3[16]), .A2(\Red_SubCellInst3_LFInst_4_LFInst_0_n12 ), 
        .ZN(\Red_SubCellInst3_LFInst_4_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_4_LFInst_0_U8  ( .A1(
        \Red_SubCellInst3_LFInst_4_LFInst_0_n11 ), .A2(PermutationOutput3[18]), 
        .ZN(\Red_SubCellInst3_LFInst_4_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_4_LFInst_0_U7  ( .A(
        \Red_SubCellInst3_LFInst_4_LFInst_0_n10 ), .B(
        \Red_SubCellInst3_LFInst_4_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst3_LFInst_4_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_4_LFInst_0_U6  ( .A1(
        PermutationOutput3[19]), .A2(\Red_SubCellInst3_LFInst_4_LFInst_0_n11 ), 
        .ZN(\Red_SubCellInst3_LFInst_4_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst3_LFInst_4_LFInst_0_U5  ( .A(PermutationOutput3[17]), 
        .ZN(\Red_SubCellInst3_LFInst_4_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_4_LFInst_0_U4  ( .A1(
        PermutationOutput3[18]), .A2(\Red_SubCellInst3_LFInst_4_LFInst_0_n8 ), 
        .ZN(\Red_SubCellInst3_LFInst_4_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst3_LFInst_4_LFInst_0_U3  ( .A(PermutationOutput3[16]), 
        .ZN(\Red_SubCellInst3_LFInst_4_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_4_LFInst_1_U8  ( .A1(
        \Red_SubCellInst3_LFInst_4_LFInst_1_n15 ), .A2(
        \Red_SubCellInst3_LFInst_4_LFInst_1_n14 ), .ZN(Red_Feedback3[17]) );
  NAND2_X1 \Red_SubCellInst3_LFInst_4_LFInst_1_U7  ( .A1(
        \Red_SubCellInst3_LFInst_4_LFInst_1_n13 ), .A2(PermutationOutput3[17]), 
        .ZN(\Red_SubCellInst3_LFInst_4_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_4_LFInst_1_U6  ( .A1(
        \Red_SubCellInst3_LFInst_4_LFInst_1_n12 ), .A2(PermutationOutput3[16]), 
        .ZN(\Red_SubCellInst3_LFInst_4_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_4_LFInst_1_U5  ( .A1(
        PermutationOutput3[19]), .A2(PermutationOutput3[18]), .ZN(
        \Red_SubCellInst3_LFInst_4_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst3_LFInst_4_LFInst_1_U4  ( .A1(PermutationOutput3[18]), 
        .A2(\Red_SubCellInst3_LFInst_4_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst3_LFInst_4_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_4_LFInst_1_U3  ( .A(PermutationOutput3[16]), .B(PermutationOutput3[19]), .ZN(\Red_SubCellInst3_LFInst_4_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_4_LFInst_2_U10  ( .A1(
        \Red_SubCellInst3_LFInst_4_LFInst_2_n19 ), .A2(
        \Red_SubCellInst3_LFInst_4_LFInst_2_n18 ), .ZN(Red_Feedback3[18]) );
  AND2_X1 \Red_SubCellInst3_LFInst_4_LFInst_2_U9  ( .A1(
        \Red_SubCellInst3_LFInst_4_LFInst_2_n17 ), .A2(PermutationOutput3[16]), 
        .ZN(\Red_SubCellInst3_LFInst_4_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_4_LFInst_2_U8  ( .A1(PermutationOutput3[18]), .A2(PermutationOutput3[17]), .ZN(\Red_SubCellInst3_LFInst_4_LFInst_2_n17 )
         );
  XNOR2_X1 \Red_SubCellInst3_LFInst_4_LFInst_2_U7  ( .A(
        \Red_SubCellInst3_LFInst_4_LFInst_2_n16 ), .B(
        \Red_SubCellInst3_LFInst_4_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst3_LFInst_4_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_4_LFInst_2_U6  ( .A1(PermutationOutput3[19]), .A2(\Red_SubCellInst3_LFInst_4_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst3_LFInst_4_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst3_LFInst_4_LFInst_2_U5  ( .A(PermutationOutput3[17]), 
        .ZN(\Red_SubCellInst3_LFInst_4_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_4_LFInst_2_U4  ( .A1(
        PermutationOutput3[18]), .A2(\Red_SubCellInst3_LFInst_4_LFInst_2_n13 ), 
        .ZN(\Red_SubCellInst3_LFInst_4_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst3_LFInst_4_LFInst_2_U3  ( .A(PermutationOutput3[16]), 
        .ZN(\Red_SubCellInst3_LFInst_4_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_4_LFInst_3_U6  ( .A(PermutationOutput3[17]), .B(\Red_SubCellInst3_LFInst_4_LFInst_3_n8 ), .ZN(Red_Feedback3[19]) );
  NOR2_X1 \Red_SubCellInst3_LFInst_4_LFInst_3_U5  ( .A1(
        \Red_SubCellInst3_LFInst_4_LFInst_3_n7 ), .A2(
        \Red_SubCellInst3_LFInst_4_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst3_LFInst_4_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_4_LFInst_3_U4  ( .A1(PermutationOutput3[18]), .A2(PermutationOutput3[19]), .ZN(\Red_SubCellInst3_LFInst_4_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst3_LFInst_4_LFInst_3_U3  ( .A1(PermutationOutput3[19]), .A2(PermutationOutput3[16]), .ZN(\Red_SubCellInst3_LFInst_4_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_5_LFInst_0_U10  ( .A1(
        \Red_SubCellInst3_LFInst_5_LFInst_0_n14 ), .A2(
        \Red_SubCellInst3_LFInst_5_LFInst_0_n13 ), .ZN(Red_Feedback3[20]) );
  NAND2_X1 \Red_SubCellInst3_LFInst_5_LFInst_0_U9  ( .A1(
        PermutationOutput3[20]), .A2(\Red_SubCellInst3_LFInst_5_LFInst_0_n12 ), 
        .ZN(\Red_SubCellInst3_LFInst_5_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_5_LFInst_0_U8  ( .A1(
        \Red_SubCellInst3_LFInst_5_LFInst_0_n11 ), .A2(PermutationOutput3[22]), 
        .ZN(\Red_SubCellInst3_LFInst_5_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_5_LFInst_0_U7  ( .A(
        \Red_SubCellInst3_LFInst_5_LFInst_0_n10 ), .B(
        \Red_SubCellInst3_LFInst_5_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst3_LFInst_5_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_5_LFInst_0_U6  ( .A1(
        PermutationOutput3[23]), .A2(\Red_SubCellInst3_LFInst_5_LFInst_0_n11 ), 
        .ZN(\Red_SubCellInst3_LFInst_5_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst3_LFInst_5_LFInst_0_U5  ( .A(PermutationOutput3[21]), 
        .ZN(\Red_SubCellInst3_LFInst_5_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_5_LFInst_0_U4  ( .A1(
        PermutationOutput3[22]), .A2(\Red_SubCellInst3_LFInst_5_LFInst_0_n8 ), 
        .ZN(\Red_SubCellInst3_LFInst_5_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst3_LFInst_5_LFInst_0_U3  ( .A(PermutationOutput3[20]), 
        .ZN(\Red_SubCellInst3_LFInst_5_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_5_LFInst_1_U8  ( .A1(
        \Red_SubCellInst3_LFInst_5_LFInst_1_n15 ), .A2(
        \Red_SubCellInst3_LFInst_5_LFInst_1_n14 ), .ZN(Red_Feedback3[21]) );
  NAND2_X1 \Red_SubCellInst3_LFInst_5_LFInst_1_U7  ( .A1(
        \Red_SubCellInst3_LFInst_5_LFInst_1_n13 ), .A2(PermutationOutput3[21]), 
        .ZN(\Red_SubCellInst3_LFInst_5_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_5_LFInst_1_U6  ( .A1(
        \Red_SubCellInst3_LFInst_5_LFInst_1_n12 ), .A2(PermutationOutput3[20]), 
        .ZN(\Red_SubCellInst3_LFInst_5_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_5_LFInst_1_U5  ( .A1(
        PermutationOutput3[23]), .A2(PermutationOutput3[22]), .ZN(
        \Red_SubCellInst3_LFInst_5_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst3_LFInst_5_LFInst_1_U4  ( .A1(PermutationOutput3[22]), 
        .A2(\Red_SubCellInst3_LFInst_5_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst3_LFInst_5_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_5_LFInst_1_U3  ( .A(PermutationOutput3[20]), .B(PermutationOutput3[23]), .ZN(\Red_SubCellInst3_LFInst_5_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_5_LFInst_2_U10  ( .A1(
        \Red_SubCellInst3_LFInst_5_LFInst_2_n19 ), .A2(
        \Red_SubCellInst3_LFInst_5_LFInst_2_n18 ), .ZN(Red_Feedback3[22]) );
  AND2_X1 \Red_SubCellInst3_LFInst_5_LFInst_2_U9  ( .A1(
        \Red_SubCellInst3_LFInst_5_LFInst_2_n17 ), .A2(PermutationOutput3[20]), 
        .ZN(\Red_SubCellInst3_LFInst_5_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_5_LFInst_2_U8  ( .A1(PermutationOutput3[22]), .A2(PermutationOutput3[21]), .ZN(\Red_SubCellInst3_LFInst_5_LFInst_2_n17 )
         );
  XNOR2_X1 \Red_SubCellInst3_LFInst_5_LFInst_2_U7  ( .A(
        \Red_SubCellInst3_LFInst_5_LFInst_2_n16 ), .B(
        \Red_SubCellInst3_LFInst_5_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst3_LFInst_5_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_5_LFInst_2_U6  ( .A1(PermutationOutput3[23]), .A2(\Red_SubCellInst3_LFInst_5_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst3_LFInst_5_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst3_LFInst_5_LFInst_2_U5  ( .A(PermutationOutput3[21]), 
        .ZN(\Red_SubCellInst3_LFInst_5_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_5_LFInst_2_U4  ( .A1(
        PermutationOutput3[22]), .A2(\Red_SubCellInst3_LFInst_5_LFInst_2_n13 ), 
        .ZN(\Red_SubCellInst3_LFInst_5_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst3_LFInst_5_LFInst_2_U3  ( .A(PermutationOutput3[20]), 
        .ZN(\Red_SubCellInst3_LFInst_5_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_5_LFInst_3_U6  ( .A(PermutationOutput3[21]), .B(\Red_SubCellInst3_LFInst_5_LFInst_3_n8 ), .ZN(Red_Feedback3[23]) );
  NOR2_X1 \Red_SubCellInst3_LFInst_5_LFInst_3_U5  ( .A1(
        \Red_SubCellInst3_LFInst_5_LFInst_3_n7 ), .A2(
        \Red_SubCellInst3_LFInst_5_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst3_LFInst_5_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_5_LFInst_3_U4  ( .A1(PermutationOutput3[22]), .A2(PermutationOutput3[23]), .ZN(\Red_SubCellInst3_LFInst_5_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst3_LFInst_5_LFInst_3_U3  ( .A1(PermutationOutput3[23]), .A2(PermutationOutput3[20]), .ZN(\Red_SubCellInst3_LFInst_5_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_6_LFInst_0_U10  ( .A1(
        \Red_SubCellInst3_LFInst_6_LFInst_0_n14 ), .A2(
        \Red_SubCellInst3_LFInst_6_LFInst_0_n13 ), .ZN(Red_Feedback3[24]) );
  NAND2_X1 \Red_SubCellInst3_LFInst_6_LFInst_0_U9  ( .A1(
        PermutationOutput3[24]), .A2(\Red_SubCellInst3_LFInst_6_LFInst_0_n12 ), 
        .ZN(\Red_SubCellInst3_LFInst_6_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_6_LFInst_0_U8  ( .A1(
        \Red_SubCellInst3_LFInst_6_LFInst_0_n11 ), .A2(PermutationOutput3[26]), 
        .ZN(\Red_SubCellInst3_LFInst_6_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_6_LFInst_0_U7  ( .A(
        \Red_SubCellInst3_LFInst_6_LFInst_0_n10 ), .B(
        \Red_SubCellInst3_LFInst_6_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst3_LFInst_6_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_6_LFInst_0_U6  ( .A1(
        PermutationOutput3[27]), .A2(\Red_SubCellInst3_LFInst_6_LFInst_0_n11 ), 
        .ZN(\Red_SubCellInst3_LFInst_6_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst3_LFInst_6_LFInst_0_U5  ( .A(PermutationOutput3[25]), 
        .ZN(\Red_SubCellInst3_LFInst_6_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_6_LFInst_0_U4  ( .A1(
        PermutationOutput3[26]), .A2(\Red_SubCellInst3_LFInst_6_LFInst_0_n8 ), 
        .ZN(\Red_SubCellInst3_LFInst_6_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst3_LFInst_6_LFInst_0_U3  ( .A(PermutationOutput3[24]), 
        .ZN(\Red_SubCellInst3_LFInst_6_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_6_LFInst_1_U8  ( .A1(
        \Red_SubCellInst3_LFInst_6_LFInst_1_n15 ), .A2(
        \Red_SubCellInst3_LFInst_6_LFInst_1_n14 ), .ZN(Red_Feedback3[25]) );
  NAND2_X1 \Red_SubCellInst3_LFInst_6_LFInst_1_U7  ( .A1(
        \Red_SubCellInst3_LFInst_6_LFInst_1_n13 ), .A2(PermutationOutput3[25]), 
        .ZN(\Red_SubCellInst3_LFInst_6_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_6_LFInst_1_U6  ( .A1(
        \Red_SubCellInst3_LFInst_6_LFInst_1_n12 ), .A2(PermutationOutput3[24]), 
        .ZN(\Red_SubCellInst3_LFInst_6_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_6_LFInst_1_U5  ( .A1(
        PermutationOutput3[27]), .A2(PermutationOutput3[26]), .ZN(
        \Red_SubCellInst3_LFInst_6_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst3_LFInst_6_LFInst_1_U4  ( .A1(PermutationOutput3[26]), 
        .A2(\Red_SubCellInst3_LFInst_6_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst3_LFInst_6_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_6_LFInst_1_U3  ( .A(PermutationOutput3[24]), .B(PermutationOutput3[27]), .ZN(\Red_SubCellInst3_LFInst_6_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_6_LFInst_2_U10  ( .A1(
        \Red_SubCellInst3_LFInst_6_LFInst_2_n19 ), .A2(
        \Red_SubCellInst3_LFInst_6_LFInst_2_n18 ), .ZN(Red_Feedback3[26]) );
  AND2_X1 \Red_SubCellInst3_LFInst_6_LFInst_2_U9  ( .A1(
        \Red_SubCellInst3_LFInst_6_LFInst_2_n17 ), .A2(PermutationOutput3[24]), 
        .ZN(\Red_SubCellInst3_LFInst_6_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_6_LFInst_2_U8  ( .A1(PermutationOutput3[26]), .A2(PermutationOutput3[25]), .ZN(\Red_SubCellInst3_LFInst_6_LFInst_2_n17 )
         );
  XNOR2_X1 \Red_SubCellInst3_LFInst_6_LFInst_2_U7  ( .A(
        \Red_SubCellInst3_LFInst_6_LFInst_2_n16 ), .B(
        \Red_SubCellInst3_LFInst_6_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst3_LFInst_6_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_6_LFInst_2_U6  ( .A1(PermutationOutput3[27]), .A2(\Red_SubCellInst3_LFInst_6_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst3_LFInst_6_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst3_LFInst_6_LFInst_2_U5  ( .A(PermutationOutput3[25]), 
        .ZN(\Red_SubCellInst3_LFInst_6_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_6_LFInst_2_U4  ( .A1(
        PermutationOutput3[26]), .A2(\Red_SubCellInst3_LFInst_6_LFInst_2_n13 ), 
        .ZN(\Red_SubCellInst3_LFInst_6_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst3_LFInst_6_LFInst_2_U3  ( .A(PermutationOutput3[24]), 
        .ZN(\Red_SubCellInst3_LFInst_6_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_6_LFInst_3_U6  ( .A(PermutationOutput3[25]), .B(\Red_SubCellInst3_LFInst_6_LFInst_3_n8 ), .ZN(Red_Feedback3[27]) );
  NOR2_X1 \Red_SubCellInst3_LFInst_6_LFInst_3_U5  ( .A1(
        \Red_SubCellInst3_LFInst_6_LFInst_3_n7 ), .A2(
        \Red_SubCellInst3_LFInst_6_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst3_LFInst_6_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_6_LFInst_3_U4  ( .A1(PermutationOutput3[26]), .A2(PermutationOutput3[27]), .ZN(\Red_SubCellInst3_LFInst_6_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst3_LFInst_6_LFInst_3_U3  ( .A1(PermutationOutput3[27]), .A2(PermutationOutput3[24]), .ZN(\Red_SubCellInst3_LFInst_6_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_7_LFInst_0_U10  ( .A1(
        \Red_SubCellInst3_LFInst_7_LFInst_0_n14 ), .A2(
        \Red_SubCellInst3_LFInst_7_LFInst_0_n13 ), .ZN(Red_Feedback3[28]) );
  NAND2_X1 \Red_SubCellInst3_LFInst_7_LFInst_0_U9  ( .A1(
        PermutationOutput3[28]), .A2(\Red_SubCellInst3_LFInst_7_LFInst_0_n12 ), 
        .ZN(\Red_SubCellInst3_LFInst_7_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_7_LFInst_0_U8  ( .A1(
        \Red_SubCellInst3_LFInst_7_LFInst_0_n11 ), .A2(PermutationOutput3[30]), 
        .ZN(\Red_SubCellInst3_LFInst_7_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_7_LFInst_0_U7  ( .A(
        \Red_SubCellInst3_LFInst_7_LFInst_0_n10 ), .B(
        \Red_SubCellInst3_LFInst_7_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst3_LFInst_7_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_7_LFInst_0_U6  ( .A1(
        PermutationOutput3[31]), .A2(\Red_SubCellInst3_LFInst_7_LFInst_0_n11 ), 
        .ZN(\Red_SubCellInst3_LFInst_7_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst3_LFInst_7_LFInst_0_U5  ( .A(PermutationOutput3[29]), 
        .ZN(\Red_SubCellInst3_LFInst_7_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_7_LFInst_0_U4  ( .A1(
        PermutationOutput3[30]), .A2(\Red_SubCellInst3_LFInst_7_LFInst_0_n8 ), 
        .ZN(\Red_SubCellInst3_LFInst_7_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst3_LFInst_7_LFInst_0_U3  ( .A(PermutationOutput3[28]), 
        .ZN(\Red_SubCellInst3_LFInst_7_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_7_LFInst_1_U8  ( .A1(
        \Red_SubCellInst3_LFInst_7_LFInst_1_n15 ), .A2(
        \Red_SubCellInst3_LFInst_7_LFInst_1_n14 ), .ZN(Red_Feedback3[29]) );
  NAND2_X1 \Red_SubCellInst3_LFInst_7_LFInst_1_U7  ( .A1(
        \Red_SubCellInst3_LFInst_7_LFInst_1_n13 ), .A2(PermutationOutput3[29]), 
        .ZN(\Red_SubCellInst3_LFInst_7_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_7_LFInst_1_U6  ( .A1(
        \Red_SubCellInst3_LFInst_7_LFInst_1_n12 ), .A2(PermutationOutput3[28]), 
        .ZN(\Red_SubCellInst3_LFInst_7_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_7_LFInst_1_U5  ( .A1(
        PermutationOutput3[31]), .A2(PermutationOutput3[30]), .ZN(
        \Red_SubCellInst3_LFInst_7_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst3_LFInst_7_LFInst_1_U4  ( .A1(PermutationOutput3[30]), 
        .A2(\Red_SubCellInst3_LFInst_7_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst3_LFInst_7_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_7_LFInst_1_U3  ( .A(PermutationOutput3[28]), .B(PermutationOutput3[31]), .ZN(\Red_SubCellInst3_LFInst_7_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_7_LFInst_2_U10  ( .A1(
        \Red_SubCellInst3_LFInst_7_LFInst_2_n19 ), .A2(
        \Red_SubCellInst3_LFInst_7_LFInst_2_n18 ), .ZN(Red_Feedback3[30]) );
  AND2_X1 \Red_SubCellInst3_LFInst_7_LFInst_2_U9  ( .A1(
        \Red_SubCellInst3_LFInst_7_LFInst_2_n17 ), .A2(PermutationOutput3[28]), 
        .ZN(\Red_SubCellInst3_LFInst_7_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_7_LFInst_2_U8  ( .A1(PermutationOutput3[30]), .A2(PermutationOutput3[29]), .ZN(\Red_SubCellInst3_LFInst_7_LFInst_2_n17 )
         );
  XNOR2_X1 \Red_SubCellInst3_LFInst_7_LFInst_2_U7  ( .A(
        \Red_SubCellInst3_LFInst_7_LFInst_2_n16 ), .B(
        \Red_SubCellInst3_LFInst_7_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst3_LFInst_7_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_7_LFInst_2_U6  ( .A1(PermutationOutput3[31]), .A2(\Red_SubCellInst3_LFInst_7_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst3_LFInst_7_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst3_LFInst_7_LFInst_2_U5  ( .A(PermutationOutput3[29]), 
        .ZN(\Red_SubCellInst3_LFInst_7_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_7_LFInst_2_U4  ( .A1(
        PermutationOutput3[30]), .A2(\Red_SubCellInst3_LFInst_7_LFInst_2_n13 ), 
        .ZN(\Red_SubCellInst3_LFInst_7_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst3_LFInst_7_LFInst_2_U3  ( .A(PermutationOutput3[28]), 
        .ZN(\Red_SubCellInst3_LFInst_7_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_7_LFInst_3_U6  ( .A(PermutationOutput3[29]), .B(\Red_SubCellInst3_LFInst_7_LFInst_3_n8 ), .ZN(Red_Feedback3[31]) );
  NOR2_X1 \Red_SubCellInst3_LFInst_7_LFInst_3_U5  ( .A1(
        \Red_SubCellInst3_LFInst_7_LFInst_3_n7 ), .A2(
        \Red_SubCellInst3_LFInst_7_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst3_LFInst_7_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_7_LFInst_3_U4  ( .A1(PermutationOutput3[30]), .A2(PermutationOutput3[31]), .ZN(\Red_SubCellInst3_LFInst_7_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst3_LFInst_7_LFInst_3_U3  ( .A1(PermutationOutput3[31]), .A2(PermutationOutput3[28]), .ZN(\Red_SubCellInst3_LFInst_7_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_8_LFInst_0_U10  ( .A1(
        \Red_SubCellInst3_LFInst_8_LFInst_0_n14 ), .A2(
        \Red_SubCellInst3_LFInst_8_LFInst_0_n13 ), .ZN(Red_Feedback3[32]) );
  NAND2_X1 \Red_SubCellInst3_LFInst_8_LFInst_0_U9  ( .A1(
        PermutationOutput3[32]), .A2(\Red_SubCellInst3_LFInst_8_LFInst_0_n12 ), 
        .ZN(\Red_SubCellInst3_LFInst_8_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_8_LFInst_0_U8  ( .A1(
        \Red_SubCellInst3_LFInst_8_LFInst_0_n11 ), .A2(PermutationOutput3[34]), 
        .ZN(\Red_SubCellInst3_LFInst_8_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_8_LFInst_0_U7  ( .A(
        \Red_SubCellInst3_LFInst_8_LFInst_0_n10 ), .B(
        \Red_SubCellInst3_LFInst_8_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst3_LFInst_8_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_8_LFInst_0_U6  ( .A1(
        PermutationOutput3[35]), .A2(\Red_SubCellInst3_LFInst_8_LFInst_0_n11 ), 
        .ZN(\Red_SubCellInst3_LFInst_8_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst3_LFInst_8_LFInst_0_U5  ( .A(PermutationOutput3[33]), 
        .ZN(\Red_SubCellInst3_LFInst_8_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_8_LFInst_0_U4  ( .A1(
        PermutationOutput3[34]), .A2(\Red_SubCellInst3_LFInst_8_LFInst_0_n8 ), 
        .ZN(\Red_SubCellInst3_LFInst_8_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst3_LFInst_8_LFInst_0_U3  ( .A(PermutationOutput3[32]), 
        .ZN(\Red_SubCellInst3_LFInst_8_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_8_LFInst_1_U8  ( .A1(
        \Red_SubCellInst3_LFInst_8_LFInst_1_n15 ), .A2(
        \Red_SubCellInst3_LFInst_8_LFInst_1_n14 ), .ZN(Red_Feedback3[33]) );
  NAND2_X1 \Red_SubCellInst3_LFInst_8_LFInst_1_U7  ( .A1(
        \Red_SubCellInst3_LFInst_8_LFInst_1_n13 ), .A2(PermutationOutput3[33]), 
        .ZN(\Red_SubCellInst3_LFInst_8_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_8_LFInst_1_U6  ( .A1(
        \Red_SubCellInst3_LFInst_8_LFInst_1_n12 ), .A2(PermutationOutput3[32]), 
        .ZN(\Red_SubCellInst3_LFInst_8_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_8_LFInst_1_U5  ( .A1(
        PermutationOutput3[35]), .A2(PermutationOutput3[34]), .ZN(
        \Red_SubCellInst3_LFInst_8_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst3_LFInst_8_LFInst_1_U4  ( .A1(PermutationOutput3[34]), 
        .A2(\Red_SubCellInst3_LFInst_8_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst3_LFInst_8_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_8_LFInst_1_U3  ( .A(PermutationOutput3[32]), .B(PermutationOutput3[35]), .ZN(\Red_SubCellInst3_LFInst_8_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_8_LFInst_2_U10  ( .A1(
        \Red_SubCellInst3_LFInst_8_LFInst_2_n19 ), .A2(
        \Red_SubCellInst3_LFInst_8_LFInst_2_n18 ), .ZN(Red_Feedback3[34]) );
  AND2_X1 \Red_SubCellInst3_LFInst_8_LFInst_2_U9  ( .A1(
        \Red_SubCellInst3_LFInst_8_LFInst_2_n17 ), .A2(PermutationOutput3[32]), 
        .ZN(\Red_SubCellInst3_LFInst_8_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_8_LFInst_2_U8  ( .A1(PermutationOutput3[34]), .A2(PermutationOutput3[33]), .ZN(\Red_SubCellInst3_LFInst_8_LFInst_2_n17 )
         );
  XNOR2_X1 \Red_SubCellInst3_LFInst_8_LFInst_2_U7  ( .A(
        \Red_SubCellInst3_LFInst_8_LFInst_2_n16 ), .B(
        \Red_SubCellInst3_LFInst_8_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst3_LFInst_8_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_8_LFInst_2_U6  ( .A1(PermutationOutput3[35]), .A2(\Red_SubCellInst3_LFInst_8_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst3_LFInst_8_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst3_LFInst_8_LFInst_2_U5  ( .A(PermutationOutput3[33]), 
        .ZN(\Red_SubCellInst3_LFInst_8_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_8_LFInst_2_U4  ( .A1(
        PermutationOutput3[34]), .A2(\Red_SubCellInst3_LFInst_8_LFInst_2_n13 ), 
        .ZN(\Red_SubCellInst3_LFInst_8_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst3_LFInst_8_LFInst_2_U3  ( .A(PermutationOutput3[32]), 
        .ZN(\Red_SubCellInst3_LFInst_8_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_8_LFInst_3_U6  ( .A(PermutationOutput3[33]), .B(\Red_SubCellInst3_LFInst_8_LFInst_3_n8 ), .ZN(Red_Feedback3[35]) );
  NOR2_X1 \Red_SubCellInst3_LFInst_8_LFInst_3_U5  ( .A1(
        \Red_SubCellInst3_LFInst_8_LFInst_3_n7 ), .A2(
        \Red_SubCellInst3_LFInst_8_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst3_LFInst_8_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_8_LFInst_3_U4  ( .A1(PermutationOutput3[34]), .A2(PermutationOutput3[35]), .ZN(\Red_SubCellInst3_LFInst_8_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst3_LFInst_8_LFInst_3_U3  ( .A1(PermutationOutput3[35]), .A2(PermutationOutput3[32]), .ZN(\Red_SubCellInst3_LFInst_8_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_9_LFInst_0_U10  ( .A1(
        \Red_SubCellInst3_LFInst_9_LFInst_0_n14 ), .A2(
        \Red_SubCellInst3_LFInst_9_LFInst_0_n13 ), .ZN(Red_Feedback3[36]) );
  NAND2_X1 \Red_SubCellInst3_LFInst_9_LFInst_0_U9  ( .A1(
        PermutationOutput3[36]), .A2(\Red_SubCellInst3_LFInst_9_LFInst_0_n12 ), 
        .ZN(\Red_SubCellInst3_LFInst_9_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_9_LFInst_0_U8  ( .A1(
        \Red_SubCellInst3_LFInst_9_LFInst_0_n11 ), .A2(PermutationOutput3[38]), 
        .ZN(\Red_SubCellInst3_LFInst_9_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_9_LFInst_0_U7  ( .A(
        \Red_SubCellInst3_LFInst_9_LFInst_0_n10 ), .B(
        \Red_SubCellInst3_LFInst_9_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst3_LFInst_9_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_9_LFInst_0_U6  ( .A1(
        PermutationOutput3[39]), .A2(\Red_SubCellInst3_LFInst_9_LFInst_0_n11 ), 
        .ZN(\Red_SubCellInst3_LFInst_9_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst3_LFInst_9_LFInst_0_U5  ( .A(PermutationOutput3[37]), 
        .ZN(\Red_SubCellInst3_LFInst_9_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_9_LFInst_0_U4  ( .A1(
        PermutationOutput3[38]), .A2(\Red_SubCellInst3_LFInst_9_LFInst_0_n8 ), 
        .ZN(\Red_SubCellInst3_LFInst_9_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst3_LFInst_9_LFInst_0_U3  ( .A(PermutationOutput3[36]), 
        .ZN(\Red_SubCellInst3_LFInst_9_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_9_LFInst_1_U8  ( .A1(
        \Red_SubCellInst3_LFInst_9_LFInst_1_n15 ), .A2(
        \Red_SubCellInst3_LFInst_9_LFInst_1_n14 ), .ZN(Red_Feedback3[37]) );
  NAND2_X1 \Red_SubCellInst3_LFInst_9_LFInst_1_U7  ( .A1(
        \Red_SubCellInst3_LFInst_9_LFInst_1_n13 ), .A2(PermutationOutput3[37]), 
        .ZN(\Red_SubCellInst3_LFInst_9_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_9_LFInst_1_U6  ( .A1(
        \Red_SubCellInst3_LFInst_9_LFInst_1_n12 ), .A2(PermutationOutput3[36]), 
        .ZN(\Red_SubCellInst3_LFInst_9_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_9_LFInst_1_U5  ( .A1(
        PermutationOutput3[39]), .A2(PermutationOutput3[38]), .ZN(
        \Red_SubCellInst3_LFInst_9_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst3_LFInst_9_LFInst_1_U4  ( .A1(PermutationOutput3[38]), 
        .A2(\Red_SubCellInst3_LFInst_9_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst3_LFInst_9_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_9_LFInst_1_U3  ( .A(PermutationOutput3[36]), .B(PermutationOutput3[39]), .ZN(\Red_SubCellInst3_LFInst_9_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_9_LFInst_2_U10  ( .A1(
        \Red_SubCellInst3_LFInst_9_LFInst_2_n19 ), .A2(
        \Red_SubCellInst3_LFInst_9_LFInst_2_n18 ), .ZN(Red_Feedback3[38]) );
  AND2_X1 \Red_SubCellInst3_LFInst_9_LFInst_2_U9  ( .A1(
        \Red_SubCellInst3_LFInst_9_LFInst_2_n17 ), .A2(PermutationOutput3[36]), 
        .ZN(\Red_SubCellInst3_LFInst_9_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_9_LFInst_2_U8  ( .A1(PermutationOutput3[38]), .A2(PermutationOutput3[37]), .ZN(\Red_SubCellInst3_LFInst_9_LFInst_2_n17 )
         );
  XNOR2_X1 \Red_SubCellInst3_LFInst_9_LFInst_2_U7  ( .A(
        \Red_SubCellInst3_LFInst_9_LFInst_2_n16 ), .B(
        \Red_SubCellInst3_LFInst_9_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst3_LFInst_9_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_9_LFInst_2_U6  ( .A1(PermutationOutput3[39]), .A2(\Red_SubCellInst3_LFInst_9_LFInst_2_n14 ), .ZN(
        \Red_SubCellInst3_LFInst_9_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst3_LFInst_9_LFInst_2_U5  ( .A(PermutationOutput3[37]), 
        .ZN(\Red_SubCellInst3_LFInst_9_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_9_LFInst_2_U4  ( .A1(
        PermutationOutput3[38]), .A2(\Red_SubCellInst3_LFInst_9_LFInst_2_n13 ), 
        .ZN(\Red_SubCellInst3_LFInst_9_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst3_LFInst_9_LFInst_2_U3  ( .A(PermutationOutput3[36]), 
        .ZN(\Red_SubCellInst3_LFInst_9_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_9_LFInst_3_U6  ( .A(PermutationOutput3[37]), .B(\Red_SubCellInst3_LFInst_9_LFInst_3_n8 ), .ZN(Red_Feedback3[39]) );
  NOR2_X1 \Red_SubCellInst3_LFInst_9_LFInst_3_U5  ( .A1(
        \Red_SubCellInst3_LFInst_9_LFInst_3_n7 ), .A2(
        \Red_SubCellInst3_LFInst_9_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst3_LFInst_9_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_9_LFInst_3_U4  ( .A1(PermutationOutput3[38]), .A2(PermutationOutput3[39]), .ZN(\Red_SubCellInst3_LFInst_9_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst3_LFInst_9_LFInst_3_U3  ( .A1(PermutationOutput3[39]), .A2(PermutationOutput3[36]), .ZN(\Red_SubCellInst3_LFInst_9_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_10_LFInst_0_U10  ( .A1(
        \Red_SubCellInst3_LFInst_10_LFInst_0_n14 ), .A2(
        \Red_SubCellInst3_LFInst_10_LFInst_0_n13 ), .ZN(Red_Feedback3[40]) );
  NAND2_X1 \Red_SubCellInst3_LFInst_10_LFInst_0_U9  ( .A1(
        PermutationOutput3[40]), .A2(\Red_SubCellInst3_LFInst_10_LFInst_0_n12 ), .ZN(\Red_SubCellInst3_LFInst_10_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_10_LFInst_0_U8  ( .A1(
        \Red_SubCellInst3_LFInst_10_LFInst_0_n11 ), .A2(PermutationOutput3[42]), .ZN(\Red_SubCellInst3_LFInst_10_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_10_LFInst_0_U7  ( .A(
        \Red_SubCellInst3_LFInst_10_LFInst_0_n10 ), .B(
        \Red_SubCellInst3_LFInst_10_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst3_LFInst_10_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_10_LFInst_0_U6  ( .A1(
        PermutationOutput3[43]), .A2(\Red_SubCellInst3_LFInst_10_LFInst_0_n11 ), .ZN(\Red_SubCellInst3_LFInst_10_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst3_LFInst_10_LFInst_0_U5  ( .A(PermutationOutput3[41]), 
        .ZN(\Red_SubCellInst3_LFInst_10_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_10_LFInst_0_U4  ( .A1(
        PermutationOutput3[42]), .A2(\Red_SubCellInst3_LFInst_10_LFInst_0_n8 ), 
        .ZN(\Red_SubCellInst3_LFInst_10_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst3_LFInst_10_LFInst_0_U3  ( .A(PermutationOutput3[40]), 
        .ZN(\Red_SubCellInst3_LFInst_10_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_10_LFInst_1_U8  ( .A1(
        \Red_SubCellInst3_LFInst_10_LFInst_1_n15 ), .A2(
        \Red_SubCellInst3_LFInst_10_LFInst_1_n14 ), .ZN(Red_Feedback3[41]) );
  NAND2_X1 \Red_SubCellInst3_LFInst_10_LFInst_1_U7  ( .A1(
        \Red_SubCellInst3_LFInst_10_LFInst_1_n13 ), .A2(PermutationOutput3[41]), .ZN(\Red_SubCellInst3_LFInst_10_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_10_LFInst_1_U6  ( .A1(
        \Red_SubCellInst3_LFInst_10_LFInst_1_n12 ), .A2(PermutationOutput3[40]), .ZN(\Red_SubCellInst3_LFInst_10_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_10_LFInst_1_U5  ( .A1(
        PermutationOutput3[43]), .A2(PermutationOutput3[42]), .ZN(
        \Red_SubCellInst3_LFInst_10_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst3_LFInst_10_LFInst_1_U4  ( .A1(PermutationOutput3[42]), .A2(\Red_SubCellInst3_LFInst_10_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst3_LFInst_10_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_10_LFInst_1_U3  ( .A(
        PermutationOutput3[40]), .B(PermutationOutput3[43]), .ZN(
        \Red_SubCellInst3_LFInst_10_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_10_LFInst_2_U10  ( .A1(
        \Red_SubCellInst3_LFInst_10_LFInst_2_n19 ), .A2(
        \Red_SubCellInst3_LFInst_10_LFInst_2_n18 ), .ZN(Red_Feedback3[42]) );
  AND2_X1 \Red_SubCellInst3_LFInst_10_LFInst_2_U9  ( .A1(
        \Red_SubCellInst3_LFInst_10_LFInst_2_n17 ), .A2(PermutationOutput3[40]), .ZN(\Red_SubCellInst3_LFInst_10_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_10_LFInst_2_U8  ( .A1(
        PermutationOutput3[42]), .A2(PermutationOutput3[41]), .ZN(
        \Red_SubCellInst3_LFInst_10_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_10_LFInst_2_U7  ( .A(
        \Red_SubCellInst3_LFInst_10_LFInst_2_n16 ), .B(
        \Red_SubCellInst3_LFInst_10_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst3_LFInst_10_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_10_LFInst_2_U6  ( .A1(
        PermutationOutput3[43]), .A2(\Red_SubCellInst3_LFInst_10_LFInst_2_n14 ), .ZN(\Red_SubCellInst3_LFInst_10_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst3_LFInst_10_LFInst_2_U5  ( .A(PermutationOutput3[41]), 
        .ZN(\Red_SubCellInst3_LFInst_10_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_10_LFInst_2_U4  ( .A1(
        PermutationOutput3[42]), .A2(\Red_SubCellInst3_LFInst_10_LFInst_2_n13 ), .ZN(\Red_SubCellInst3_LFInst_10_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst3_LFInst_10_LFInst_2_U3  ( .A(PermutationOutput3[40]), 
        .ZN(\Red_SubCellInst3_LFInst_10_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_10_LFInst_3_U6  ( .A(
        PermutationOutput3[41]), .B(\Red_SubCellInst3_LFInst_10_LFInst_3_n8 ), 
        .ZN(Red_Feedback3[43]) );
  NOR2_X1 \Red_SubCellInst3_LFInst_10_LFInst_3_U5  ( .A1(
        \Red_SubCellInst3_LFInst_10_LFInst_3_n7 ), .A2(
        \Red_SubCellInst3_LFInst_10_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst3_LFInst_10_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_10_LFInst_3_U4  ( .A1(
        PermutationOutput3[42]), .A2(PermutationOutput3[43]), .ZN(
        \Red_SubCellInst3_LFInst_10_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst3_LFInst_10_LFInst_3_U3  ( .A1(
        PermutationOutput3[43]), .A2(PermutationOutput3[40]), .ZN(
        \Red_SubCellInst3_LFInst_10_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_11_LFInst_0_U10  ( .A1(
        \Red_SubCellInst3_LFInst_11_LFInst_0_n14 ), .A2(
        \Red_SubCellInst3_LFInst_11_LFInst_0_n13 ), .ZN(Red_Feedback3[44]) );
  NAND2_X1 \Red_SubCellInst3_LFInst_11_LFInst_0_U9  ( .A1(
        PermutationOutput3[44]), .A2(\Red_SubCellInst3_LFInst_11_LFInst_0_n12 ), .ZN(\Red_SubCellInst3_LFInst_11_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_11_LFInst_0_U8  ( .A1(
        \Red_SubCellInst3_LFInst_11_LFInst_0_n11 ), .A2(PermutationOutput3[46]), .ZN(\Red_SubCellInst3_LFInst_11_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_11_LFInst_0_U7  ( .A(
        \Red_SubCellInst3_LFInst_11_LFInst_0_n10 ), .B(
        \Red_SubCellInst3_LFInst_11_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst3_LFInst_11_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_11_LFInst_0_U6  ( .A1(
        PermutationOutput3[47]), .A2(\Red_SubCellInst3_LFInst_11_LFInst_0_n11 ), .ZN(\Red_SubCellInst3_LFInst_11_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst3_LFInst_11_LFInst_0_U5  ( .A(PermutationOutput3[45]), 
        .ZN(\Red_SubCellInst3_LFInst_11_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_11_LFInst_0_U4  ( .A1(
        PermutationOutput3[46]), .A2(\Red_SubCellInst3_LFInst_11_LFInst_0_n8 ), 
        .ZN(\Red_SubCellInst3_LFInst_11_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst3_LFInst_11_LFInst_0_U3  ( .A(PermutationOutput3[44]), 
        .ZN(\Red_SubCellInst3_LFInst_11_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_11_LFInst_1_U8  ( .A1(
        \Red_SubCellInst3_LFInst_11_LFInst_1_n15 ), .A2(
        \Red_SubCellInst3_LFInst_11_LFInst_1_n14 ), .ZN(Red_Feedback3[45]) );
  NAND2_X1 \Red_SubCellInst3_LFInst_11_LFInst_1_U7  ( .A1(
        \Red_SubCellInst3_LFInst_11_LFInst_1_n13 ), .A2(PermutationOutput3[45]), .ZN(\Red_SubCellInst3_LFInst_11_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_11_LFInst_1_U6  ( .A1(
        \Red_SubCellInst3_LFInst_11_LFInst_1_n12 ), .A2(PermutationOutput3[44]), .ZN(\Red_SubCellInst3_LFInst_11_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_11_LFInst_1_U5  ( .A1(
        PermutationOutput3[47]), .A2(PermutationOutput3[46]), .ZN(
        \Red_SubCellInst3_LFInst_11_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst3_LFInst_11_LFInst_1_U4  ( .A1(PermutationOutput3[46]), .A2(\Red_SubCellInst3_LFInst_11_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst3_LFInst_11_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_11_LFInst_1_U3  ( .A(
        PermutationOutput3[44]), .B(PermutationOutput3[47]), .ZN(
        \Red_SubCellInst3_LFInst_11_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_11_LFInst_2_U10  ( .A1(
        \Red_SubCellInst3_LFInst_11_LFInst_2_n19 ), .A2(
        \Red_SubCellInst3_LFInst_11_LFInst_2_n18 ), .ZN(Red_Feedback3[46]) );
  AND2_X1 \Red_SubCellInst3_LFInst_11_LFInst_2_U9  ( .A1(
        \Red_SubCellInst3_LFInst_11_LFInst_2_n17 ), .A2(PermutationOutput3[44]), .ZN(\Red_SubCellInst3_LFInst_11_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_11_LFInst_2_U8  ( .A1(
        PermutationOutput3[46]), .A2(PermutationOutput3[45]), .ZN(
        \Red_SubCellInst3_LFInst_11_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_11_LFInst_2_U7  ( .A(
        \Red_SubCellInst3_LFInst_11_LFInst_2_n16 ), .B(
        \Red_SubCellInst3_LFInst_11_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst3_LFInst_11_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_11_LFInst_2_U6  ( .A1(
        PermutationOutput3[47]), .A2(\Red_SubCellInst3_LFInst_11_LFInst_2_n14 ), .ZN(\Red_SubCellInst3_LFInst_11_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst3_LFInst_11_LFInst_2_U5  ( .A(PermutationOutput3[45]), 
        .ZN(\Red_SubCellInst3_LFInst_11_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_11_LFInst_2_U4  ( .A1(
        PermutationOutput3[46]), .A2(\Red_SubCellInst3_LFInst_11_LFInst_2_n13 ), .ZN(\Red_SubCellInst3_LFInst_11_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst3_LFInst_11_LFInst_2_U3  ( .A(PermutationOutput3[44]), 
        .ZN(\Red_SubCellInst3_LFInst_11_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_11_LFInst_3_U6  ( .A(
        PermutationOutput3[45]), .B(\Red_SubCellInst3_LFInst_11_LFInst_3_n8 ), 
        .ZN(Red_Feedback3[47]) );
  NOR2_X1 \Red_SubCellInst3_LFInst_11_LFInst_3_U5  ( .A1(
        \Red_SubCellInst3_LFInst_11_LFInst_3_n7 ), .A2(
        \Red_SubCellInst3_LFInst_11_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst3_LFInst_11_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_11_LFInst_3_U4  ( .A1(
        PermutationOutput3[46]), .A2(PermutationOutput3[47]), .ZN(
        \Red_SubCellInst3_LFInst_11_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst3_LFInst_11_LFInst_3_U3  ( .A1(
        PermutationOutput3[47]), .A2(PermutationOutput3[44]), .ZN(
        \Red_SubCellInst3_LFInst_11_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_12_LFInst_0_U10  ( .A1(
        \Red_SubCellInst3_LFInst_12_LFInst_0_n14 ), .A2(
        \Red_SubCellInst3_LFInst_12_LFInst_0_n13 ), .ZN(Red_Feedback3[48]) );
  NAND2_X1 \Red_SubCellInst3_LFInst_12_LFInst_0_U9  ( .A1(
        PermutationOutput3[48]), .A2(\Red_SubCellInst3_LFInst_12_LFInst_0_n12 ), .ZN(\Red_SubCellInst3_LFInst_12_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_12_LFInst_0_U8  ( .A1(
        \Red_SubCellInst3_LFInst_12_LFInst_0_n11 ), .A2(PermutationOutput3[50]), .ZN(\Red_SubCellInst3_LFInst_12_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_12_LFInst_0_U7  ( .A(
        \Red_SubCellInst3_LFInst_12_LFInst_0_n10 ), .B(
        \Red_SubCellInst3_LFInst_12_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst3_LFInst_12_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_12_LFInst_0_U6  ( .A1(
        PermutationOutput3[51]), .A2(\Red_SubCellInst3_LFInst_12_LFInst_0_n11 ), .ZN(\Red_SubCellInst3_LFInst_12_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst3_LFInst_12_LFInst_0_U5  ( .A(PermutationOutput3[49]), 
        .ZN(\Red_SubCellInst3_LFInst_12_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_12_LFInst_0_U4  ( .A1(
        PermutationOutput3[50]), .A2(\Red_SubCellInst3_LFInst_12_LFInst_0_n8 ), 
        .ZN(\Red_SubCellInst3_LFInst_12_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst3_LFInst_12_LFInst_0_U3  ( .A(PermutationOutput3[48]), 
        .ZN(\Red_SubCellInst3_LFInst_12_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_12_LFInst_1_U8  ( .A1(
        \Red_SubCellInst3_LFInst_12_LFInst_1_n15 ), .A2(
        \Red_SubCellInst3_LFInst_12_LFInst_1_n14 ), .ZN(Red_Feedback3[49]) );
  NAND2_X1 \Red_SubCellInst3_LFInst_12_LFInst_1_U7  ( .A1(
        \Red_SubCellInst3_LFInst_12_LFInst_1_n13 ), .A2(PermutationOutput3[49]), .ZN(\Red_SubCellInst3_LFInst_12_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_12_LFInst_1_U6  ( .A1(
        \Red_SubCellInst3_LFInst_12_LFInst_1_n12 ), .A2(PermutationOutput3[48]), .ZN(\Red_SubCellInst3_LFInst_12_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_12_LFInst_1_U5  ( .A1(
        PermutationOutput3[51]), .A2(PermutationOutput3[50]), .ZN(
        \Red_SubCellInst3_LFInst_12_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst3_LFInst_12_LFInst_1_U4  ( .A1(PermutationOutput3[50]), .A2(\Red_SubCellInst3_LFInst_12_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst3_LFInst_12_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_12_LFInst_1_U3  ( .A(
        PermutationOutput3[48]), .B(PermutationOutput3[51]), .ZN(
        \Red_SubCellInst3_LFInst_12_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_12_LFInst_2_U10  ( .A1(
        \Red_SubCellInst3_LFInst_12_LFInst_2_n19 ), .A2(
        \Red_SubCellInst3_LFInst_12_LFInst_2_n18 ), .ZN(Red_Feedback3[50]) );
  AND2_X1 \Red_SubCellInst3_LFInst_12_LFInst_2_U9  ( .A1(
        \Red_SubCellInst3_LFInst_12_LFInst_2_n17 ), .A2(PermutationOutput3[48]), .ZN(\Red_SubCellInst3_LFInst_12_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_12_LFInst_2_U8  ( .A1(
        PermutationOutput3[50]), .A2(PermutationOutput3[49]), .ZN(
        \Red_SubCellInst3_LFInst_12_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_12_LFInst_2_U7  ( .A(
        \Red_SubCellInst3_LFInst_12_LFInst_2_n16 ), .B(
        \Red_SubCellInst3_LFInst_12_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst3_LFInst_12_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_12_LFInst_2_U6  ( .A1(
        PermutationOutput3[51]), .A2(\Red_SubCellInst3_LFInst_12_LFInst_2_n14 ), .ZN(\Red_SubCellInst3_LFInst_12_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst3_LFInst_12_LFInst_2_U5  ( .A(PermutationOutput3[49]), 
        .ZN(\Red_SubCellInst3_LFInst_12_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_12_LFInst_2_U4  ( .A1(
        PermutationOutput3[50]), .A2(\Red_SubCellInst3_LFInst_12_LFInst_2_n13 ), .ZN(\Red_SubCellInst3_LFInst_12_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst3_LFInst_12_LFInst_2_U3  ( .A(PermutationOutput3[48]), 
        .ZN(\Red_SubCellInst3_LFInst_12_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_12_LFInst_3_U6  ( .A(
        PermutationOutput3[49]), .B(\Red_SubCellInst3_LFInst_12_LFInst_3_n8 ), 
        .ZN(Red_Feedback3[51]) );
  NOR2_X1 \Red_SubCellInst3_LFInst_12_LFInst_3_U5  ( .A1(
        \Red_SubCellInst3_LFInst_12_LFInst_3_n7 ), .A2(
        \Red_SubCellInst3_LFInst_12_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst3_LFInst_12_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_12_LFInst_3_U4  ( .A1(
        PermutationOutput3[50]), .A2(PermutationOutput3[51]), .ZN(
        \Red_SubCellInst3_LFInst_12_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst3_LFInst_12_LFInst_3_U3  ( .A1(
        PermutationOutput3[51]), .A2(PermutationOutput3[48]), .ZN(
        \Red_SubCellInst3_LFInst_12_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_13_LFInst_0_U10  ( .A1(
        \Red_SubCellInst3_LFInst_13_LFInst_0_n14 ), .A2(
        \Red_SubCellInst3_LFInst_13_LFInst_0_n13 ), .ZN(Red_Feedback3[52]) );
  NAND2_X1 \Red_SubCellInst3_LFInst_13_LFInst_0_U9  ( .A1(
        PermutationOutput3[52]), .A2(\Red_SubCellInst3_LFInst_13_LFInst_0_n12 ), .ZN(\Red_SubCellInst3_LFInst_13_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_13_LFInst_0_U8  ( .A1(
        \Red_SubCellInst3_LFInst_13_LFInst_0_n11 ), .A2(PermutationOutput3[54]), .ZN(\Red_SubCellInst3_LFInst_13_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_13_LFInst_0_U7  ( .A(
        \Red_SubCellInst3_LFInst_13_LFInst_0_n10 ), .B(
        \Red_SubCellInst3_LFInst_13_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst3_LFInst_13_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_13_LFInst_0_U6  ( .A1(
        PermutationOutput3[55]), .A2(\Red_SubCellInst3_LFInst_13_LFInst_0_n11 ), .ZN(\Red_SubCellInst3_LFInst_13_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst3_LFInst_13_LFInst_0_U5  ( .A(PermutationOutput3[53]), 
        .ZN(\Red_SubCellInst3_LFInst_13_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_13_LFInst_0_U4  ( .A1(
        PermutationOutput3[54]), .A2(\Red_SubCellInst3_LFInst_13_LFInst_0_n8 ), 
        .ZN(\Red_SubCellInst3_LFInst_13_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst3_LFInst_13_LFInst_0_U3  ( .A(PermutationOutput3[52]), 
        .ZN(\Red_SubCellInst3_LFInst_13_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_13_LFInst_1_U8  ( .A1(
        \Red_SubCellInst3_LFInst_13_LFInst_1_n15 ), .A2(
        \Red_SubCellInst3_LFInst_13_LFInst_1_n14 ), .ZN(Red_Feedback3[53]) );
  NAND2_X1 \Red_SubCellInst3_LFInst_13_LFInst_1_U7  ( .A1(
        \Red_SubCellInst3_LFInst_13_LFInst_1_n13 ), .A2(PermutationOutput3[53]), .ZN(\Red_SubCellInst3_LFInst_13_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_13_LFInst_1_U6  ( .A1(
        \Red_SubCellInst3_LFInst_13_LFInst_1_n12 ), .A2(PermutationOutput3[52]), .ZN(\Red_SubCellInst3_LFInst_13_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_13_LFInst_1_U5  ( .A1(
        PermutationOutput3[55]), .A2(PermutationOutput3[54]), .ZN(
        \Red_SubCellInst3_LFInst_13_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst3_LFInst_13_LFInst_1_U4  ( .A1(PermutationOutput3[54]), .A2(\Red_SubCellInst3_LFInst_13_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst3_LFInst_13_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_13_LFInst_1_U3  ( .A(
        PermutationOutput3[52]), .B(PermutationOutput3[55]), .ZN(
        \Red_SubCellInst3_LFInst_13_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_13_LFInst_2_U10  ( .A1(
        \Red_SubCellInst3_LFInst_13_LFInst_2_n19 ), .A2(
        \Red_SubCellInst3_LFInst_13_LFInst_2_n18 ), .ZN(Red_Feedback3[54]) );
  AND2_X1 \Red_SubCellInst3_LFInst_13_LFInst_2_U9  ( .A1(
        \Red_SubCellInst3_LFInst_13_LFInst_2_n17 ), .A2(PermutationOutput3[52]), .ZN(\Red_SubCellInst3_LFInst_13_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_13_LFInst_2_U8  ( .A1(
        PermutationOutput3[54]), .A2(PermutationOutput3[53]), .ZN(
        \Red_SubCellInst3_LFInst_13_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_13_LFInst_2_U7  ( .A(
        \Red_SubCellInst3_LFInst_13_LFInst_2_n16 ), .B(
        \Red_SubCellInst3_LFInst_13_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst3_LFInst_13_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_13_LFInst_2_U6  ( .A1(
        PermutationOutput3[55]), .A2(\Red_SubCellInst3_LFInst_13_LFInst_2_n14 ), .ZN(\Red_SubCellInst3_LFInst_13_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst3_LFInst_13_LFInst_2_U5  ( .A(PermutationOutput3[53]), 
        .ZN(\Red_SubCellInst3_LFInst_13_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_13_LFInst_2_U4  ( .A1(
        PermutationOutput3[54]), .A2(\Red_SubCellInst3_LFInst_13_LFInst_2_n13 ), .ZN(\Red_SubCellInst3_LFInst_13_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst3_LFInst_13_LFInst_2_U3  ( .A(PermutationOutput3[52]), 
        .ZN(\Red_SubCellInst3_LFInst_13_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_13_LFInst_3_U6  ( .A(
        PermutationOutput3[53]), .B(\Red_SubCellInst3_LFInst_13_LFInst_3_n8 ), 
        .ZN(Red_Feedback3[55]) );
  NOR2_X1 \Red_SubCellInst3_LFInst_13_LFInst_3_U5  ( .A1(
        \Red_SubCellInst3_LFInst_13_LFInst_3_n7 ), .A2(
        \Red_SubCellInst3_LFInst_13_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst3_LFInst_13_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_13_LFInst_3_U4  ( .A1(
        PermutationOutput3[54]), .A2(PermutationOutput3[55]), .ZN(
        \Red_SubCellInst3_LFInst_13_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst3_LFInst_13_LFInst_3_U3  ( .A1(
        PermutationOutput3[55]), .A2(PermutationOutput3[52]), .ZN(
        \Red_SubCellInst3_LFInst_13_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_14_LFInst_0_U10  ( .A1(
        \Red_SubCellInst3_LFInst_14_LFInst_0_n14 ), .A2(
        \Red_SubCellInst3_LFInst_14_LFInst_0_n13 ), .ZN(Red_Feedback3[56]) );
  NAND2_X1 \Red_SubCellInst3_LFInst_14_LFInst_0_U9  ( .A1(
        PermutationOutput3[56]), .A2(\Red_SubCellInst3_LFInst_14_LFInst_0_n12 ), .ZN(\Red_SubCellInst3_LFInst_14_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_14_LFInst_0_U8  ( .A1(
        \Red_SubCellInst3_LFInst_14_LFInst_0_n11 ), .A2(PermutationOutput3[58]), .ZN(\Red_SubCellInst3_LFInst_14_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_14_LFInst_0_U7  ( .A(
        \Red_SubCellInst3_LFInst_14_LFInst_0_n10 ), .B(
        \Red_SubCellInst3_LFInst_14_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst3_LFInst_14_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_14_LFInst_0_U6  ( .A1(
        PermutationOutput3[59]), .A2(\Red_SubCellInst3_LFInst_14_LFInst_0_n11 ), .ZN(\Red_SubCellInst3_LFInst_14_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst3_LFInst_14_LFInst_0_U5  ( .A(PermutationOutput3[57]), 
        .ZN(\Red_SubCellInst3_LFInst_14_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_14_LFInst_0_U4  ( .A1(
        PermutationOutput3[58]), .A2(\Red_SubCellInst3_LFInst_14_LFInst_0_n8 ), 
        .ZN(\Red_SubCellInst3_LFInst_14_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst3_LFInst_14_LFInst_0_U3  ( .A(PermutationOutput3[56]), 
        .ZN(\Red_SubCellInst3_LFInst_14_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_14_LFInst_1_U8  ( .A1(
        \Red_SubCellInst3_LFInst_14_LFInst_1_n15 ), .A2(
        \Red_SubCellInst3_LFInst_14_LFInst_1_n14 ), .ZN(Red_Feedback3[57]) );
  NAND2_X1 \Red_SubCellInst3_LFInst_14_LFInst_1_U7  ( .A1(
        \Red_SubCellInst3_LFInst_14_LFInst_1_n13 ), .A2(PermutationOutput3[57]), .ZN(\Red_SubCellInst3_LFInst_14_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_14_LFInst_1_U6  ( .A1(
        \Red_SubCellInst3_LFInst_14_LFInst_1_n12 ), .A2(PermutationOutput3[56]), .ZN(\Red_SubCellInst3_LFInst_14_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_14_LFInst_1_U5  ( .A1(
        PermutationOutput3[59]), .A2(PermutationOutput3[58]), .ZN(
        \Red_SubCellInst3_LFInst_14_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst3_LFInst_14_LFInst_1_U4  ( .A1(PermutationOutput3[58]), .A2(\Red_SubCellInst3_LFInst_14_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst3_LFInst_14_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_14_LFInst_1_U3  ( .A(
        PermutationOutput3[56]), .B(PermutationOutput3[59]), .ZN(
        \Red_SubCellInst3_LFInst_14_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_14_LFInst_2_U10  ( .A1(
        \Red_SubCellInst3_LFInst_14_LFInst_2_n19 ), .A2(
        \Red_SubCellInst3_LFInst_14_LFInst_2_n18 ), .ZN(Red_Feedback3[58]) );
  AND2_X1 \Red_SubCellInst3_LFInst_14_LFInst_2_U9  ( .A1(
        \Red_SubCellInst3_LFInst_14_LFInst_2_n17 ), .A2(PermutationOutput3[56]), .ZN(\Red_SubCellInst3_LFInst_14_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_14_LFInst_2_U8  ( .A1(
        PermutationOutput3[58]), .A2(PermutationOutput3[57]), .ZN(
        \Red_SubCellInst3_LFInst_14_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_14_LFInst_2_U7  ( .A(
        \Red_SubCellInst3_LFInst_14_LFInst_2_n16 ), .B(
        \Red_SubCellInst3_LFInst_14_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst3_LFInst_14_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_14_LFInst_2_U6  ( .A1(
        PermutationOutput3[59]), .A2(\Red_SubCellInst3_LFInst_14_LFInst_2_n14 ), .ZN(\Red_SubCellInst3_LFInst_14_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst3_LFInst_14_LFInst_2_U5  ( .A(PermutationOutput3[57]), 
        .ZN(\Red_SubCellInst3_LFInst_14_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_14_LFInst_2_U4  ( .A1(
        PermutationOutput3[58]), .A2(\Red_SubCellInst3_LFInst_14_LFInst_2_n13 ), .ZN(\Red_SubCellInst3_LFInst_14_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst3_LFInst_14_LFInst_2_U3  ( .A(PermutationOutput3[56]), 
        .ZN(\Red_SubCellInst3_LFInst_14_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_14_LFInst_3_U6  ( .A(
        PermutationOutput3[57]), .B(\Red_SubCellInst3_LFInst_14_LFInst_3_n8 ), 
        .ZN(Red_Feedback3[59]) );
  NOR2_X1 \Red_SubCellInst3_LFInst_14_LFInst_3_U5  ( .A1(
        \Red_SubCellInst3_LFInst_14_LFInst_3_n7 ), .A2(
        \Red_SubCellInst3_LFInst_14_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst3_LFInst_14_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_14_LFInst_3_U4  ( .A1(
        PermutationOutput3[58]), .A2(PermutationOutput3[59]), .ZN(
        \Red_SubCellInst3_LFInst_14_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst3_LFInst_14_LFInst_3_U3  ( .A1(
        PermutationOutput3[59]), .A2(PermutationOutput3[56]), .ZN(
        \Red_SubCellInst3_LFInst_14_LFInst_3_n7 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_15_LFInst_0_U10  ( .A1(
        \Red_SubCellInst3_LFInst_15_LFInst_0_n14 ), .A2(
        \Red_SubCellInst3_LFInst_15_LFInst_0_n13 ), .ZN(Red_Feedback3[60]) );
  NAND2_X1 \Red_SubCellInst3_LFInst_15_LFInst_0_U9  ( .A1(
        PermutationOutput3[60]), .A2(\Red_SubCellInst3_LFInst_15_LFInst_0_n12 ), .ZN(\Red_SubCellInst3_LFInst_15_LFInst_0_n13 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_15_LFInst_0_U8  ( .A1(
        \Red_SubCellInst3_LFInst_15_LFInst_0_n11 ), .A2(PermutationOutput3[62]), .ZN(\Red_SubCellInst3_LFInst_15_LFInst_0_n12 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_15_LFInst_0_U7  ( .A(
        \Red_SubCellInst3_LFInst_15_LFInst_0_n10 ), .B(
        \Red_SubCellInst3_LFInst_15_LFInst_0_n9 ), .ZN(
        \Red_SubCellInst3_LFInst_15_LFInst_0_n14 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_15_LFInst_0_U6  ( .A1(
        PermutationOutput3[63]), .A2(\Red_SubCellInst3_LFInst_15_LFInst_0_n11 ), .ZN(\Red_SubCellInst3_LFInst_15_LFInst_0_n9 ) );
  INV_X1 \Red_SubCellInst3_LFInst_15_LFInst_0_U5  ( .A(PermutationOutput3[61]), 
        .ZN(\Red_SubCellInst3_LFInst_15_LFInst_0_n11 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_15_LFInst_0_U4  ( .A1(
        PermutationOutput3[62]), .A2(\Red_SubCellInst3_LFInst_15_LFInst_0_n8 ), 
        .ZN(\Red_SubCellInst3_LFInst_15_LFInst_0_n10 ) );
  INV_X1 \Red_SubCellInst3_LFInst_15_LFInst_0_U3  ( .A(PermutationOutput3[60]), 
        .ZN(\Red_SubCellInst3_LFInst_15_LFInst_0_n8 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_15_LFInst_1_U8  ( .A1(
        \Red_SubCellInst3_LFInst_15_LFInst_1_n15 ), .A2(
        \Red_SubCellInst3_LFInst_15_LFInst_1_n14 ), .ZN(Red_Feedback3[61]) );
  NAND2_X1 \Red_SubCellInst3_LFInst_15_LFInst_1_U7  ( .A1(
        \Red_SubCellInst3_LFInst_15_LFInst_1_n13 ), .A2(PermutationOutput3[61]), .ZN(\Red_SubCellInst3_LFInst_15_LFInst_1_n14 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_15_LFInst_1_U6  ( .A1(
        \Red_SubCellInst3_LFInst_15_LFInst_1_n12 ), .A2(PermutationOutput3[60]), .ZN(\Red_SubCellInst3_LFInst_15_LFInst_1_n13 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_15_LFInst_1_U5  ( .A1(
        PermutationOutput3[63]), .A2(PermutationOutput3[62]), .ZN(
        \Red_SubCellInst3_LFInst_15_LFInst_1_n12 ) );
  OR2_X1 \Red_SubCellInst3_LFInst_15_LFInst_1_U4  ( .A1(PermutationOutput3[62]), .A2(\Red_SubCellInst3_LFInst_15_LFInst_1_n11 ), .ZN(
        \Red_SubCellInst3_LFInst_15_LFInst_1_n15 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_15_LFInst_1_U3  ( .A(
        PermutationOutput3[60]), .B(PermutationOutput3[63]), .ZN(
        \Red_SubCellInst3_LFInst_15_LFInst_1_n11 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_15_LFInst_2_U10  ( .A1(
        \Red_SubCellInst3_LFInst_15_LFInst_2_n19 ), .A2(
        \Red_SubCellInst3_LFInst_15_LFInst_2_n18 ), .ZN(Red_Feedback3[62]) );
  AND2_X1 \Red_SubCellInst3_LFInst_15_LFInst_2_U9  ( .A1(
        \Red_SubCellInst3_LFInst_15_LFInst_2_n17 ), .A2(PermutationOutput3[60]), .ZN(\Red_SubCellInst3_LFInst_15_LFInst_2_n18 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_15_LFInst_2_U8  ( .A1(
        PermutationOutput3[62]), .A2(PermutationOutput3[61]), .ZN(
        \Red_SubCellInst3_LFInst_15_LFInst_2_n17 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_15_LFInst_2_U7  ( .A(
        \Red_SubCellInst3_LFInst_15_LFInst_2_n16 ), .B(
        \Red_SubCellInst3_LFInst_15_LFInst_2_n15 ), .ZN(
        \Red_SubCellInst3_LFInst_15_LFInst_2_n19 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_15_LFInst_2_U6  ( .A1(
        PermutationOutput3[63]), .A2(\Red_SubCellInst3_LFInst_15_LFInst_2_n14 ), .ZN(\Red_SubCellInst3_LFInst_15_LFInst_2_n15 ) );
  INV_X1 \Red_SubCellInst3_LFInst_15_LFInst_2_U5  ( .A(PermutationOutput3[61]), 
        .ZN(\Red_SubCellInst3_LFInst_15_LFInst_2_n14 ) );
  NAND2_X1 \Red_SubCellInst3_LFInst_15_LFInst_2_U4  ( .A1(
        PermutationOutput3[62]), .A2(\Red_SubCellInst3_LFInst_15_LFInst_2_n13 ), .ZN(\Red_SubCellInst3_LFInst_15_LFInst_2_n16 ) );
  INV_X1 \Red_SubCellInst3_LFInst_15_LFInst_2_U3  ( .A(PermutationOutput3[60]), 
        .ZN(\Red_SubCellInst3_LFInst_15_LFInst_2_n13 ) );
  XNOR2_X1 \Red_SubCellInst3_LFInst_15_LFInst_3_U6  ( .A(
        PermutationOutput3[61]), .B(\Red_SubCellInst3_LFInst_15_LFInst_3_n8 ), 
        .ZN(Red_Feedback3[63]) );
  NOR2_X1 \Red_SubCellInst3_LFInst_15_LFInst_3_U5  ( .A1(
        \Red_SubCellInst3_LFInst_15_LFInst_3_n7 ), .A2(
        \Red_SubCellInst3_LFInst_15_LFInst_3_n6 ), .ZN(
        \Red_SubCellInst3_LFInst_15_LFInst_3_n8 ) );
  NOR2_X1 \Red_SubCellInst3_LFInst_15_LFInst_3_U4  ( .A1(
        PermutationOutput3[62]), .A2(PermutationOutput3[63]), .ZN(
        \Red_SubCellInst3_LFInst_15_LFInst_3_n6 ) );
  AND2_X1 \Red_SubCellInst3_LFInst_15_LFInst_3_U3  ( .A1(
        PermutationOutput3[63]), .A2(PermutationOutput3[60]), .ZN(
        \Red_SubCellInst3_LFInst_15_LFInst_3_n7 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_0_LFInst_0_U4  ( .A(
        \Red_K0Inst_LFInst_0_LFInst_0_n2 ), .B(Key[130]), .ZN(Red_K0[0]) );
  XNOR2_X1 \Red_K0Inst_LFInst_0_LFInst_0_U3  ( .A(Key[131]), .B(Key[129]), 
        .ZN(\Red_K0Inst_LFInst_0_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_0_LFInst_1_U4  ( .A(
        \Red_K0Inst_LFInst_0_LFInst_1_n2 ), .B(Key[130]), .ZN(Red_K0[1]) );
  XNOR2_X1 \Red_K0Inst_LFInst_0_LFInst_1_U3  ( .A(Key[131]), .B(Key[128]), 
        .ZN(\Red_K0Inst_LFInst_0_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_0_LFInst_2_U4  ( .A(
        \Red_K0Inst_LFInst_0_LFInst_2_n2 ), .B(Key[129]), .ZN(Red_K0[2]) );
  XNOR2_X1 \Red_K0Inst_LFInst_0_LFInst_2_U3  ( .A(Key[131]), .B(Key[128]), 
        .ZN(\Red_K0Inst_LFInst_0_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_0_LFInst_3_U4  ( .A(
        \Red_K0Inst_LFInst_0_LFInst_3_n2 ), .B(Key[129]), .ZN(Red_K0[3]) );
  XNOR2_X1 \Red_K0Inst_LFInst_0_LFInst_3_U3  ( .A(Key[130]), .B(Key[128]), 
        .ZN(\Red_K0Inst_LFInst_0_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_1_LFInst_0_U4  ( .A(
        \Red_K0Inst_LFInst_1_LFInst_0_n2 ), .B(Key[134]), .ZN(Red_K0[4]) );
  XNOR2_X1 \Red_K0Inst_LFInst_1_LFInst_0_U3  ( .A(Key[135]), .B(Key[133]), 
        .ZN(\Red_K0Inst_LFInst_1_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_1_LFInst_1_U4  ( .A(
        \Red_K0Inst_LFInst_1_LFInst_1_n2 ), .B(Key[134]), .ZN(Red_K0[5]) );
  XNOR2_X1 \Red_K0Inst_LFInst_1_LFInst_1_U3  ( .A(Key[135]), .B(Key[132]), 
        .ZN(\Red_K0Inst_LFInst_1_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_1_LFInst_2_U4  ( .A(
        \Red_K0Inst_LFInst_1_LFInst_2_n2 ), .B(Key[133]), .ZN(Red_K0[6]) );
  XNOR2_X1 \Red_K0Inst_LFInst_1_LFInst_2_U3  ( .A(Key[135]), .B(Key[132]), 
        .ZN(\Red_K0Inst_LFInst_1_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_1_LFInst_3_U4  ( .A(
        \Red_K0Inst_LFInst_1_LFInst_3_n2 ), .B(Key[133]), .ZN(Red_K0[7]) );
  XNOR2_X1 \Red_K0Inst_LFInst_1_LFInst_3_U3  ( .A(Key[134]), .B(Key[132]), 
        .ZN(\Red_K0Inst_LFInst_1_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_2_LFInst_0_U4  ( .A(
        \Red_K0Inst_LFInst_2_LFInst_0_n2 ), .B(Key[138]), .ZN(Red_K0[8]) );
  XNOR2_X1 \Red_K0Inst_LFInst_2_LFInst_0_U3  ( .A(Key[139]), .B(Key[137]), 
        .ZN(\Red_K0Inst_LFInst_2_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_2_LFInst_1_U4  ( .A(
        \Red_K0Inst_LFInst_2_LFInst_1_n2 ), .B(Key[138]), .ZN(Red_K0[9]) );
  XNOR2_X1 \Red_K0Inst_LFInst_2_LFInst_1_U3  ( .A(Key[139]), .B(Key[136]), 
        .ZN(\Red_K0Inst_LFInst_2_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_2_LFInst_2_U4  ( .A(
        \Red_K0Inst_LFInst_2_LFInst_2_n2 ), .B(Key[137]), .ZN(Red_K0[10]) );
  XNOR2_X1 \Red_K0Inst_LFInst_2_LFInst_2_U3  ( .A(Key[139]), .B(Key[136]), 
        .ZN(\Red_K0Inst_LFInst_2_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_2_LFInst_3_U4  ( .A(
        \Red_K0Inst_LFInst_2_LFInst_3_n2 ), .B(Key[137]), .ZN(Red_K0[11]) );
  XNOR2_X1 \Red_K0Inst_LFInst_2_LFInst_3_U3  ( .A(Key[138]), .B(Key[136]), 
        .ZN(\Red_K0Inst_LFInst_2_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_3_LFInst_0_U4  ( .A(
        \Red_K0Inst_LFInst_3_LFInst_0_n2 ), .B(Key[142]), .ZN(Red_K0[12]) );
  XNOR2_X1 \Red_K0Inst_LFInst_3_LFInst_0_U3  ( .A(Key[143]), .B(Key[141]), 
        .ZN(\Red_K0Inst_LFInst_3_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_3_LFInst_1_U4  ( .A(
        \Red_K0Inst_LFInst_3_LFInst_1_n2 ), .B(Key[142]), .ZN(Red_K0[13]) );
  XNOR2_X1 \Red_K0Inst_LFInst_3_LFInst_1_U3  ( .A(Key[143]), .B(Key[140]), 
        .ZN(\Red_K0Inst_LFInst_3_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_3_LFInst_2_U4  ( .A(
        \Red_K0Inst_LFInst_3_LFInst_2_n2 ), .B(Key[141]), .ZN(Red_K0[14]) );
  XNOR2_X1 \Red_K0Inst_LFInst_3_LFInst_2_U3  ( .A(Key[143]), .B(Key[140]), 
        .ZN(\Red_K0Inst_LFInst_3_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_3_LFInst_3_U4  ( .A(
        \Red_K0Inst_LFInst_3_LFInst_3_n2 ), .B(Key[141]), .ZN(Red_K0[15]) );
  XNOR2_X1 \Red_K0Inst_LFInst_3_LFInst_3_U3  ( .A(Key[142]), .B(Key[140]), 
        .ZN(\Red_K0Inst_LFInst_3_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_4_LFInst_0_U4  ( .A(
        \Red_K0Inst_LFInst_4_LFInst_0_n2 ), .B(Key[146]), .ZN(Red_K0[16]) );
  XNOR2_X1 \Red_K0Inst_LFInst_4_LFInst_0_U3  ( .A(Key[147]), .B(Key[145]), 
        .ZN(\Red_K0Inst_LFInst_4_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_4_LFInst_1_U4  ( .A(
        \Red_K0Inst_LFInst_4_LFInst_1_n2 ), .B(Key[146]), .ZN(Red_K0[17]) );
  XNOR2_X1 \Red_K0Inst_LFInst_4_LFInst_1_U3  ( .A(Key[147]), .B(Key[144]), 
        .ZN(\Red_K0Inst_LFInst_4_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_4_LFInst_2_U4  ( .A(
        \Red_K0Inst_LFInst_4_LFInst_2_n2 ), .B(Key[145]), .ZN(Red_K0[18]) );
  XNOR2_X1 \Red_K0Inst_LFInst_4_LFInst_2_U3  ( .A(Key[147]), .B(Key[144]), 
        .ZN(\Red_K0Inst_LFInst_4_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_4_LFInst_3_U4  ( .A(
        \Red_K0Inst_LFInst_4_LFInst_3_n2 ), .B(Key[145]), .ZN(Red_K0[19]) );
  XNOR2_X1 \Red_K0Inst_LFInst_4_LFInst_3_U3  ( .A(Key[146]), .B(Key[144]), 
        .ZN(\Red_K0Inst_LFInst_4_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_5_LFInst_0_U4  ( .A(
        \Red_K0Inst_LFInst_5_LFInst_0_n2 ), .B(Key[150]), .ZN(Red_K0[20]) );
  XNOR2_X1 \Red_K0Inst_LFInst_5_LFInst_0_U3  ( .A(Key[151]), .B(Key[149]), 
        .ZN(\Red_K0Inst_LFInst_5_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_5_LFInst_1_U4  ( .A(
        \Red_K0Inst_LFInst_5_LFInst_1_n2 ), .B(Key[150]), .ZN(Red_K0[21]) );
  XNOR2_X1 \Red_K0Inst_LFInst_5_LFInst_1_U3  ( .A(Key[151]), .B(Key[148]), 
        .ZN(\Red_K0Inst_LFInst_5_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_5_LFInst_2_U4  ( .A(
        \Red_K0Inst_LFInst_5_LFInst_2_n2 ), .B(Key[149]), .ZN(Red_K0[22]) );
  XNOR2_X1 \Red_K0Inst_LFInst_5_LFInst_2_U3  ( .A(Key[151]), .B(Key[148]), 
        .ZN(\Red_K0Inst_LFInst_5_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_5_LFInst_3_U4  ( .A(
        \Red_K0Inst_LFInst_5_LFInst_3_n2 ), .B(Key[149]), .ZN(Red_K0[23]) );
  XNOR2_X1 \Red_K0Inst_LFInst_5_LFInst_3_U3  ( .A(Key[150]), .B(Key[148]), 
        .ZN(\Red_K0Inst_LFInst_5_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_6_LFInst_0_U4  ( .A(
        \Red_K0Inst_LFInst_6_LFInst_0_n2 ), .B(Key[154]), .ZN(Red_K0[24]) );
  XNOR2_X1 \Red_K0Inst_LFInst_6_LFInst_0_U3  ( .A(Key[155]), .B(Key[153]), 
        .ZN(\Red_K0Inst_LFInst_6_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_6_LFInst_1_U4  ( .A(
        \Red_K0Inst_LFInst_6_LFInst_1_n2 ), .B(Key[154]), .ZN(Red_K0[25]) );
  XNOR2_X1 \Red_K0Inst_LFInst_6_LFInst_1_U3  ( .A(Key[155]), .B(Key[152]), 
        .ZN(\Red_K0Inst_LFInst_6_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_6_LFInst_2_U4  ( .A(
        \Red_K0Inst_LFInst_6_LFInst_2_n2 ), .B(Key[153]), .ZN(Red_K0[26]) );
  XNOR2_X1 \Red_K0Inst_LFInst_6_LFInst_2_U3  ( .A(Key[155]), .B(Key[152]), 
        .ZN(\Red_K0Inst_LFInst_6_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_6_LFInst_3_U4  ( .A(
        \Red_K0Inst_LFInst_6_LFInst_3_n2 ), .B(Key[153]), .ZN(Red_K0[27]) );
  XNOR2_X1 \Red_K0Inst_LFInst_6_LFInst_3_U3  ( .A(Key[154]), .B(Key[152]), 
        .ZN(\Red_K0Inst_LFInst_6_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_7_LFInst_0_U4  ( .A(
        \Red_K0Inst_LFInst_7_LFInst_0_n2 ), .B(Key[158]), .ZN(Red_K0[28]) );
  XNOR2_X1 \Red_K0Inst_LFInst_7_LFInst_0_U3  ( .A(Key[159]), .B(Key[157]), 
        .ZN(\Red_K0Inst_LFInst_7_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_7_LFInst_1_U4  ( .A(
        \Red_K0Inst_LFInst_7_LFInst_1_n2 ), .B(Key[158]), .ZN(Red_K0[29]) );
  XNOR2_X1 \Red_K0Inst_LFInst_7_LFInst_1_U3  ( .A(Key[159]), .B(Key[156]), 
        .ZN(\Red_K0Inst_LFInst_7_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_7_LFInst_2_U4  ( .A(
        \Red_K0Inst_LFInst_7_LFInst_2_n2 ), .B(Key[157]), .ZN(Red_K0[30]) );
  XNOR2_X1 \Red_K0Inst_LFInst_7_LFInst_2_U3  ( .A(Key[159]), .B(Key[156]), 
        .ZN(\Red_K0Inst_LFInst_7_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_7_LFInst_3_U4  ( .A(
        \Red_K0Inst_LFInst_7_LFInst_3_n2 ), .B(Key[157]), .ZN(Red_K0[31]) );
  XNOR2_X1 \Red_K0Inst_LFInst_7_LFInst_3_U3  ( .A(Key[158]), .B(Key[156]), 
        .ZN(\Red_K0Inst_LFInst_7_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_8_LFInst_0_U4  ( .A(
        \Red_K0Inst_LFInst_8_LFInst_0_n2 ), .B(Key[162]), .ZN(Red_K0[32]) );
  XNOR2_X1 \Red_K0Inst_LFInst_8_LFInst_0_U3  ( .A(Key[163]), .B(Key[161]), 
        .ZN(\Red_K0Inst_LFInst_8_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_8_LFInst_1_U4  ( .A(
        \Red_K0Inst_LFInst_8_LFInst_1_n2 ), .B(Key[162]), .ZN(Red_K0[33]) );
  XNOR2_X1 \Red_K0Inst_LFInst_8_LFInst_1_U3  ( .A(Key[163]), .B(Key[160]), 
        .ZN(\Red_K0Inst_LFInst_8_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_8_LFInst_2_U4  ( .A(
        \Red_K0Inst_LFInst_8_LFInst_2_n2 ), .B(Key[161]), .ZN(Red_K0[34]) );
  XNOR2_X1 \Red_K0Inst_LFInst_8_LFInst_2_U3  ( .A(Key[163]), .B(Key[160]), 
        .ZN(\Red_K0Inst_LFInst_8_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_8_LFInst_3_U4  ( .A(
        \Red_K0Inst_LFInst_8_LFInst_3_n2 ), .B(Key[161]), .ZN(Red_K0[35]) );
  XNOR2_X1 \Red_K0Inst_LFInst_8_LFInst_3_U3  ( .A(Key[162]), .B(Key[160]), 
        .ZN(\Red_K0Inst_LFInst_8_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_9_LFInst_0_U4  ( .A(
        \Red_K0Inst_LFInst_9_LFInst_0_n2 ), .B(Key[166]), .ZN(Red_K0[36]) );
  XNOR2_X1 \Red_K0Inst_LFInst_9_LFInst_0_U3  ( .A(Key[167]), .B(Key[165]), 
        .ZN(\Red_K0Inst_LFInst_9_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_9_LFInst_1_U4  ( .A(
        \Red_K0Inst_LFInst_9_LFInst_1_n2 ), .B(Key[166]), .ZN(Red_K0[37]) );
  XNOR2_X1 \Red_K0Inst_LFInst_9_LFInst_1_U3  ( .A(Key[167]), .B(Key[164]), 
        .ZN(\Red_K0Inst_LFInst_9_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_9_LFInst_2_U4  ( .A(
        \Red_K0Inst_LFInst_9_LFInst_2_n2 ), .B(Key[165]), .ZN(Red_K0[38]) );
  XNOR2_X1 \Red_K0Inst_LFInst_9_LFInst_2_U3  ( .A(Key[167]), .B(Key[164]), 
        .ZN(\Red_K0Inst_LFInst_9_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_9_LFInst_3_U4  ( .A(
        \Red_K0Inst_LFInst_9_LFInst_3_n2 ), .B(Key[165]), .ZN(Red_K0[39]) );
  XNOR2_X1 \Red_K0Inst_LFInst_9_LFInst_3_U3  ( .A(Key[166]), .B(Key[164]), 
        .ZN(\Red_K0Inst_LFInst_9_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_10_LFInst_0_U4  ( .A(
        \Red_K0Inst_LFInst_10_LFInst_0_n2 ), .B(Key[170]), .ZN(Red_K0[40]) );
  XNOR2_X1 \Red_K0Inst_LFInst_10_LFInst_0_U3  ( .A(Key[171]), .B(Key[169]), 
        .ZN(\Red_K0Inst_LFInst_10_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_10_LFInst_1_U4  ( .A(
        \Red_K0Inst_LFInst_10_LFInst_1_n2 ), .B(Key[170]), .ZN(Red_K0[41]) );
  XNOR2_X1 \Red_K0Inst_LFInst_10_LFInst_1_U3  ( .A(Key[171]), .B(Key[168]), 
        .ZN(\Red_K0Inst_LFInst_10_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_10_LFInst_2_U4  ( .A(
        \Red_K0Inst_LFInst_10_LFInst_2_n2 ), .B(Key[169]), .ZN(Red_K0[42]) );
  XNOR2_X1 \Red_K0Inst_LFInst_10_LFInst_2_U3  ( .A(Key[171]), .B(Key[168]), 
        .ZN(\Red_K0Inst_LFInst_10_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_10_LFInst_3_U4  ( .A(
        \Red_K0Inst_LFInst_10_LFInst_3_n2 ), .B(Key[169]), .ZN(Red_K0[43]) );
  XNOR2_X1 \Red_K0Inst_LFInst_10_LFInst_3_U3  ( .A(Key[170]), .B(Key[168]), 
        .ZN(\Red_K0Inst_LFInst_10_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_11_LFInst_0_U4  ( .A(
        \Red_K0Inst_LFInst_11_LFInst_0_n2 ), .B(Key[174]), .ZN(Red_K0[44]) );
  XNOR2_X1 \Red_K0Inst_LFInst_11_LFInst_0_U3  ( .A(Key[175]), .B(Key[173]), 
        .ZN(\Red_K0Inst_LFInst_11_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_11_LFInst_1_U4  ( .A(
        \Red_K0Inst_LFInst_11_LFInst_1_n2 ), .B(Key[174]), .ZN(Red_K0[45]) );
  XNOR2_X1 \Red_K0Inst_LFInst_11_LFInst_1_U3  ( .A(Key[175]), .B(Key[172]), 
        .ZN(\Red_K0Inst_LFInst_11_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_11_LFInst_2_U4  ( .A(
        \Red_K0Inst_LFInst_11_LFInst_2_n2 ), .B(Key[173]), .ZN(Red_K0[46]) );
  XNOR2_X1 \Red_K0Inst_LFInst_11_LFInst_2_U3  ( .A(Key[175]), .B(Key[172]), 
        .ZN(\Red_K0Inst_LFInst_11_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_11_LFInst_3_U4  ( .A(
        \Red_K0Inst_LFInst_11_LFInst_3_n2 ), .B(Key[173]), .ZN(Red_K0[47]) );
  XNOR2_X1 \Red_K0Inst_LFInst_11_LFInst_3_U3  ( .A(Key[174]), .B(Key[172]), 
        .ZN(\Red_K0Inst_LFInst_11_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_12_LFInst_0_U4  ( .A(
        \Red_K0Inst_LFInst_12_LFInst_0_n2 ), .B(Key[178]), .ZN(Red_K0[48]) );
  XNOR2_X1 \Red_K0Inst_LFInst_12_LFInst_0_U3  ( .A(Key[179]), .B(Key[177]), 
        .ZN(\Red_K0Inst_LFInst_12_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_12_LFInst_1_U4  ( .A(
        \Red_K0Inst_LFInst_12_LFInst_1_n2 ), .B(Key[178]), .ZN(Red_K0[49]) );
  XNOR2_X1 \Red_K0Inst_LFInst_12_LFInst_1_U3  ( .A(Key[179]), .B(Key[176]), 
        .ZN(\Red_K0Inst_LFInst_12_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_12_LFInst_2_U4  ( .A(
        \Red_K0Inst_LFInst_12_LFInst_2_n2 ), .B(Key[177]), .ZN(Red_K0[50]) );
  XNOR2_X1 \Red_K0Inst_LFInst_12_LFInst_2_U3  ( .A(Key[179]), .B(Key[176]), 
        .ZN(\Red_K0Inst_LFInst_12_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_12_LFInst_3_U4  ( .A(
        \Red_K0Inst_LFInst_12_LFInst_3_n2 ), .B(Key[177]), .ZN(Red_K0[51]) );
  XNOR2_X1 \Red_K0Inst_LFInst_12_LFInst_3_U3  ( .A(Key[178]), .B(Key[176]), 
        .ZN(\Red_K0Inst_LFInst_12_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_13_LFInst_0_U4  ( .A(
        \Red_K0Inst_LFInst_13_LFInst_0_n2 ), .B(Key[182]), .ZN(Red_K0[52]) );
  XNOR2_X1 \Red_K0Inst_LFInst_13_LFInst_0_U3  ( .A(Key[183]), .B(Key[181]), 
        .ZN(\Red_K0Inst_LFInst_13_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_13_LFInst_1_U4  ( .A(
        \Red_K0Inst_LFInst_13_LFInst_1_n2 ), .B(Key[182]), .ZN(Red_K0[53]) );
  XNOR2_X1 \Red_K0Inst_LFInst_13_LFInst_1_U3  ( .A(Key[183]), .B(Key[180]), 
        .ZN(\Red_K0Inst_LFInst_13_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_13_LFInst_2_U4  ( .A(
        \Red_K0Inst_LFInst_13_LFInst_2_n2 ), .B(Key[181]), .ZN(Red_K0[54]) );
  XNOR2_X1 \Red_K0Inst_LFInst_13_LFInst_2_U3  ( .A(Key[183]), .B(Key[180]), 
        .ZN(\Red_K0Inst_LFInst_13_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_13_LFInst_3_U4  ( .A(
        \Red_K0Inst_LFInst_13_LFInst_3_n2 ), .B(Key[181]), .ZN(Red_K0[55]) );
  XNOR2_X1 \Red_K0Inst_LFInst_13_LFInst_3_U3  ( .A(Key[182]), .B(Key[180]), 
        .ZN(\Red_K0Inst_LFInst_13_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_14_LFInst_0_U4  ( .A(
        \Red_K0Inst_LFInst_14_LFInst_0_n2 ), .B(Key[186]), .ZN(Red_K0[56]) );
  XNOR2_X1 \Red_K0Inst_LFInst_14_LFInst_0_U3  ( .A(Key[187]), .B(Key[185]), 
        .ZN(\Red_K0Inst_LFInst_14_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_14_LFInst_1_U4  ( .A(
        \Red_K0Inst_LFInst_14_LFInst_1_n2 ), .B(Key[186]), .ZN(Red_K0[57]) );
  XNOR2_X1 \Red_K0Inst_LFInst_14_LFInst_1_U3  ( .A(Key[187]), .B(Key[184]), 
        .ZN(\Red_K0Inst_LFInst_14_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_14_LFInst_2_U4  ( .A(
        \Red_K0Inst_LFInst_14_LFInst_2_n2 ), .B(Key[185]), .ZN(Red_K0[58]) );
  XNOR2_X1 \Red_K0Inst_LFInst_14_LFInst_2_U3  ( .A(Key[187]), .B(Key[184]), 
        .ZN(\Red_K0Inst_LFInst_14_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_14_LFInst_3_U4  ( .A(
        \Red_K0Inst_LFInst_14_LFInst_3_n2 ), .B(Key[185]), .ZN(Red_K0[59]) );
  XNOR2_X1 \Red_K0Inst_LFInst_14_LFInst_3_U3  ( .A(Key[186]), .B(Key[184]), 
        .ZN(\Red_K0Inst_LFInst_14_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_15_LFInst_0_U4  ( .A(
        \Red_K0Inst_LFInst_15_LFInst_0_n2 ), .B(Key[190]), .ZN(Red_K0[60]) );
  XNOR2_X1 \Red_K0Inst_LFInst_15_LFInst_0_U3  ( .A(Key[191]), .B(Key[189]), 
        .ZN(\Red_K0Inst_LFInst_15_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_15_LFInst_1_U4  ( .A(
        \Red_K0Inst_LFInst_15_LFInst_1_n2 ), .B(Key[190]), .ZN(Red_K0[61]) );
  XNOR2_X1 \Red_K0Inst_LFInst_15_LFInst_1_U3  ( .A(Key[191]), .B(Key[188]), 
        .ZN(\Red_K0Inst_LFInst_15_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_15_LFInst_2_U4  ( .A(
        \Red_K0Inst_LFInst_15_LFInst_2_n2 ), .B(Key[189]), .ZN(Red_K0[62]) );
  XNOR2_X1 \Red_K0Inst_LFInst_15_LFInst_2_U3  ( .A(Key[191]), .B(Key[188]), 
        .ZN(\Red_K0Inst_LFInst_15_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K0Inst_LFInst_15_LFInst_3_U4  ( .A(
        \Red_K0Inst_LFInst_15_LFInst_3_n2 ), .B(Key[189]), .ZN(Red_K0[63]) );
  XNOR2_X1 \Red_K0Inst_LFInst_15_LFInst_3_U3  ( .A(Key[190]), .B(Key[188]), 
        .ZN(\Red_K0Inst_LFInst_15_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_0_LFInst_0_U4  ( .A(
        \Red_K1Inst_LFInst_0_LFInst_0_n2 ), .B(Key[66]), .ZN(Red_K1[0]) );
  XNOR2_X1 \Red_K1Inst_LFInst_0_LFInst_0_U3  ( .A(Key[67]), .B(Key[65]), .ZN(
        \Red_K1Inst_LFInst_0_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_0_LFInst_1_U4  ( .A(
        \Red_K1Inst_LFInst_0_LFInst_1_n2 ), .B(Key[66]), .ZN(Red_K1[1]) );
  XNOR2_X1 \Red_K1Inst_LFInst_0_LFInst_1_U3  ( .A(Key[67]), .B(Key[64]), .ZN(
        \Red_K1Inst_LFInst_0_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_0_LFInst_2_U4  ( .A(
        \Red_K1Inst_LFInst_0_LFInst_2_n2 ), .B(Key[65]), .ZN(Red_K1[2]) );
  XNOR2_X1 \Red_K1Inst_LFInst_0_LFInst_2_U3  ( .A(Key[67]), .B(Key[64]), .ZN(
        \Red_K1Inst_LFInst_0_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_0_LFInst_3_U4  ( .A(
        \Red_K1Inst_LFInst_0_LFInst_3_n2 ), .B(Key[65]), .ZN(Red_K1[3]) );
  XNOR2_X1 \Red_K1Inst_LFInst_0_LFInst_3_U3  ( .A(Key[66]), .B(Key[64]), .ZN(
        \Red_K1Inst_LFInst_0_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_1_LFInst_0_U4  ( .A(
        \Red_K1Inst_LFInst_1_LFInst_0_n2 ), .B(Key[70]), .ZN(Red_K1[4]) );
  XNOR2_X1 \Red_K1Inst_LFInst_1_LFInst_0_U3  ( .A(Key[71]), .B(Key[69]), .ZN(
        \Red_K1Inst_LFInst_1_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_1_LFInst_1_U4  ( .A(
        \Red_K1Inst_LFInst_1_LFInst_1_n2 ), .B(Key[70]), .ZN(Red_K1[5]) );
  XNOR2_X1 \Red_K1Inst_LFInst_1_LFInst_1_U3  ( .A(Key[71]), .B(Key[68]), .ZN(
        \Red_K1Inst_LFInst_1_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_1_LFInst_2_U4  ( .A(
        \Red_K1Inst_LFInst_1_LFInst_2_n2 ), .B(Key[69]), .ZN(Red_K1[6]) );
  XNOR2_X1 \Red_K1Inst_LFInst_1_LFInst_2_U3  ( .A(Key[71]), .B(Key[68]), .ZN(
        \Red_K1Inst_LFInst_1_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_1_LFInst_3_U4  ( .A(
        \Red_K1Inst_LFInst_1_LFInst_3_n2 ), .B(Key[69]), .ZN(Red_K1[7]) );
  XNOR2_X1 \Red_K1Inst_LFInst_1_LFInst_3_U3  ( .A(Key[70]), .B(Key[68]), .ZN(
        \Red_K1Inst_LFInst_1_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_2_LFInst_0_U4  ( .A(
        \Red_K1Inst_LFInst_2_LFInst_0_n2 ), .B(Key[74]), .ZN(Red_K1[8]) );
  XNOR2_X1 \Red_K1Inst_LFInst_2_LFInst_0_U3  ( .A(Key[75]), .B(Key[73]), .ZN(
        \Red_K1Inst_LFInst_2_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_2_LFInst_1_U4  ( .A(
        \Red_K1Inst_LFInst_2_LFInst_1_n2 ), .B(Key[74]), .ZN(Red_K1[9]) );
  XNOR2_X1 \Red_K1Inst_LFInst_2_LFInst_1_U3  ( .A(Key[75]), .B(Key[72]), .ZN(
        \Red_K1Inst_LFInst_2_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_2_LFInst_2_U4  ( .A(
        \Red_K1Inst_LFInst_2_LFInst_2_n2 ), .B(Key[73]), .ZN(Red_K1[10]) );
  XNOR2_X1 \Red_K1Inst_LFInst_2_LFInst_2_U3  ( .A(Key[75]), .B(Key[72]), .ZN(
        \Red_K1Inst_LFInst_2_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_2_LFInst_3_U4  ( .A(
        \Red_K1Inst_LFInst_2_LFInst_3_n2 ), .B(Key[73]), .ZN(Red_K1[11]) );
  XNOR2_X1 \Red_K1Inst_LFInst_2_LFInst_3_U3  ( .A(Key[74]), .B(Key[72]), .ZN(
        \Red_K1Inst_LFInst_2_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_3_LFInst_0_U4  ( .A(
        \Red_K1Inst_LFInst_3_LFInst_0_n2 ), .B(Key[78]), .ZN(Red_K1[12]) );
  XNOR2_X1 \Red_K1Inst_LFInst_3_LFInst_0_U3  ( .A(Key[79]), .B(Key[77]), .ZN(
        \Red_K1Inst_LFInst_3_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_3_LFInst_1_U4  ( .A(
        \Red_K1Inst_LFInst_3_LFInst_1_n2 ), .B(Key[78]), .ZN(Red_K1[13]) );
  XNOR2_X1 \Red_K1Inst_LFInst_3_LFInst_1_U3  ( .A(Key[79]), .B(Key[76]), .ZN(
        \Red_K1Inst_LFInst_3_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_3_LFInst_2_U4  ( .A(
        \Red_K1Inst_LFInst_3_LFInst_2_n2 ), .B(Key[77]), .ZN(Red_K1[14]) );
  XNOR2_X1 \Red_K1Inst_LFInst_3_LFInst_2_U3  ( .A(Key[79]), .B(Key[76]), .ZN(
        \Red_K1Inst_LFInst_3_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_3_LFInst_3_U4  ( .A(
        \Red_K1Inst_LFInst_3_LFInst_3_n2 ), .B(Key[77]), .ZN(Red_K1[15]) );
  XNOR2_X1 \Red_K1Inst_LFInst_3_LFInst_3_U3  ( .A(Key[78]), .B(Key[76]), .ZN(
        \Red_K1Inst_LFInst_3_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_4_LFInst_0_U4  ( .A(
        \Red_K1Inst_LFInst_4_LFInst_0_n2 ), .B(Key[82]), .ZN(Red_K1[16]) );
  XNOR2_X1 \Red_K1Inst_LFInst_4_LFInst_0_U3  ( .A(Key[83]), .B(Key[81]), .ZN(
        \Red_K1Inst_LFInst_4_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_4_LFInst_1_U4  ( .A(
        \Red_K1Inst_LFInst_4_LFInst_1_n2 ), .B(Key[82]), .ZN(Red_K1[17]) );
  XNOR2_X1 \Red_K1Inst_LFInst_4_LFInst_1_U3  ( .A(Key[83]), .B(Key[80]), .ZN(
        \Red_K1Inst_LFInst_4_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_4_LFInst_2_U4  ( .A(
        \Red_K1Inst_LFInst_4_LFInst_2_n2 ), .B(Key[81]), .ZN(Red_K1[18]) );
  XNOR2_X1 \Red_K1Inst_LFInst_4_LFInst_2_U3  ( .A(Key[83]), .B(Key[80]), .ZN(
        \Red_K1Inst_LFInst_4_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_4_LFInst_3_U4  ( .A(
        \Red_K1Inst_LFInst_4_LFInst_3_n2 ), .B(Key[81]), .ZN(Red_K1[19]) );
  XNOR2_X1 \Red_K1Inst_LFInst_4_LFInst_3_U3  ( .A(Key[82]), .B(Key[80]), .ZN(
        \Red_K1Inst_LFInst_4_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_5_LFInst_0_U4  ( .A(
        \Red_K1Inst_LFInst_5_LFInst_0_n2 ), .B(Key[86]), .ZN(Red_K1[20]) );
  XNOR2_X1 \Red_K1Inst_LFInst_5_LFInst_0_U3  ( .A(Key[87]), .B(Key[85]), .ZN(
        \Red_K1Inst_LFInst_5_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_5_LFInst_1_U4  ( .A(
        \Red_K1Inst_LFInst_5_LFInst_1_n2 ), .B(Key[86]), .ZN(Red_K1[21]) );
  XNOR2_X1 \Red_K1Inst_LFInst_5_LFInst_1_U3  ( .A(Key[87]), .B(Key[84]), .ZN(
        \Red_K1Inst_LFInst_5_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_5_LFInst_2_U4  ( .A(
        \Red_K1Inst_LFInst_5_LFInst_2_n2 ), .B(Key[85]), .ZN(Red_K1[22]) );
  XNOR2_X1 \Red_K1Inst_LFInst_5_LFInst_2_U3  ( .A(Key[87]), .B(Key[84]), .ZN(
        \Red_K1Inst_LFInst_5_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_5_LFInst_3_U4  ( .A(
        \Red_K1Inst_LFInst_5_LFInst_3_n2 ), .B(Key[85]), .ZN(Red_K1[23]) );
  XNOR2_X1 \Red_K1Inst_LFInst_5_LFInst_3_U3  ( .A(Key[86]), .B(Key[84]), .ZN(
        \Red_K1Inst_LFInst_5_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_6_LFInst_0_U4  ( .A(
        \Red_K1Inst_LFInst_6_LFInst_0_n2 ), .B(Key[90]), .ZN(Red_K1[24]) );
  XNOR2_X1 \Red_K1Inst_LFInst_6_LFInst_0_U3  ( .A(Key[91]), .B(Key[89]), .ZN(
        \Red_K1Inst_LFInst_6_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_6_LFInst_1_U4  ( .A(
        \Red_K1Inst_LFInst_6_LFInst_1_n2 ), .B(Key[90]), .ZN(Red_K1[25]) );
  XNOR2_X1 \Red_K1Inst_LFInst_6_LFInst_1_U3  ( .A(Key[91]), .B(Key[88]), .ZN(
        \Red_K1Inst_LFInst_6_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_6_LFInst_2_U4  ( .A(
        \Red_K1Inst_LFInst_6_LFInst_2_n2 ), .B(Key[89]), .ZN(Red_K1[26]) );
  XNOR2_X1 \Red_K1Inst_LFInst_6_LFInst_2_U3  ( .A(Key[91]), .B(Key[88]), .ZN(
        \Red_K1Inst_LFInst_6_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_6_LFInst_3_U4  ( .A(
        \Red_K1Inst_LFInst_6_LFInst_3_n2 ), .B(Key[89]), .ZN(Red_K1[27]) );
  XNOR2_X1 \Red_K1Inst_LFInst_6_LFInst_3_U3  ( .A(Key[90]), .B(Key[88]), .ZN(
        \Red_K1Inst_LFInst_6_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_7_LFInst_0_U4  ( .A(
        \Red_K1Inst_LFInst_7_LFInst_0_n2 ), .B(Key[94]), .ZN(Red_K1[28]) );
  XNOR2_X1 \Red_K1Inst_LFInst_7_LFInst_0_U3  ( .A(Key[95]), .B(Key[93]), .ZN(
        \Red_K1Inst_LFInst_7_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_7_LFInst_1_U4  ( .A(
        \Red_K1Inst_LFInst_7_LFInst_1_n2 ), .B(Key[94]), .ZN(Red_K1[29]) );
  XNOR2_X1 \Red_K1Inst_LFInst_7_LFInst_1_U3  ( .A(Key[95]), .B(Key[92]), .ZN(
        \Red_K1Inst_LFInst_7_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_7_LFInst_2_U4  ( .A(
        \Red_K1Inst_LFInst_7_LFInst_2_n2 ), .B(Key[93]), .ZN(Red_K1[30]) );
  XNOR2_X1 \Red_K1Inst_LFInst_7_LFInst_2_U3  ( .A(Key[95]), .B(Key[92]), .ZN(
        \Red_K1Inst_LFInst_7_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_7_LFInst_3_U4  ( .A(
        \Red_K1Inst_LFInst_7_LFInst_3_n2 ), .B(Key[93]), .ZN(Red_K1[31]) );
  XNOR2_X1 \Red_K1Inst_LFInst_7_LFInst_3_U3  ( .A(Key[94]), .B(Key[92]), .ZN(
        \Red_K1Inst_LFInst_7_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_8_LFInst_0_U4  ( .A(
        \Red_K1Inst_LFInst_8_LFInst_0_n2 ), .B(Key[98]), .ZN(Red_K1[32]) );
  XNOR2_X1 \Red_K1Inst_LFInst_8_LFInst_0_U3  ( .A(Key[99]), .B(Key[97]), .ZN(
        \Red_K1Inst_LFInst_8_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_8_LFInst_1_U4  ( .A(
        \Red_K1Inst_LFInst_8_LFInst_1_n2 ), .B(Key[98]), .ZN(Red_K1[33]) );
  XNOR2_X1 \Red_K1Inst_LFInst_8_LFInst_1_U3  ( .A(Key[99]), .B(Key[96]), .ZN(
        \Red_K1Inst_LFInst_8_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_8_LFInst_2_U4  ( .A(
        \Red_K1Inst_LFInst_8_LFInst_2_n2 ), .B(Key[97]), .ZN(Red_K1[34]) );
  XNOR2_X1 \Red_K1Inst_LFInst_8_LFInst_2_U3  ( .A(Key[99]), .B(Key[96]), .ZN(
        \Red_K1Inst_LFInst_8_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_8_LFInst_3_U4  ( .A(
        \Red_K1Inst_LFInst_8_LFInst_3_n2 ), .B(Key[97]), .ZN(Red_K1[35]) );
  XNOR2_X1 \Red_K1Inst_LFInst_8_LFInst_3_U3  ( .A(Key[98]), .B(Key[96]), .ZN(
        \Red_K1Inst_LFInst_8_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_9_LFInst_0_U4  ( .A(
        \Red_K1Inst_LFInst_9_LFInst_0_n2 ), .B(Key[102]), .ZN(Red_K1[36]) );
  XNOR2_X1 \Red_K1Inst_LFInst_9_LFInst_0_U3  ( .A(Key[103]), .B(Key[101]), 
        .ZN(\Red_K1Inst_LFInst_9_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_9_LFInst_1_U4  ( .A(
        \Red_K1Inst_LFInst_9_LFInst_1_n2 ), .B(Key[102]), .ZN(Red_K1[37]) );
  XNOR2_X1 \Red_K1Inst_LFInst_9_LFInst_1_U3  ( .A(Key[103]), .B(Key[100]), 
        .ZN(\Red_K1Inst_LFInst_9_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_9_LFInst_2_U4  ( .A(
        \Red_K1Inst_LFInst_9_LFInst_2_n2 ), .B(Key[101]), .ZN(Red_K1[38]) );
  XNOR2_X1 \Red_K1Inst_LFInst_9_LFInst_2_U3  ( .A(Key[103]), .B(Key[100]), 
        .ZN(\Red_K1Inst_LFInst_9_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_9_LFInst_3_U4  ( .A(
        \Red_K1Inst_LFInst_9_LFInst_3_n2 ), .B(Key[101]), .ZN(Red_K1[39]) );
  XNOR2_X1 \Red_K1Inst_LFInst_9_LFInst_3_U3  ( .A(Key[102]), .B(Key[100]), 
        .ZN(\Red_K1Inst_LFInst_9_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_10_LFInst_0_U4  ( .A(
        \Red_K1Inst_LFInst_10_LFInst_0_n2 ), .B(Key[106]), .ZN(Red_K1[40]) );
  XNOR2_X1 \Red_K1Inst_LFInst_10_LFInst_0_U3  ( .A(Key[107]), .B(Key[105]), 
        .ZN(\Red_K1Inst_LFInst_10_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_10_LFInst_1_U4  ( .A(
        \Red_K1Inst_LFInst_10_LFInst_1_n2 ), .B(Key[106]), .ZN(Red_K1[41]) );
  XNOR2_X1 \Red_K1Inst_LFInst_10_LFInst_1_U3  ( .A(Key[107]), .B(Key[104]), 
        .ZN(\Red_K1Inst_LFInst_10_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_10_LFInst_2_U4  ( .A(
        \Red_K1Inst_LFInst_10_LFInst_2_n2 ), .B(Key[105]), .ZN(Red_K1[42]) );
  XNOR2_X1 \Red_K1Inst_LFInst_10_LFInst_2_U3  ( .A(Key[107]), .B(Key[104]), 
        .ZN(\Red_K1Inst_LFInst_10_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_10_LFInst_3_U4  ( .A(
        \Red_K1Inst_LFInst_10_LFInst_3_n2 ), .B(Key[105]), .ZN(Red_K1[43]) );
  XNOR2_X1 \Red_K1Inst_LFInst_10_LFInst_3_U3  ( .A(Key[106]), .B(Key[104]), 
        .ZN(\Red_K1Inst_LFInst_10_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_11_LFInst_0_U4  ( .A(
        \Red_K1Inst_LFInst_11_LFInst_0_n2 ), .B(Key[110]), .ZN(Red_K1[44]) );
  XNOR2_X1 \Red_K1Inst_LFInst_11_LFInst_0_U3  ( .A(Key[111]), .B(Key[109]), 
        .ZN(\Red_K1Inst_LFInst_11_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_11_LFInst_1_U4  ( .A(
        \Red_K1Inst_LFInst_11_LFInst_1_n2 ), .B(Key[110]), .ZN(Red_K1[45]) );
  XNOR2_X1 \Red_K1Inst_LFInst_11_LFInst_1_U3  ( .A(Key[111]), .B(Key[108]), 
        .ZN(\Red_K1Inst_LFInst_11_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_11_LFInst_2_U4  ( .A(
        \Red_K1Inst_LFInst_11_LFInst_2_n2 ), .B(Key[109]), .ZN(Red_K1[46]) );
  XNOR2_X1 \Red_K1Inst_LFInst_11_LFInst_2_U3  ( .A(Key[111]), .B(Key[108]), 
        .ZN(\Red_K1Inst_LFInst_11_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_11_LFInst_3_U4  ( .A(
        \Red_K1Inst_LFInst_11_LFInst_3_n2 ), .B(Key[109]), .ZN(Red_K1[47]) );
  XNOR2_X1 \Red_K1Inst_LFInst_11_LFInst_3_U3  ( .A(Key[110]), .B(Key[108]), 
        .ZN(\Red_K1Inst_LFInst_11_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_12_LFInst_0_U4  ( .A(
        \Red_K1Inst_LFInst_12_LFInst_0_n2 ), .B(Key[114]), .ZN(Red_K1[48]) );
  XNOR2_X1 \Red_K1Inst_LFInst_12_LFInst_0_U3  ( .A(Key[115]), .B(Key[113]), 
        .ZN(\Red_K1Inst_LFInst_12_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_12_LFInst_1_U4  ( .A(
        \Red_K1Inst_LFInst_12_LFInst_1_n2 ), .B(Key[114]), .ZN(Red_K1[49]) );
  XNOR2_X1 \Red_K1Inst_LFInst_12_LFInst_1_U3  ( .A(Key[115]), .B(Key[112]), 
        .ZN(\Red_K1Inst_LFInst_12_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_12_LFInst_2_U4  ( .A(
        \Red_K1Inst_LFInst_12_LFInst_2_n2 ), .B(Key[113]), .ZN(Red_K1[50]) );
  XNOR2_X1 \Red_K1Inst_LFInst_12_LFInst_2_U3  ( .A(Key[115]), .B(Key[112]), 
        .ZN(\Red_K1Inst_LFInst_12_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_12_LFInst_3_U4  ( .A(
        \Red_K1Inst_LFInst_12_LFInst_3_n2 ), .B(Key[113]), .ZN(Red_K1[51]) );
  XNOR2_X1 \Red_K1Inst_LFInst_12_LFInst_3_U3  ( .A(Key[114]), .B(Key[112]), 
        .ZN(\Red_K1Inst_LFInst_12_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_13_LFInst_0_U4  ( .A(
        \Red_K1Inst_LFInst_13_LFInst_0_n2 ), .B(Key[118]), .ZN(Red_K1[52]) );
  XNOR2_X1 \Red_K1Inst_LFInst_13_LFInst_0_U3  ( .A(Key[119]), .B(Key[117]), 
        .ZN(\Red_K1Inst_LFInst_13_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_13_LFInst_1_U4  ( .A(
        \Red_K1Inst_LFInst_13_LFInst_1_n2 ), .B(Key[118]), .ZN(Red_K1[53]) );
  XNOR2_X1 \Red_K1Inst_LFInst_13_LFInst_1_U3  ( .A(Key[119]), .B(Key[116]), 
        .ZN(\Red_K1Inst_LFInst_13_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_13_LFInst_2_U4  ( .A(
        \Red_K1Inst_LFInst_13_LFInst_2_n2 ), .B(Key[117]), .ZN(Red_K1[54]) );
  XNOR2_X1 \Red_K1Inst_LFInst_13_LFInst_2_U3  ( .A(Key[119]), .B(Key[116]), 
        .ZN(\Red_K1Inst_LFInst_13_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_13_LFInst_3_U4  ( .A(
        \Red_K1Inst_LFInst_13_LFInst_3_n2 ), .B(Key[117]), .ZN(Red_K1[55]) );
  XNOR2_X1 \Red_K1Inst_LFInst_13_LFInst_3_U3  ( .A(Key[118]), .B(Key[116]), 
        .ZN(\Red_K1Inst_LFInst_13_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_14_LFInst_0_U4  ( .A(
        \Red_K1Inst_LFInst_14_LFInst_0_n2 ), .B(Key[122]), .ZN(Red_K1[56]) );
  XNOR2_X1 \Red_K1Inst_LFInst_14_LFInst_0_U3  ( .A(Key[123]), .B(Key[121]), 
        .ZN(\Red_K1Inst_LFInst_14_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_14_LFInst_1_U4  ( .A(
        \Red_K1Inst_LFInst_14_LFInst_1_n2 ), .B(Key[122]), .ZN(Red_K1[57]) );
  XNOR2_X1 \Red_K1Inst_LFInst_14_LFInst_1_U3  ( .A(Key[123]), .B(Key[120]), 
        .ZN(\Red_K1Inst_LFInst_14_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_14_LFInst_2_U4  ( .A(
        \Red_K1Inst_LFInst_14_LFInst_2_n2 ), .B(Key[121]), .ZN(Red_K1[58]) );
  XNOR2_X1 \Red_K1Inst_LFInst_14_LFInst_2_U3  ( .A(Key[123]), .B(Key[120]), 
        .ZN(\Red_K1Inst_LFInst_14_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_14_LFInst_3_U4  ( .A(
        \Red_K1Inst_LFInst_14_LFInst_3_n2 ), .B(Key[121]), .ZN(Red_K1[59]) );
  XNOR2_X1 \Red_K1Inst_LFInst_14_LFInst_3_U3  ( .A(Key[122]), .B(Key[120]), 
        .ZN(\Red_K1Inst_LFInst_14_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_15_LFInst_0_U4  ( .A(
        \Red_K1Inst_LFInst_15_LFInst_0_n2 ), .B(Key[126]), .ZN(Red_K1[60]) );
  XNOR2_X1 \Red_K1Inst_LFInst_15_LFInst_0_U3  ( .A(Key[127]), .B(Key[125]), 
        .ZN(\Red_K1Inst_LFInst_15_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_15_LFInst_1_U4  ( .A(
        \Red_K1Inst_LFInst_15_LFInst_1_n2 ), .B(Key[126]), .ZN(Red_K1[61]) );
  XNOR2_X1 \Red_K1Inst_LFInst_15_LFInst_1_U3  ( .A(Key[127]), .B(Key[124]), 
        .ZN(\Red_K1Inst_LFInst_15_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_15_LFInst_2_U4  ( .A(
        \Red_K1Inst_LFInst_15_LFInst_2_n2 ), .B(Key[125]), .ZN(Red_K1[62]) );
  XNOR2_X1 \Red_K1Inst_LFInst_15_LFInst_2_U3  ( .A(Key[127]), .B(Key[124]), 
        .ZN(\Red_K1Inst_LFInst_15_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K1Inst_LFInst_15_LFInst_3_U4  ( .A(
        \Red_K1Inst_LFInst_15_LFInst_3_n2 ), .B(Key[125]), .ZN(Red_K1[63]) );
  XNOR2_X1 \Red_K1Inst_LFInst_15_LFInst_3_U3  ( .A(Key[126]), .B(Key[124]), 
        .ZN(\Red_K1Inst_LFInst_15_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_0_LFInst_0_U4  ( .A(
        \Red_K2Inst_LFInst_0_LFInst_0_n2 ), .B(Key[2]), .ZN(Red_K2[0]) );
  XNOR2_X1 \Red_K2Inst_LFInst_0_LFInst_0_U3  ( .A(Key[3]), .B(Key[1]), .ZN(
        \Red_K2Inst_LFInst_0_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_0_LFInst_1_U4  ( .A(
        \Red_K2Inst_LFInst_0_LFInst_1_n2 ), .B(Key[2]), .ZN(Red_K2[1]) );
  XNOR2_X1 \Red_K2Inst_LFInst_0_LFInst_1_U3  ( .A(Key[3]), .B(Key[0]), .ZN(
        \Red_K2Inst_LFInst_0_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_0_LFInst_2_U4  ( .A(
        \Red_K2Inst_LFInst_0_LFInst_2_n2 ), .B(Key[1]), .ZN(Red_K2[2]) );
  XNOR2_X1 \Red_K2Inst_LFInst_0_LFInst_2_U3  ( .A(Key[3]), .B(Key[0]), .ZN(
        \Red_K2Inst_LFInst_0_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_0_LFInst_3_U4  ( .A(
        \Red_K2Inst_LFInst_0_LFInst_3_n2 ), .B(Key[1]), .ZN(Red_K2[3]) );
  XNOR2_X1 \Red_K2Inst_LFInst_0_LFInst_3_U3  ( .A(Key[2]), .B(Key[0]), .ZN(
        \Red_K2Inst_LFInst_0_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_1_LFInst_0_U4  ( .A(
        \Red_K2Inst_LFInst_1_LFInst_0_n2 ), .B(Key[6]), .ZN(Red_K2[4]) );
  XNOR2_X1 \Red_K2Inst_LFInst_1_LFInst_0_U3  ( .A(Key[7]), .B(Key[5]), .ZN(
        \Red_K2Inst_LFInst_1_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_1_LFInst_1_U4  ( .A(
        \Red_K2Inst_LFInst_1_LFInst_1_n2 ), .B(Key[6]), .ZN(Red_K2[5]) );
  XNOR2_X1 \Red_K2Inst_LFInst_1_LFInst_1_U3  ( .A(Key[7]), .B(Key[4]), .ZN(
        \Red_K2Inst_LFInst_1_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_1_LFInst_2_U4  ( .A(
        \Red_K2Inst_LFInst_1_LFInst_2_n2 ), .B(Key[5]), .ZN(Red_K2[6]) );
  XNOR2_X1 \Red_K2Inst_LFInst_1_LFInst_2_U3  ( .A(Key[7]), .B(Key[4]), .ZN(
        \Red_K2Inst_LFInst_1_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_1_LFInst_3_U4  ( .A(
        \Red_K2Inst_LFInst_1_LFInst_3_n2 ), .B(Key[5]), .ZN(Red_K2[7]) );
  XNOR2_X1 \Red_K2Inst_LFInst_1_LFInst_3_U3  ( .A(Key[6]), .B(Key[4]), .ZN(
        \Red_K2Inst_LFInst_1_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_2_LFInst_0_U4  ( .A(
        \Red_K2Inst_LFInst_2_LFInst_0_n2 ), .B(Key[10]), .ZN(Red_K2[8]) );
  XNOR2_X1 \Red_K2Inst_LFInst_2_LFInst_0_U3  ( .A(Key[11]), .B(Key[9]), .ZN(
        \Red_K2Inst_LFInst_2_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_2_LFInst_1_U4  ( .A(
        \Red_K2Inst_LFInst_2_LFInst_1_n2 ), .B(Key[10]), .ZN(Red_K2[9]) );
  XNOR2_X1 \Red_K2Inst_LFInst_2_LFInst_1_U3  ( .A(Key[11]), .B(Key[8]), .ZN(
        \Red_K2Inst_LFInst_2_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_2_LFInst_2_U4  ( .A(
        \Red_K2Inst_LFInst_2_LFInst_2_n2 ), .B(Key[9]), .ZN(Red_K2[10]) );
  XNOR2_X1 \Red_K2Inst_LFInst_2_LFInst_2_U3  ( .A(Key[11]), .B(Key[8]), .ZN(
        \Red_K2Inst_LFInst_2_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_2_LFInst_3_U4  ( .A(
        \Red_K2Inst_LFInst_2_LFInst_3_n2 ), .B(Key[9]), .ZN(Red_K2[11]) );
  XNOR2_X1 \Red_K2Inst_LFInst_2_LFInst_3_U3  ( .A(Key[10]), .B(Key[8]), .ZN(
        \Red_K2Inst_LFInst_2_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_3_LFInst_0_U4  ( .A(
        \Red_K2Inst_LFInst_3_LFInst_0_n2 ), .B(Key[14]), .ZN(Red_K2[12]) );
  XNOR2_X1 \Red_K2Inst_LFInst_3_LFInst_0_U3  ( .A(Key[15]), .B(Key[13]), .ZN(
        \Red_K2Inst_LFInst_3_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_3_LFInst_1_U4  ( .A(
        \Red_K2Inst_LFInst_3_LFInst_1_n2 ), .B(Key[14]), .ZN(Red_K2[13]) );
  XNOR2_X1 \Red_K2Inst_LFInst_3_LFInst_1_U3  ( .A(Key[15]), .B(Key[12]), .ZN(
        \Red_K2Inst_LFInst_3_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_3_LFInst_2_U4  ( .A(
        \Red_K2Inst_LFInst_3_LFInst_2_n2 ), .B(Key[13]), .ZN(Red_K2[14]) );
  XNOR2_X1 \Red_K2Inst_LFInst_3_LFInst_2_U3  ( .A(Key[15]), .B(Key[12]), .ZN(
        \Red_K2Inst_LFInst_3_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_3_LFInst_3_U4  ( .A(
        \Red_K2Inst_LFInst_3_LFInst_3_n2 ), .B(Key[13]), .ZN(Red_K2[15]) );
  XNOR2_X1 \Red_K2Inst_LFInst_3_LFInst_3_U3  ( .A(Key[14]), .B(Key[12]), .ZN(
        \Red_K2Inst_LFInst_3_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_4_LFInst_0_U4  ( .A(
        \Red_K2Inst_LFInst_4_LFInst_0_n2 ), .B(Key[18]), .ZN(Red_K2[16]) );
  XNOR2_X1 \Red_K2Inst_LFInst_4_LFInst_0_U3  ( .A(Key[19]), .B(Key[17]), .ZN(
        \Red_K2Inst_LFInst_4_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_4_LFInst_1_U4  ( .A(
        \Red_K2Inst_LFInst_4_LFInst_1_n2 ), .B(Key[18]), .ZN(Red_K2[17]) );
  XNOR2_X1 \Red_K2Inst_LFInst_4_LFInst_1_U3  ( .A(Key[19]), .B(Key[16]), .ZN(
        \Red_K2Inst_LFInst_4_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_4_LFInst_2_U4  ( .A(
        \Red_K2Inst_LFInst_4_LFInst_2_n2 ), .B(Key[17]), .ZN(Red_K2[18]) );
  XNOR2_X1 \Red_K2Inst_LFInst_4_LFInst_2_U3  ( .A(Key[19]), .B(Key[16]), .ZN(
        \Red_K2Inst_LFInst_4_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_4_LFInst_3_U4  ( .A(
        \Red_K2Inst_LFInst_4_LFInst_3_n2 ), .B(Key[17]), .ZN(Red_K2[19]) );
  XNOR2_X1 \Red_K2Inst_LFInst_4_LFInst_3_U3  ( .A(Key[18]), .B(Key[16]), .ZN(
        \Red_K2Inst_LFInst_4_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_5_LFInst_0_U4  ( .A(
        \Red_K2Inst_LFInst_5_LFInst_0_n2 ), .B(Key[22]), .ZN(Red_K2[20]) );
  XNOR2_X1 \Red_K2Inst_LFInst_5_LFInst_0_U3  ( .A(Key[23]), .B(Key[21]), .ZN(
        \Red_K2Inst_LFInst_5_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_5_LFInst_1_U4  ( .A(
        \Red_K2Inst_LFInst_5_LFInst_1_n2 ), .B(Key[22]), .ZN(Red_K2[21]) );
  XNOR2_X1 \Red_K2Inst_LFInst_5_LFInst_1_U3  ( .A(Key[23]), .B(Key[20]), .ZN(
        \Red_K2Inst_LFInst_5_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_5_LFInst_2_U4  ( .A(
        \Red_K2Inst_LFInst_5_LFInst_2_n2 ), .B(Key[21]), .ZN(Red_K2[22]) );
  XNOR2_X1 \Red_K2Inst_LFInst_5_LFInst_2_U3  ( .A(Key[23]), .B(Key[20]), .ZN(
        \Red_K2Inst_LFInst_5_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_5_LFInst_3_U4  ( .A(
        \Red_K2Inst_LFInst_5_LFInst_3_n2 ), .B(Key[21]), .ZN(Red_K2[23]) );
  XNOR2_X1 \Red_K2Inst_LFInst_5_LFInst_3_U3  ( .A(Key[22]), .B(Key[20]), .ZN(
        \Red_K2Inst_LFInst_5_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_6_LFInst_0_U4  ( .A(
        \Red_K2Inst_LFInst_6_LFInst_0_n2 ), .B(Key[26]), .ZN(Red_K2[24]) );
  XNOR2_X1 \Red_K2Inst_LFInst_6_LFInst_0_U3  ( .A(Key[27]), .B(Key[25]), .ZN(
        \Red_K2Inst_LFInst_6_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_6_LFInst_1_U4  ( .A(
        \Red_K2Inst_LFInst_6_LFInst_1_n2 ), .B(Key[26]), .ZN(Red_K2[25]) );
  XNOR2_X1 \Red_K2Inst_LFInst_6_LFInst_1_U3  ( .A(Key[27]), .B(Key[24]), .ZN(
        \Red_K2Inst_LFInst_6_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_6_LFInst_2_U4  ( .A(
        \Red_K2Inst_LFInst_6_LFInst_2_n2 ), .B(Key[25]), .ZN(Red_K2[26]) );
  XNOR2_X1 \Red_K2Inst_LFInst_6_LFInst_2_U3  ( .A(Key[27]), .B(Key[24]), .ZN(
        \Red_K2Inst_LFInst_6_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_6_LFInst_3_U4  ( .A(
        \Red_K2Inst_LFInst_6_LFInst_3_n2 ), .B(Key[25]), .ZN(Red_K2[27]) );
  XNOR2_X1 \Red_K2Inst_LFInst_6_LFInst_3_U3  ( .A(Key[26]), .B(Key[24]), .ZN(
        \Red_K2Inst_LFInst_6_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_7_LFInst_0_U4  ( .A(
        \Red_K2Inst_LFInst_7_LFInst_0_n2 ), .B(Key[30]), .ZN(Red_K2[28]) );
  XNOR2_X1 \Red_K2Inst_LFInst_7_LFInst_0_U3  ( .A(Key[31]), .B(Key[29]), .ZN(
        \Red_K2Inst_LFInst_7_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_7_LFInst_1_U4  ( .A(
        \Red_K2Inst_LFInst_7_LFInst_1_n2 ), .B(Key[30]), .ZN(Red_K2[29]) );
  XNOR2_X1 \Red_K2Inst_LFInst_7_LFInst_1_U3  ( .A(Key[31]), .B(Key[28]), .ZN(
        \Red_K2Inst_LFInst_7_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_7_LFInst_2_U4  ( .A(
        \Red_K2Inst_LFInst_7_LFInst_2_n2 ), .B(Key[29]), .ZN(Red_K2[30]) );
  XNOR2_X1 \Red_K2Inst_LFInst_7_LFInst_2_U3  ( .A(Key[31]), .B(Key[28]), .ZN(
        \Red_K2Inst_LFInst_7_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_7_LFInst_3_U4  ( .A(
        \Red_K2Inst_LFInst_7_LFInst_3_n2 ), .B(Key[29]), .ZN(Red_K2[31]) );
  XNOR2_X1 \Red_K2Inst_LFInst_7_LFInst_3_U3  ( .A(Key[30]), .B(Key[28]), .ZN(
        \Red_K2Inst_LFInst_7_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_8_LFInst_0_U4  ( .A(
        \Red_K2Inst_LFInst_8_LFInst_0_n2 ), .B(Key[34]), .ZN(Red_K2[32]) );
  XNOR2_X1 \Red_K2Inst_LFInst_8_LFInst_0_U3  ( .A(Key[35]), .B(Key[33]), .ZN(
        \Red_K2Inst_LFInst_8_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_8_LFInst_1_U4  ( .A(
        \Red_K2Inst_LFInst_8_LFInst_1_n2 ), .B(Key[34]), .ZN(Red_K2[33]) );
  XNOR2_X1 \Red_K2Inst_LFInst_8_LFInst_1_U3  ( .A(Key[35]), .B(Key[32]), .ZN(
        \Red_K2Inst_LFInst_8_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_8_LFInst_2_U4  ( .A(
        \Red_K2Inst_LFInst_8_LFInst_2_n2 ), .B(Key[33]), .ZN(Red_K2[34]) );
  XNOR2_X1 \Red_K2Inst_LFInst_8_LFInst_2_U3  ( .A(Key[35]), .B(Key[32]), .ZN(
        \Red_K2Inst_LFInst_8_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_8_LFInst_3_U4  ( .A(
        \Red_K2Inst_LFInst_8_LFInst_3_n2 ), .B(Key[33]), .ZN(Red_K2[35]) );
  XNOR2_X1 \Red_K2Inst_LFInst_8_LFInst_3_U3  ( .A(Key[34]), .B(Key[32]), .ZN(
        \Red_K2Inst_LFInst_8_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_9_LFInst_0_U4  ( .A(
        \Red_K2Inst_LFInst_9_LFInst_0_n2 ), .B(Key[38]), .ZN(Red_K2[36]) );
  XNOR2_X1 \Red_K2Inst_LFInst_9_LFInst_0_U3  ( .A(Key[39]), .B(Key[37]), .ZN(
        \Red_K2Inst_LFInst_9_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_9_LFInst_1_U4  ( .A(
        \Red_K2Inst_LFInst_9_LFInst_1_n2 ), .B(Key[38]), .ZN(Red_K2[37]) );
  XNOR2_X1 \Red_K2Inst_LFInst_9_LFInst_1_U3  ( .A(Key[39]), .B(Key[36]), .ZN(
        \Red_K2Inst_LFInst_9_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_9_LFInst_2_U4  ( .A(
        \Red_K2Inst_LFInst_9_LFInst_2_n2 ), .B(Key[37]), .ZN(Red_K2[38]) );
  XNOR2_X1 \Red_K2Inst_LFInst_9_LFInst_2_U3  ( .A(Key[39]), .B(Key[36]), .ZN(
        \Red_K2Inst_LFInst_9_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_9_LFInst_3_U4  ( .A(
        \Red_K2Inst_LFInst_9_LFInst_3_n2 ), .B(Key[37]), .ZN(Red_K2[39]) );
  XNOR2_X1 \Red_K2Inst_LFInst_9_LFInst_3_U3  ( .A(Key[38]), .B(Key[36]), .ZN(
        \Red_K2Inst_LFInst_9_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_10_LFInst_0_U4  ( .A(
        \Red_K2Inst_LFInst_10_LFInst_0_n2 ), .B(Key[42]), .ZN(Red_K2[40]) );
  XNOR2_X1 \Red_K2Inst_LFInst_10_LFInst_0_U3  ( .A(Key[43]), .B(Key[41]), .ZN(
        \Red_K2Inst_LFInst_10_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_10_LFInst_1_U4  ( .A(
        \Red_K2Inst_LFInst_10_LFInst_1_n2 ), .B(Key[42]), .ZN(Red_K2[41]) );
  XNOR2_X1 \Red_K2Inst_LFInst_10_LFInst_1_U3  ( .A(Key[43]), .B(Key[40]), .ZN(
        \Red_K2Inst_LFInst_10_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_10_LFInst_2_U4  ( .A(
        \Red_K2Inst_LFInst_10_LFInst_2_n2 ), .B(Key[41]), .ZN(Red_K2[42]) );
  XNOR2_X1 \Red_K2Inst_LFInst_10_LFInst_2_U3  ( .A(Key[43]), .B(Key[40]), .ZN(
        \Red_K2Inst_LFInst_10_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_10_LFInst_3_U4  ( .A(
        \Red_K2Inst_LFInst_10_LFInst_3_n2 ), .B(Key[41]), .ZN(Red_K2[43]) );
  XNOR2_X1 \Red_K2Inst_LFInst_10_LFInst_3_U3  ( .A(Key[42]), .B(Key[40]), .ZN(
        \Red_K2Inst_LFInst_10_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_11_LFInst_0_U4  ( .A(
        \Red_K2Inst_LFInst_11_LFInst_0_n2 ), .B(Key[46]), .ZN(Red_K2[44]) );
  XNOR2_X1 \Red_K2Inst_LFInst_11_LFInst_0_U3  ( .A(Key[47]), .B(Key[45]), .ZN(
        \Red_K2Inst_LFInst_11_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_11_LFInst_1_U4  ( .A(
        \Red_K2Inst_LFInst_11_LFInst_1_n2 ), .B(Key[46]), .ZN(Red_K2[45]) );
  XNOR2_X1 \Red_K2Inst_LFInst_11_LFInst_1_U3  ( .A(Key[47]), .B(Key[44]), .ZN(
        \Red_K2Inst_LFInst_11_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_11_LFInst_2_U4  ( .A(
        \Red_K2Inst_LFInst_11_LFInst_2_n2 ), .B(Key[45]), .ZN(Red_K2[46]) );
  XNOR2_X1 \Red_K2Inst_LFInst_11_LFInst_2_U3  ( .A(Key[47]), .B(Key[44]), .ZN(
        \Red_K2Inst_LFInst_11_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_11_LFInst_3_U4  ( .A(
        \Red_K2Inst_LFInst_11_LFInst_3_n2 ), .B(Key[45]), .ZN(Red_K2[47]) );
  XNOR2_X1 \Red_K2Inst_LFInst_11_LFInst_3_U3  ( .A(Key[46]), .B(Key[44]), .ZN(
        \Red_K2Inst_LFInst_11_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_12_LFInst_0_U4  ( .A(
        \Red_K2Inst_LFInst_12_LFInst_0_n2 ), .B(Key[50]), .ZN(Red_K2[48]) );
  XNOR2_X1 \Red_K2Inst_LFInst_12_LFInst_0_U3  ( .A(Key[51]), .B(Key[49]), .ZN(
        \Red_K2Inst_LFInst_12_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_12_LFInst_1_U4  ( .A(
        \Red_K2Inst_LFInst_12_LFInst_1_n2 ), .B(Key[50]), .ZN(Red_K2[49]) );
  XNOR2_X1 \Red_K2Inst_LFInst_12_LFInst_1_U3  ( .A(Key[51]), .B(Key[48]), .ZN(
        \Red_K2Inst_LFInst_12_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_12_LFInst_2_U4  ( .A(
        \Red_K2Inst_LFInst_12_LFInst_2_n2 ), .B(Key[49]), .ZN(Red_K2[50]) );
  XNOR2_X1 \Red_K2Inst_LFInst_12_LFInst_2_U3  ( .A(Key[51]), .B(Key[48]), .ZN(
        \Red_K2Inst_LFInst_12_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_12_LFInst_3_U4  ( .A(
        \Red_K2Inst_LFInst_12_LFInst_3_n2 ), .B(Key[49]), .ZN(Red_K2[51]) );
  XNOR2_X1 \Red_K2Inst_LFInst_12_LFInst_3_U3  ( .A(Key[50]), .B(Key[48]), .ZN(
        \Red_K2Inst_LFInst_12_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_13_LFInst_0_U4  ( .A(
        \Red_K2Inst_LFInst_13_LFInst_0_n2 ), .B(Key[54]), .ZN(Red_K2[52]) );
  XNOR2_X1 \Red_K2Inst_LFInst_13_LFInst_0_U3  ( .A(Key[55]), .B(Key[53]), .ZN(
        \Red_K2Inst_LFInst_13_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_13_LFInst_1_U4  ( .A(
        \Red_K2Inst_LFInst_13_LFInst_1_n2 ), .B(Key[54]), .ZN(Red_K2[53]) );
  XNOR2_X1 \Red_K2Inst_LFInst_13_LFInst_1_U3  ( .A(Key[55]), .B(Key[52]), .ZN(
        \Red_K2Inst_LFInst_13_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_13_LFInst_2_U4  ( .A(
        \Red_K2Inst_LFInst_13_LFInst_2_n2 ), .B(Key[53]), .ZN(Red_K2[54]) );
  XNOR2_X1 \Red_K2Inst_LFInst_13_LFInst_2_U3  ( .A(Key[55]), .B(Key[52]), .ZN(
        \Red_K2Inst_LFInst_13_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_13_LFInst_3_U4  ( .A(
        \Red_K2Inst_LFInst_13_LFInst_3_n2 ), .B(Key[53]), .ZN(Red_K2[55]) );
  XNOR2_X1 \Red_K2Inst_LFInst_13_LFInst_3_U3  ( .A(Key[54]), .B(Key[52]), .ZN(
        \Red_K2Inst_LFInst_13_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_14_LFInst_0_U4  ( .A(
        \Red_K2Inst_LFInst_14_LFInst_0_n2 ), .B(Key[58]), .ZN(Red_K2[56]) );
  XNOR2_X1 \Red_K2Inst_LFInst_14_LFInst_0_U3  ( .A(Key[59]), .B(Key[57]), .ZN(
        \Red_K2Inst_LFInst_14_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_14_LFInst_1_U4  ( .A(
        \Red_K2Inst_LFInst_14_LFInst_1_n2 ), .B(Key[58]), .ZN(Red_K2[57]) );
  XNOR2_X1 \Red_K2Inst_LFInst_14_LFInst_1_U3  ( .A(Key[59]), .B(Key[56]), .ZN(
        \Red_K2Inst_LFInst_14_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_14_LFInst_2_U4  ( .A(
        \Red_K2Inst_LFInst_14_LFInst_2_n2 ), .B(Key[57]), .ZN(Red_K2[58]) );
  XNOR2_X1 \Red_K2Inst_LFInst_14_LFInst_2_U3  ( .A(Key[59]), .B(Key[56]), .ZN(
        \Red_K2Inst_LFInst_14_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_14_LFInst_3_U4  ( .A(
        \Red_K2Inst_LFInst_14_LFInst_3_n2 ), .B(Key[57]), .ZN(Red_K2[59]) );
  XNOR2_X1 \Red_K2Inst_LFInst_14_LFInst_3_U3  ( .A(Key[58]), .B(Key[56]), .ZN(
        \Red_K2Inst_LFInst_14_LFInst_3_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_15_LFInst_0_U4  ( .A(
        \Red_K2Inst_LFInst_15_LFInst_0_n2 ), .B(Key[62]), .ZN(Red_K2[60]) );
  XNOR2_X1 \Red_K2Inst_LFInst_15_LFInst_0_U3  ( .A(Key[63]), .B(Key[61]), .ZN(
        \Red_K2Inst_LFInst_15_LFInst_0_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_15_LFInst_1_U4  ( .A(
        \Red_K2Inst_LFInst_15_LFInst_1_n2 ), .B(Key[62]), .ZN(Red_K2[61]) );
  XNOR2_X1 \Red_K2Inst_LFInst_15_LFInst_1_U3  ( .A(Key[63]), .B(Key[60]), .ZN(
        \Red_K2Inst_LFInst_15_LFInst_1_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_15_LFInst_2_U4  ( .A(
        \Red_K2Inst_LFInst_15_LFInst_2_n2 ), .B(Key[61]), .ZN(Red_K2[62]) );
  XNOR2_X1 \Red_K2Inst_LFInst_15_LFInst_2_U3  ( .A(Key[63]), .B(Key[60]), .ZN(
        \Red_K2Inst_LFInst_15_LFInst_2_n2 ) );
  XNOR2_X1 \Red_K2Inst_LFInst_15_LFInst_3_U4  ( .A(
        \Red_K2Inst_LFInst_15_LFInst_3_n2 ), .B(Key[61]), .ZN(Red_K2[63]) );
  XNOR2_X1 \Red_K2Inst_LFInst_15_LFInst_3_U3  ( .A(Key[62]), .B(Key[60]), .ZN(
        \Red_K2Inst_LFInst_15_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_0_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_0_LFInst_0_n2 ), .B(AddRoundKeyOutput3[2]), 
        .ZN(Red_SignaltoCheck[0]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_0_LFInst_0_U3  ( .A(AddRoundKeyOutput3[3]), 
        .B(AddRoundKeyOutput3[1]), .ZN(\Red_ToCheckInst_LFInst_0_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_0_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_0_LFInst_1_n2 ), .B(AddRoundKeyOutput3[2]), 
        .ZN(Red_SignaltoCheck[1]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_0_LFInst_1_U3  ( .A(AddRoundKeyOutput3[3]), 
        .B(AddRoundKeyOutput3[0]), .ZN(\Red_ToCheckInst_LFInst_0_LFInst_1_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_0_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_0_LFInst_2_n2 ), .B(AddRoundKeyOutput3[1]), 
        .ZN(Red_SignaltoCheck[2]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_0_LFInst_2_U3  ( .A(AddRoundKeyOutput3[3]), 
        .B(AddRoundKeyOutput3[0]), .ZN(\Red_ToCheckInst_LFInst_0_LFInst_2_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_0_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_0_LFInst_3_n2 ), .B(AddRoundKeyOutput3[1]), 
        .ZN(Red_SignaltoCheck[3]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_0_LFInst_3_U3  ( .A(AddRoundKeyOutput3[2]), 
        .B(AddRoundKeyOutput3[0]), .ZN(\Red_ToCheckInst_LFInst_0_LFInst_3_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_1_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_1_LFInst_0_n2 ), .B(AddRoundKeyOutput3[6]), 
        .ZN(Red_SignaltoCheck[4]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_1_LFInst_0_U3  ( .A(AddRoundKeyOutput3[7]), 
        .B(AddRoundKeyOutput3[5]), .ZN(\Red_ToCheckInst_LFInst_1_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_1_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_1_LFInst_1_n2 ), .B(AddRoundKeyOutput3[6]), 
        .ZN(Red_SignaltoCheck[5]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_1_LFInst_1_U3  ( .A(AddRoundKeyOutput3[7]), 
        .B(AddRoundKeyOutput3[4]), .ZN(\Red_ToCheckInst_LFInst_1_LFInst_1_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_1_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_1_LFInst_2_n2 ), .B(AddRoundKeyOutput3[5]), 
        .ZN(Red_SignaltoCheck[6]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_1_LFInst_2_U3  ( .A(AddRoundKeyOutput3[7]), 
        .B(AddRoundKeyOutput3[4]), .ZN(\Red_ToCheckInst_LFInst_1_LFInst_2_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_1_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_1_LFInst_3_n2 ), .B(AddRoundKeyOutput3[5]), 
        .ZN(Red_SignaltoCheck[7]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_1_LFInst_3_U3  ( .A(AddRoundKeyOutput3[6]), 
        .B(AddRoundKeyOutput3[4]), .ZN(\Red_ToCheckInst_LFInst_1_LFInst_3_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_2_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_2_LFInst_0_n2 ), .B(AddRoundKeyOutput3[10]), 
        .ZN(Red_SignaltoCheck[8]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_2_LFInst_0_U3  ( .A(AddRoundKeyOutput3[11]), 
        .B(AddRoundKeyOutput3[9]), .ZN(\Red_ToCheckInst_LFInst_2_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_2_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_2_LFInst_1_n2 ), .B(AddRoundKeyOutput3[10]), 
        .ZN(Red_SignaltoCheck[9]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_2_LFInst_1_U3  ( .A(AddRoundKeyOutput3[11]), 
        .B(AddRoundKeyOutput3[8]), .ZN(\Red_ToCheckInst_LFInst_2_LFInst_1_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_2_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_2_LFInst_2_n2 ), .B(AddRoundKeyOutput3[9]), 
        .ZN(Red_SignaltoCheck[10]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_2_LFInst_2_U3  ( .A(AddRoundKeyOutput3[11]), 
        .B(AddRoundKeyOutput3[8]), .ZN(\Red_ToCheckInst_LFInst_2_LFInst_2_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_2_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_2_LFInst_3_n2 ), .B(AddRoundKeyOutput3[9]), 
        .ZN(Red_SignaltoCheck[11]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_2_LFInst_3_U3  ( .A(AddRoundKeyOutput3[10]), 
        .B(AddRoundKeyOutput3[8]), .ZN(\Red_ToCheckInst_LFInst_2_LFInst_3_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_3_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_3_LFInst_0_n2 ), .B(AddRoundKeyOutput3[14]), 
        .ZN(Red_SignaltoCheck[12]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_3_LFInst_0_U3  ( .A(AddRoundKeyOutput3[15]), 
        .B(AddRoundKeyOutput3[13]), .ZN(\Red_ToCheckInst_LFInst_3_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_3_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_3_LFInst_1_n2 ), .B(AddRoundKeyOutput3[14]), 
        .ZN(Red_SignaltoCheck[13]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_3_LFInst_1_U3  ( .A(AddRoundKeyOutput3[15]), 
        .B(AddRoundKeyOutput3[12]), .ZN(\Red_ToCheckInst_LFInst_3_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_3_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_3_LFInst_2_n2 ), .B(AddRoundKeyOutput3[13]), 
        .ZN(Red_SignaltoCheck[14]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_3_LFInst_2_U3  ( .A(AddRoundKeyOutput3[15]), 
        .B(AddRoundKeyOutput3[12]), .ZN(\Red_ToCheckInst_LFInst_3_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_3_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_3_LFInst_3_n2 ), .B(AddRoundKeyOutput3[13]), 
        .ZN(Red_SignaltoCheck[15]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_3_LFInst_3_U3  ( .A(AddRoundKeyOutput3[14]), 
        .B(AddRoundKeyOutput3[12]), .ZN(\Red_ToCheckInst_LFInst_3_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_4_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_4_LFInst_0_n2 ), .B(AddRoundKeyOutput3[18]), 
        .ZN(Red_SignaltoCheck[16]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_4_LFInst_0_U3  ( .A(AddRoundKeyOutput3[19]), 
        .B(AddRoundKeyOutput3[17]), .ZN(\Red_ToCheckInst_LFInst_4_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_4_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_4_LFInst_1_n2 ), .B(AddRoundKeyOutput3[18]), 
        .ZN(Red_SignaltoCheck[17]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_4_LFInst_1_U3  ( .A(AddRoundKeyOutput3[19]), 
        .B(AddRoundKeyOutput3[16]), .ZN(\Red_ToCheckInst_LFInst_4_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_4_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_4_LFInst_2_n2 ), .B(AddRoundKeyOutput3[17]), 
        .ZN(Red_SignaltoCheck[18]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_4_LFInst_2_U3  ( .A(AddRoundKeyOutput3[19]), 
        .B(AddRoundKeyOutput3[16]), .ZN(\Red_ToCheckInst_LFInst_4_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_4_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_4_LFInst_3_n2 ), .B(AddRoundKeyOutput3[17]), 
        .ZN(Red_SignaltoCheck[19]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_4_LFInst_3_U3  ( .A(AddRoundKeyOutput3[18]), 
        .B(AddRoundKeyOutput3[16]), .ZN(\Red_ToCheckInst_LFInst_4_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_5_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_5_LFInst_0_n2 ), .B(AddRoundKeyOutput3[22]), 
        .ZN(Red_SignaltoCheck[20]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_5_LFInst_0_U3  ( .A(AddRoundKeyOutput3[23]), 
        .B(AddRoundKeyOutput3[21]), .ZN(\Red_ToCheckInst_LFInst_5_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_5_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_5_LFInst_1_n2 ), .B(AddRoundKeyOutput3[22]), 
        .ZN(Red_SignaltoCheck[21]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_5_LFInst_1_U3  ( .A(AddRoundKeyOutput3[23]), 
        .B(AddRoundKeyOutput3[20]), .ZN(\Red_ToCheckInst_LFInst_5_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_5_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_5_LFInst_2_n2 ), .B(AddRoundKeyOutput3[21]), 
        .ZN(Red_SignaltoCheck[22]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_5_LFInst_2_U3  ( .A(AddRoundKeyOutput3[23]), 
        .B(AddRoundKeyOutput3[20]), .ZN(\Red_ToCheckInst_LFInst_5_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_5_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_5_LFInst_3_n2 ), .B(AddRoundKeyOutput3[21]), 
        .ZN(Red_SignaltoCheck[23]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_5_LFInst_3_U3  ( .A(AddRoundKeyOutput3[22]), 
        .B(AddRoundKeyOutput3[20]), .ZN(\Red_ToCheckInst_LFInst_5_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_6_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_6_LFInst_0_n2 ), .B(AddRoundKeyOutput3[26]), 
        .ZN(Red_SignaltoCheck[24]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_6_LFInst_0_U3  ( .A(AddRoundKeyOutput3[27]), 
        .B(AddRoundKeyOutput3[25]), .ZN(\Red_ToCheckInst_LFInst_6_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_6_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_6_LFInst_1_n2 ), .B(AddRoundKeyOutput3[26]), 
        .ZN(Red_SignaltoCheck[25]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_6_LFInst_1_U3  ( .A(AddRoundKeyOutput3[27]), 
        .B(AddRoundKeyOutput3[24]), .ZN(\Red_ToCheckInst_LFInst_6_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_6_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_6_LFInst_2_n2 ), .B(AddRoundKeyOutput3[25]), 
        .ZN(Red_SignaltoCheck[26]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_6_LFInst_2_U3  ( .A(AddRoundKeyOutput3[27]), 
        .B(AddRoundKeyOutput3[24]), .ZN(\Red_ToCheckInst_LFInst_6_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_6_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_6_LFInst_3_n2 ), .B(AddRoundKeyOutput3[25]), 
        .ZN(Red_SignaltoCheck[27]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_6_LFInst_3_U3  ( .A(AddRoundKeyOutput3[26]), 
        .B(AddRoundKeyOutput3[24]), .ZN(\Red_ToCheckInst_LFInst_6_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_7_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_7_LFInst_0_n2 ), .B(AddRoundKeyOutput3[30]), 
        .ZN(Red_SignaltoCheck[28]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_7_LFInst_0_U3  ( .A(AddRoundKeyOutput3[31]), 
        .B(AddRoundKeyOutput3[29]), .ZN(\Red_ToCheckInst_LFInst_7_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_7_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_7_LFInst_1_n2 ), .B(AddRoundKeyOutput3[30]), 
        .ZN(Red_SignaltoCheck[29]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_7_LFInst_1_U3  ( .A(AddRoundKeyOutput3[31]), 
        .B(AddRoundKeyOutput3[28]), .ZN(\Red_ToCheckInst_LFInst_7_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_7_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_7_LFInst_2_n2 ), .B(AddRoundKeyOutput3[29]), 
        .ZN(Red_SignaltoCheck[30]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_7_LFInst_2_U3  ( .A(AddRoundKeyOutput3[31]), 
        .B(AddRoundKeyOutput3[28]), .ZN(\Red_ToCheckInst_LFInst_7_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_7_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_7_LFInst_3_n2 ), .B(AddRoundKeyOutput3[29]), 
        .ZN(Red_SignaltoCheck[31]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_7_LFInst_3_U3  ( .A(AddRoundKeyOutput3[30]), 
        .B(AddRoundKeyOutput3[28]), .ZN(\Red_ToCheckInst_LFInst_7_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_8_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_8_LFInst_0_n2 ), .B(AddRoundKeyOutput3[34]), 
        .ZN(Red_SignaltoCheck[32]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_8_LFInst_0_U3  ( .A(AddRoundKeyOutput3[35]), 
        .B(AddRoundKeyOutput3[33]), .ZN(\Red_ToCheckInst_LFInst_8_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_8_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_8_LFInst_1_n2 ), .B(AddRoundKeyOutput3[34]), 
        .ZN(Red_SignaltoCheck[33]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_8_LFInst_1_U3  ( .A(AddRoundKeyOutput3[35]), 
        .B(AddRoundKeyOutput3[32]), .ZN(\Red_ToCheckInst_LFInst_8_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_8_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_8_LFInst_2_n2 ), .B(AddRoundKeyOutput3[33]), 
        .ZN(Red_SignaltoCheck[34]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_8_LFInst_2_U3  ( .A(AddRoundKeyOutput3[35]), 
        .B(AddRoundKeyOutput3[32]), .ZN(\Red_ToCheckInst_LFInst_8_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_8_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_8_LFInst_3_n2 ), .B(AddRoundKeyOutput3[33]), 
        .ZN(Red_SignaltoCheck[35]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_8_LFInst_3_U3  ( .A(AddRoundKeyOutput3[34]), 
        .B(AddRoundKeyOutput3[32]), .ZN(\Red_ToCheckInst_LFInst_8_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_9_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_9_LFInst_0_n2 ), .B(AddRoundKeyOutput3[38]), 
        .ZN(Red_SignaltoCheck[36]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_9_LFInst_0_U3  ( .A(AddRoundKeyOutput3[39]), 
        .B(AddRoundKeyOutput3[37]), .ZN(\Red_ToCheckInst_LFInst_9_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_9_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_9_LFInst_1_n2 ), .B(AddRoundKeyOutput3[38]), 
        .ZN(Red_SignaltoCheck[37]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_9_LFInst_1_U3  ( .A(AddRoundKeyOutput3[39]), 
        .B(AddRoundKeyOutput3[36]), .ZN(\Red_ToCheckInst_LFInst_9_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_9_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_9_LFInst_2_n2 ), .B(AddRoundKeyOutput3[37]), 
        .ZN(Red_SignaltoCheck[38]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_9_LFInst_2_U3  ( .A(AddRoundKeyOutput3[39]), 
        .B(AddRoundKeyOutput3[36]), .ZN(\Red_ToCheckInst_LFInst_9_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_9_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_9_LFInst_3_n2 ), .B(AddRoundKeyOutput3[37]), 
        .ZN(Red_SignaltoCheck[39]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_9_LFInst_3_U3  ( .A(AddRoundKeyOutput3[38]), 
        .B(AddRoundKeyOutput3[36]), .ZN(\Red_ToCheckInst_LFInst_9_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_10_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_10_LFInst_0_n2 ), .B(AddRoundKeyOutput3[42]), 
        .ZN(Red_SignaltoCheck[40]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_10_LFInst_0_U3  ( .A(AddRoundKeyOutput3[43]), .B(AddRoundKeyOutput3[41]), .ZN(\Red_ToCheckInst_LFInst_10_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_10_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_10_LFInst_1_n2 ), .B(AddRoundKeyOutput3[42]), 
        .ZN(Red_SignaltoCheck[41]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_10_LFInst_1_U3  ( .A(AddRoundKeyOutput3[43]), .B(AddRoundKeyOutput3[40]), .ZN(\Red_ToCheckInst_LFInst_10_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_10_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_10_LFInst_2_n2 ), .B(AddRoundKeyOutput3[41]), 
        .ZN(Red_SignaltoCheck[42]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_10_LFInst_2_U3  ( .A(AddRoundKeyOutput3[43]), .B(AddRoundKeyOutput3[40]), .ZN(\Red_ToCheckInst_LFInst_10_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_10_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_10_LFInst_3_n2 ), .B(AddRoundKeyOutput3[41]), 
        .ZN(Red_SignaltoCheck[43]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_10_LFInst_3_U3  ( .A(AddRoundKeyOutput3[42]), .B(AddRoundKeyOutput3[40]), .ZN(\Red_ToCheckInst_LFInst_10_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_11_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_11_LFInst_0_n2 ), .B(AddRoundKeyOutput3[46]), 
        .ZN(Red_SignaltoCheck[44]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_11_LFInst_0_U3  ( .A(AddRoundKeyOutput3[47]), .B(AddRoundKeyOutput3[45]), .ZN(\Red_ToCheckInst_LFInst_11_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_11_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_11_LFInst_1_n2 ), .B(AddRoundKeyOutput3[46]), 
        .ZN(Red_SignaltoCheck[45]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_11_LFInst_1_U3  ( .A(AddRoundKeyOutput3[47]), .B(AddRoundKeyOutput3[44]), .ZN(\Red_ToCheckInst_LFInst_11_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_11_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_11_LFInst_2_n2 ), .B(AddRoundKeyOutput3[45]), 
        .ZN(Red_SignaltoCheck[46]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_11_LFInst_2_U3  ( .A(AddRoundKeyOutput3[47]), .B(AddRoundKeyOutput3[44]), .ZN(\Red_ToCheckInst_LFInst_11_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_11_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_11_LFInst_3_n2 ), .B(AddRoundKeyOutput3[45]), 
        .ZN(Red_SignaltoCheck[47]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_11_LFInst_3_U3  ( .A(AddRoundKeyOutput3[46]), .B(AddRoundKeyOutput3[44]), .ZN(\Red_ToCheckInst_LFInst_11_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_12_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_12_LFInst_0_n2 ), .B(AddRoundKeyOutput3[50]), 
        .ZN(Red_SignaltoCheck[48]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_12_LFInst_0_U3  ( .A(AddRoundKeyOutput3[51]), .B(AddRoundKeyOutput3[49]), .ZN(\Red_ToCheckInst_LFInst_12_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_12_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_12_LFInst_1_n2 ), .B(AddRoundKeyOutput3[50]), 
        .ZN(Red_SignaltoCheck[49]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_12_LFInst_1_U3  ( .A(AddRoundKeyOutput3[51]), .B(AddRoundKeyOutput3[48]), .ZN(\Red_ToCheckInst_LFInst_12_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_12_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_12_LFInst_2_n2 ), .B(AddRoundKeyOutput3[49]), 
        .ZN(Red_SignaltoCheck[50]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_12_LFInst_2_U3  ( .A(AddRoundKeyOutput3[51]), .B(AddRoundKeyOutput3[48]), .ZN(\Red_ToCheckInst_LFInst_12_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_12_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_12_LFInst_3_n2 ), .B(AddRoundKeyOutput3[49]), 
        .ZN(Red_SignaltoCheck[51]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_12_LFInst_3_U3  ( .A(AddRoundKeyOutput3[50]), .B(AddRoundKeyOutput3[48]), .ZN(\Red_ToCheckInst_LFInst_12_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_13_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_13_LFInst_0_n2 ), .B(AddRoundKeyOutput3[54]), 
        .ZN(Red_SignaltoCheck[52]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_13_LFInst_0_U3  ( .A(AddRoundKeyOutput3[55]), .B(AddRoundKeyOutput3[53]), .ZN(\Red_ToCheckInst_LFInst_13_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_13_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_13_LFInst_1_n2 ), .B(AddRoundKeyOutput3[54]), 
        .ZN(Red_SignaltoCheck[53]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_13_LFInst_1_U3  ( .A(AddRoundKeyOutput3[55]), .B(AddRoundKeyOutput3[52]), .ZN(\Red_ToCheckInst_LFInst_13_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_13_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_13_LFInst_2_n2 ), .B(AddRoundKeyOutput3[53]), 
        .ZN(Red_SignaltoCheck[54]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_13_LFInst_2_U3  ( .A(AddRoundKeyOutput3[55]), .B(AddRoundKeyOutput3[52]), .ZN(\Red_ToCheckInst_LFInst_13_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_13_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_13_LFInst_3_n2 ), .B(AddRoundKeyOutput3[53]), 
        .ZN(Red_SignaltoCheck[55]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_13_LFInst_3_U3  ( .A(AddRoundKeyOutput3[54]), .B(AddRoundKeyOutput3[52]), .ZN(\Red_ToCheckInst_LFInst_13_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_14_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_14_LFInst_0_n2 ), .B(AddRoundKeyOutput3[58]), 
        .ZN(Red_SignaltoCheck[56]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_14_LFInst_0_U3  ( .A(AddRoundKeyOutput3[59]), .B(AddRoundKeyOutput3[57]), .ZN(\Red_ToCheckInst_LFInst_14_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_14_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_14_LFInst_1_n2 ), .B(AddRoundKeyOutput3[58]), 
        .ZN(Red_SignaltoCheck[57]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_14_LFInst_1_U3  ( .A(AddRoundKeyOutput3[59]), .B(AddRoundKeyOutput3[56]), .ZN(\Red_ToCheckInst_LFInst_14_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_14_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_14_LFInst_2_n2 ), .B(AddRoundKeyOutput3[57]), 
        .ZN(Red_SignaltoCheck[58]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_14_LFInst_2_U3  ( .A(AddRoundKeyOutput3[59]), .B(AddRoundKeyOutput3[56]), .ZN(\Red_ToCheckInst_LFInst_14_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_14_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_14_LFInst_3_n2 ), .B(AddRoundKeyOutput3[57]), 
        .ZN(Red_SignaltoCheck[59]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_14_LFInst_3_U3  ( .A(AddRoundKeyOutput3[58]), .B(AddRoundKeyOutput3[56]), .ZN(\Red_ToCheckInst_LFInst_14_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_15_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_15_LFInst_0_n2 ), .B(AddRoundKeyOutput3[62]), 
        .ZN(Red_SignaltoCheck[60]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_15_LFInst_0_U3  ( .A(AddRoundKeyOutput3[63]), .B(AddRoundKeyOutput3[61]), .ZN(\Red_ToCheckInst_LFInst_15_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_15_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_15_LFInst_1_n2 ), .B(AddRoundKeyOutput3[62]), 
        .ZN(Red_SignaltoCheck[61]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_15_LFInst_1_U3  ( .A(AddRoundKeyOutput3[63]), .B(AddRoundKeyOutput3[60]), .ZN(\Red_ToCheckInst_LFInst_15_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_15_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_15_LFInst_2_n2 ), .B(AddRoundKeyOutput3[61]), 
        .ZN(Red_SignaltoCheck[62]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_15_LFInst_2_U3  ( .A(AddRoundKeyOutput3[63]), .B(AddRoundKeyOutput3[60]), .ZN(\Red_ToCheckInst_LFInst_15_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_15_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_15_LFInst_3_n2 ), .B(AddRoundKeyOutput3[61]), 
        .ZN(Red_SignaltoCheck[63]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_15_LFInst_3_U3  ( .A(AddRoundKeyOutput3[62]), .B(AddRoundKeyOutput3[60]), .ZN(\Red_ToCheckInst_LFInst_15_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_16_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_16_LFInst_0_n2 ), .B(AddRoundKeyOutput2[2]), 
        .ZN(Red_SignaltoCheck[64]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_16_LFInst_0_U3  ( .A(AddRoundKeyOutput2[3]), 
        .B(AddRoundKeyOutput2[1]), .ZN(\Red_ToCheckInst_LFInst_16_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_16_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_16_LFInst_1_n2 ), .B(AddRoundKeyOutput2[2]), 
        .ZN(Red_SignaltoCheck[65]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_16_LFInst_1_U3  ( .A(AddRoundKeyOutput2[3]), 
        .B(AddRoundKeyOutput2[0]), .ZN(\Red_ToCheckInst_LFInst_16_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_16_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_16_LFInst_2_n2 ), .B(AddRoundKeyOutput2[1]), 
        .ZN(Red_SignaltoCheck[66]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_16_LFInst_2_U3  ( .A(AddRoundKeyOutput2[3]), 
        .B(AddRoundKeyOutput2[0]), .ZN(\Red_ToCheckInst_LFInst_16_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_16_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_16_LFInst_3_n2 ), .B(AddRoundKeyOutput2[1]), 
        .ZN(Red_SignaltoCheck[67]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_16_LFInst_3_U3  ( .A(AddRoundKeyOutput2[2]), 
        .B(AddRoundKeyOutput2[0]), .ZN(\Red_ToCheckInst_LFInst_16_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_17_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_17_LFInst_0_n2 ), .B(AddRoundKeyOutput2[6]), 
        .ZN(Red_SignaltoCheck[68]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_17_LFInst_0_U3  ( .A(AddRoundKeyOutput2[7]), 
        .B(AddRoundKeyOutput2[5]), .ZN(\Red_ToCheckInst_LFInst_17_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_17_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_17_LFInst_1_n2 ), .B(AddRoundKeyOutput2[6]), 
        .ZN(Red_SignaltoCheck[69]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_17_LFInst_1_U3  ( .A(AddRoundKeyOutput2[7]), 
        .B(AddRoundKeyOutput2[4]), .ZN(\Red_ToCheckInst_LFInst_17_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_17_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_17_LFInst_2_n2 ), .B(AddRoundKeyOutput2[5]), 
        .ZN(Red_SignaltoCheck[70]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_17_LFInst_2_U3  ( .A(AddRoundKeyOutput2[7]), 
        .B(AddRoundKeyOutput2[4]), .ZN(\Red_ToCheckInst_LFInst_17_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_17_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_17_LFInst_3_n2 ), .B(AddRoundKeyOutput2[5]), 
        .ZN(Red_SignaltoCheck[71]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_17_LFInst_3_U3  ( .A(AddRoundKeyOutput2[6]), 
        .B(AddRoundKeyOutput2[4]), .ZN(\Red_ToCheckInst_LFInst_17_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_18_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_18_LFInst_0_n2 ), .B(AddRoundKeyOutput2[10]), 
        .ZN(Red_SignaltoCheck[72]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_18_LFInst_0_U3  ( .A(AddRoundKeyOutput2[11]), .B(AddRoundKeyOutput2[9]), .ZN(\Red_ToCheckInst_LFInst_18_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_18_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_18_LFInst_1_n2 ), .B(AddRoundKeyOutput2[10]), 
        .ZN(Red_SignaltoCheck[73]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_18_LFInst_1_U3  ( .A(AddRoundKeyOutput2[11]), .B(AddRoundKeyOutput2[8]), .ZN(\Red_ToCheckInst_LFInst_18_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_18_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_18_LFInst_2_n2 ), .B(AddRoundKeyOutput2[9]), 
        .ZN(Red_SignaltoCheck[74]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_18_LFInst_2_U3  ( .A(AddRoundKeyOutput2[11]), .B(AddRoundKeyOutput2[8]), .ZN(\Red_ToCheckInst_LFInst_18_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_18_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_18_LFInst_3_n2 ), .B(AddRoundKeyOutput2[9]), 
        .ZN(Red_SignaltoCheck[75]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_18_LFInst_3_U3  ( .A(AddRoundKeyOutput2[10]), .B(AddRoundKeyOutput2[8]), .ZN(\Red_ToCheckInst_LFInst_18_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_19_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_19_LFInst_0_n2 ), .B(AddRoundKeyOutput2[14]), 
        .ZN(Red_SignaltoCheck[76]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_19_LFInst_0_U3  ( .A(AddRoundKeyOutput2[15]), .B(AddRoundKeyOutput2[13]), .ZN(\Red_ToCheckInst_LFInst_19_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_19_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_19_LFInst_1_n2 ), .B(AddRoundKeyOutput2[14]), 
        .ZN(Red_SignaltoCheck[77]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_19_LFInst_1_U3  ( .A(AddRoundKeyOutput2[15]), .B(AddRoundKeyOutput2[12]), .ZN(\Red_ToCheckInst_LFInst_19_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_19_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_19_LFInst_2_n2 ), .B(AddRoundKeyOutput2[13]), 
        .ZN(Red_SignaltoCheck[78]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_19_LFInst_2_U3  ( .A(AddRoundKeyOutput2[15]), .B(AddRoundKeyOutput2[12]), .ZN(\Red_ToCheckInst_LFInst_19_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_19_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_19_LFInst_3_n2 ), .B(AddRoundKeyOutput2[13]), 
        .ZN(Red_SignaltoCheck[79]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_19_LFInst_3_U3  ( .A(AddRoundKeyOutput2[14]), .B(AddRoundKeyOutput2[12]), .ZN(\Red_ToCheckInst_LFInst_19_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_20_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_20_LFInst_0_n2 ), .B(AddRoundKeyOutput2[18]), 
        .ZN(Red_SignaltoCheck[80]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_20_LFInst_0_U3  ( .A(AddRoundKeyOutput2[19]), .B(AddRoundKeyOutput2[17]), .ZN(\Red_ToCheckInst_LFInst_20_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_20_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_20_LFInst_1_n2 ), .B(AddRoundKeyOutput2[18]), 
        .ZN(Red_SignaltoCheck[81]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_20_LFInst_1_U3  ( .A(AddRoundKeyOutput2[19]), .B(AddRoundKeyOutput2[16]), .ZN(\Red_ToCheckInst_LFInst_20_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_20_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_20_LFInst_2_n2 ), .B(AddRoundKeyOutput2[17]), 
        .ZN(Red_SignaltoCheck[82]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_20_LFInst_2_U3  ( .A(AddRoundKeyOutput2[19]), .B(AddRoundKeyOutput2[16]), .ZN(\Red_ToCheckInst_LFInst_20_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_20_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_20_LFInst_3_n2 ), .B(AddRoundKeyOutput2[17]), 
        .ZN(Red_SignaltoCheck[83]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_20_LFInst_3_U3  ( .A(AddRoundKeyOutput2[18]), .B(AddRoundKeyOutput2[16]), .ZN(\Red_ToCheckInst_LFInst_20_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_21_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_21_LFInst_0_n2 ), .B(AddRoundKeyOutput2[22]), 
        .ZN(Red_SignaltoCheck[84]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_21_LFInst_0_U3  ( .A(AddRoundKeyOutput2[23]), .B(AddRoundKeyOutput2[21]), .ZN(\Red_ToCheckInst_LFInst_21_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_21_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_21_LFInst_1_n2 ), .B(AddRoundKeyOutput2[22]), 
        .ZN(Red_SignaltoCheck[85]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_21_LFInst_1_U3  ( .A(AddRoundKeyOutput2[23]), .B(AddRoundKeyOutput2[20]), .ZN(\Red_ToCheckInst_LFInst_21_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_21_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_21_LFInst_2_n2 ), .B(AddRoundKeyOutput2[21]), 
        .ZN(Red_SignaltoCheck[86]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_21_LFInst_2_U3  ( .A(AddRoundKeyOutput2[23]), .B(AddRoundKeyOutput2[20]), .ZN(\Red_ToCheckInst_LFInst_21_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_21_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_21_LFInst_3_n2 ), .B(AddRoundKeyOutput2[21]), 
        .ZN(Red_SignaltoCheck[87]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_21_LFInst_3_U3  ( .A(AddRoundKeyOutput2[22]), .B(AddRoundKeyOutput2[20]), .ZN(\Red_ToCheckInst_LFInst_21_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_22_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_22_LFInst_0_n2 ), .B(AddRoundKeyOutput2[26]), 
        .ZN(Red_SignaltoCheck[88]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_22_LFInst_0_U3  ( .A(AddRoundKeyOutput2[27]), .B(AddRoundKeyOutput2[25]), .ZN(\Red_ToCheckInst_LFInst_22_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_22_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_22_LFInst_1_n2 ), .B(AddRoundKeyOutput2[26]), 
        .ZN(Red_SignaltoCheck[89]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_22_LFInst_1_U3  ( .A(AddRoundKeyOutput2[27]), .B(AddRoundKeyOutput2[24]), .ZN(\Red_ToCheckInst_LFInst_22_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_22_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_22_LFInst_2_n2 ), .B(AddRoundKeyOutput2[25]), 
        .ZN(Red_SignaltoCheck[90]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_22_LFInst_2_U3  ( .A(AddRoundKeyOutput2[27]), .B(AddRoundKeyOutput2[24]), .ZN(\Red_ToCheckInst_LFInst_22_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_22_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_22_LFInst_3_n2 ), .B(AddRoundKeyOutput2[25]), 
        .ZN(Red_SignaltoCheck[91]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_22_LFInst_3_U3  ( .A(AddRoundKeyOutput2[26]), .B(AddRoundKeyOutput2[24]), .ZN(\Red_ToCheckInst_LFInst_22_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_23_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_23_LFInst_0_n2 ), .B(AddRoundKeyOutput2[30]), 
        .ZN(Red_SignaltoCheck[92]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_23_LFInst_0_U3  ( .A(AddRoundKeyOutput2[31]), .B(AddRoundKeyOutput2[29]), .ZN(\Red_ToCheckInst_LFInst_23_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_23_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_23_LFInst_1_n2 ), .B(AddRoundKeyOutput2[30]), 
        .ZN(Red_SignaltoCheck[93]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_23_LFInst_1_U3  ( .A(AddRoundKeyOutput2[31]), .B(AddRoundKeyOutput2[28]), .ZN(\Red_ToCheckInst_LFInst_23_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_23_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_23_LFInst_2_n2 ), .B(AddRoundKeyOutput2[29]), 
        .ZN(Red_SignaltoCheck[94]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_23_LFInst_2_U3  ( .A(AddRoundKeyOutput2[31]), .B(AddRoundKeyOutput2[28]), .ZN(\Red_ToCheckInst_LFInst_23_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_23_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_23_LFInst_3_n2 ), .B(AddRoundKeyOutput2[29]), 
        .ZN(Red_SignaltoCheck[95]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_23_LFInst_3_U3  ( .A(AddRoundKeyOutput2[30]), .B(AddRoundKeyOutput2[28]), .ZN(\Red_ToCheckInst_LFInst_23_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_24_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_24_LFInst_0_n2 ), .B(AddRoundKeyOutput2[34]), 
        .ZN(Red_SignaltoCheck[96]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_24_LFInst_0_U3  ( .A(AddRoundKeyOutput2[35]), .B(AddRoundKeyOutput2[33]), .ZN(\Red_ToCheckInst_LFInst_24_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_24_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_24_LFInst_1_n2 ), .B(AddRoundKeyOutput2[34]), 
        .ZN(Red_SignaltoCheck[97]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_24_LFInst_1_U3  ( .A(AddRoundKeyOutput2[35]), .B(AddRoundKeyOutput2[32]), .ZN(\Red_ToCheckInst_LFInst_24_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_24_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_24_LFInst_2_n2 ), .B(AddRoundKeyOutput2[33]), 
        .ZN(Red_SignaltoCheck[98]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_24_LFInst_2_U3  ( .A(AddRoundKeyOutput2[35]), .B(AddRoundKeyOutput2[32]), .ZN(\Red_ToCheckInst_LFInst_24_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_24_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_24_LFInst_3_n2 ), .B(AddRoundKeyOutput2[33]), 
        .ZN(Red_SignaltoCheck[99]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_24_LFInst_3_U3  ( .A(AddRoundKeyOutput2[34]), .B(AddRoundKeyOutput2[32]), .ZN(\Red_ToCheckInst_LFInst_24_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_25_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_25_LFInst_0_n2 ), .B(AddRoundKeyOutput2[38]), 
        .ZN(Red_SignaltoCheck[100]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_25_LFInst_0_U3  ( .A(AddRoundKeyOutput2[39]), .B(AddRoundKeyOutput2[37]), .ZN(\Red_ToCheckInst_LFInst_25_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_25_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_25_LFInst_1_n2 ), .B(AddRoundKeyOutput2[38]), 
        .ZN(Red_SignaltoCheck[101]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_25_LFInst_1_U3  ( .A(AddRoundKeyOutput2[39]), .B(AddRoundKeyOutput2[36]), .ZN(\Red_ToCheckInst_LFInst_25_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_25_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_25_LFInst_2_n2 ), .B(AddRoundKeyOutput2[37]), 
        .ZN(Red_SignaltoCheck[102]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_25_LFInst_2_U3  ( .A(AddRoundKeyOutput2[39]), .B(AddRoundKeyOutput2[36]), .ZN(\Red_ToCheckInst_LFInst_25_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_25_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_25_LFInst_3_n2 ), .B(AddRoundKeyOutput2[37]), 
        .ZN(Red_SignaltoCheck[103]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_25_LFInst_3_U3  ( .A(AddRoundKeyOutput2[38]), .B(AddRoundKeyOutput2[36]), .ZN(\Red_ToCheckInst_LFInst_25_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_26_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_26_LFInst_0_n2 ), .B(AddRoundKeyOutput2[42]), 
        .ZN(Red_SignaltoCheck[104]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_26_LFInst_0_U3  ( .A(AddRoundKeyOutput2[43]), .B(AddRoundKeyOutput2[41]), .ZN(\Red_ToCheckInst_LFInst_26_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_26_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_26_LFInst_1_n2 ), .B(AddRoundKeyOutput2[42]), 
        .ZN(Red_SignaltoCheck[105]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_26_LFInst_1_U3  ( .A(AddRoundKeyOutput2[43]), .B(AddRoundKeyOutput2[40]), .ZN(\Red_ToCheckInst_LFInst_26_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_26_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_26_LFInst_2_n2 ), .B(AddRoundKeyOutput2[41]), 
        .ZN(Red_SignaltoCheck[106]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_26_LFInst_2_U3  ( .A(AddRoundKeyOutput2[43]), .B(AddRoundKeyOutput2[40]), .ZN(\Red_ToCheckInst_LFInst_26_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_26_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_26_LFInst_3_n2 ), .B(AddRoundKeyOutput2[41]), 
        .ZN(Red_SignaltoCheck[107]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_26_LFInst_3_U3  ( .A(AddRoundKeyOutput2[42]), .B(AddRoundKeyOutput2[40]), .ZN(\Red_ToCheckInst_LFInst_26_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_27_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_27_LFInst_0_n2 ), .B(AddRoundKeyOutput2[46]), 
        .ZN(Red_SignaltoCheck[108]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_27_LFInst_0_U3  ( .A(AddRoundKeyOutput2[47]), .B(AddRoundKeyOutput2[45]), .ZN(\Red_ToCheckInst_LFInst_27_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_27_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_27_LFInst_1_n2 ), .B(AddRoundKeyOutput2[46]), 
        .ZN(Red_SignaltoCheck[109]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_27_LFInst_1_U3  ( .A(AddRoundKeyOutput2[47]), .B(AddRoundKeyOutput2[44]), .ZN(\Red_ToCheckInst_LFInst_27_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_27_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_27_LFInst_2_n2 ), .B(AddRoundKeyOutput2[45]), 
        .ZN(Red_SignaltoCheck[110]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_27_LFInst_2_U3  ( .A(AddRoundKeyOutput2[47]), .B(AddRoundKeyOutput2[44]), .ZN(\Red_ToCheckInst_LFInst_27_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_27_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_27_LFInst_3_n2 ), .B(AddRoundKeyOutput2[45]), 
        .ZN(Red_SignaltoCheck[111]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_27_LFInst_3_U3  ( .A(AddRoundKeyOutput2[46]), .B(AddRoundKeyOutput2[44]), .ZN(\Red_ToCheckInst_LFInst_27_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_28_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_28_LFInst_0_n2 ), .B(AddRoundKeyOutput2[50]), 
        .ZN(Red_SignaltoCheck[112]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_28_LFInst_0_U3  ( .A(AddRoundKeyOutput2[51]), .B(AddRoundKeyOutput2[49]), .ZN(\Red_ToCheckInst_LFInst_28_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_28_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_28_LFInst_1_n2 ), .B(AddRoundKeyOutput2[50]), 
        .ZN(Red_SignaltoCheck[113]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_28_LFInst_1_U3  ( .A(AddRoundKeyOutput2[51]), .B(AddRoundKeyOutput2[48]), .ZN(\Red_ToCheckInst_LFInst_28_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_28_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_28_LFInst_2_n2 ), .B(AddRoundKeyOutput2[49]), 
        .ZN(Red_SignaltoCheck[114]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_28_LFInst_2_U3  ( .A(AddRoundKeyOutput2[51]), .B(AddRoundKeyOutput2[48]), .ZN(\Red_ToCheckInst_LFInst_28_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_28_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_28_LFInst_3_n2 ), .B(AddRoundKeyOutput2[49]), 
        .ZN(Red_SignaltoCheck[115]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_28_LFInst_3_U3  ( .A(AddRoundKeyOutput2[50]), .B(AddRoundKeyOutput2[48]), .ZN(\Red_ToCheckInst_LFInst_28_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_29_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_29_LFInst_0_n2 ), .B(AddRoundKeyOutput2[54]), 
        .ZN(Red_SignaltoCheck[116]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_29_LFInst_0_U3  ( .A(AddRoundKeyOutput2[55]), .B(AddRoundKeyOutput2[53]), .ZN(\Red_ToCheckInst_LFInst_29_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_29_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_29_LFInst_1_n2 ), .B(AddRoundKeyOutput2[54]), 
        .ZN(Red_SignaltoCheck[117]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_29_LFInst_1_U3  ( .A(AddRoundKeyOutput2[55]), .B(AddRoundKeyOutput2[52]), .ZN(\Red_ToCheckInst_LFInst_29_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_29_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_29_LFInst_2_n2 ), .B(AddRoundKeyOutput2[53]), 
        .ZN(Red_SignaltoCheck[118]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_29_LFInst_2_U3  ( .A(AddRoundKeyOutput2[55]), .B(AddRoundKeyOutput2[52]), .ZN(\Red_ToCheckInst_LFInst_29_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_29_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_29_LFInst_3_n2 ), .B(AddRoundKeyOutput2[53]), 
        .ZN(Red_SignaltoCheck[119]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_29_LFInst_3_U3  ( .A(AddRoundKeyOutput2[54]), .B(AddRoundKeyOutput2[52]), .ZN(\Red_ToCheckInst_LFInst_29_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_30_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_30_LFInst_0_n2 ), .B(AddRoundKeyOutput2[58]), 
        .ZN(Red_SignaltoCheck[120]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_30_LFInst_0_U3  ( .A(AddRoundKeyOutput2[59]), .B(AddRoundKeyOutput2[57]), .ZN(\Red_ToCheckInst_LFInst_30_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_30_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_30_LFInst_1_n2 ), .B(AddRoundKeyOutput2[58]), 
        .ZN(Red_SignaltoCheck[121]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_30_LFInst_1_U3  ( .A(AddRoundKeyOutput2[59]), .B(AddRoundKeyOutput2[56]), .ZN(\Red_ToCheckInst_LFInst_30_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_30_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_30_LFInst_2_n2 ), .B(AddRoundKeyOutput2[57]), 
        .ZN(Red_SignaltoCheck[122]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_30_LFInst_2_U3  ( .A(AddRoundKeyOutput2[59]), .B(AddRoundKeyOutput2[56]), .ZN(\Red_ToCheckInst_LFInst_30_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_30_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_30_LFInst_3_n2 ), .B(AddRoundKeyOutput2[57]), 
        .ZN(Red_SignaltoCheck[123]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_30_LFInst_3_U3  ( .A(AddRoundKeyOutput2[58]), .B(AddRoundKeyOutput2[56]), .ZN(\Red_ToCheckInst_LFInst_30_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_31_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_31_LFInst_0_n2 ), .B(AddRoundKeyOutput2[62]), 
        .ZN(Red_SignaltoCheck[124]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_31_LFInst_0_U3  ( .A(AddRoundKeyOutput2[63]), .B(AddRoundKeyOutput2[61]), .ZN(\Red_ToCheckInst_LFInst_31_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_31_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_31_LFInst_1_n2 ), .B(AddRoundKeyOutput2[62]), 
        .ZN(Red_SignaltoCheck[125]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_31_LFInst_1_U3  ( .A(AddRoundKeyOutput2[63]), .B(AddRoundKeyOutput2[60]), .ZN(\Red_ToCheckInst_LFInst_31_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_31_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_31_LFInst_2_n2 ), .B(AddRoundKeyOutput2[61]), 
        .ZN(Red_SignaltoCheck[126]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_31_LFInst_2_U3  ( .A(AddRoundKeyOutput2[63]), .B(AddRoundKeyOutput2[60]), .ZN(\Red_ToCheckInst_LFInst_31_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_31_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_31_LFInst_3_n2 ), .B(AddRoundKeyOutput2[61]), 
        .ZN(Red_SignaltoCheck[127]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_31_LFInst_3_U3  ( .A(AddRoundKeyOutput2[62]), .B(AddRoundKeyOutput2[60]), .ZN(\Red_ToCheckInst_LFInst_31_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_32_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_32_LFInst_0_n2 ), .B(AddRoundKeyOutput[2]), 
        .ZN(Red_SignaltoCheck[128]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_32_LFInst_0_U3  ( .A(AddRoundKeyOutput[3]), 
        .B(AddRoundKeyOutput[1]), .ZN(\Red_ToCheckInst_LFInst_32_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_32_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_32_LFInst_1_n2 ), .B(AddRoundKeyOutput[2]), 
        .ZN(Red_SignaltoCheck[129]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_32_LFInst_1_U3  ( .A(AddRoundKeyOutput[3]), 
        .B(AddRoundKeyOutput[0]), .ZN(\Red_ToCheckInst_LFInst_32_LFInst_1_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_32_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_32_LFInst_2_n2 ), .B(AddRoundKeyOutput[1]), 
        .ZN(Red_SignaltoCheck[130]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_32_LFInst_2_U3  ( .A(AddRoundKeyOutput[3]), 
        .B(AddRoundKeyOutput[0]), .ZN(\Red_ToCheckInst_LFInst_32_LFInst_2_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_32_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_32_LFInst_3_n2 ), .B(AddRoundKeyOutput[1]), 
        .ZN(Red_SignaltoCheck[131]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_32_LFInst_3_U3  ( .A(AddRoundKeyOutput[2]), 
        .B(AddRoundKeyOutput[0]), .ZN(\Red_ToCheckInst_LFInst_32_LFInst_3_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_33_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_33_LFInst_0_n2 ), .B(AddRoundKeyOutput[6]), 
        .ZN(Red_SignaltoCheck[132]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_33_LFInst_0_U3  ( .A(AddRoundKeyOutput[7]), 
        .B(AddRoundKeyOutput[5]), .ZN(\Red_ToCheckInst_LFInst_33_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_33_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_33_LFInst_1_n2 ), .B(AddRoundKeyOutput[6]), 
        .ZN(Red_SignaltoCheck[133]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_33_LFInst_1_U3  ( .A(AddRoundKeyOutput[7]), 
        .B(AddRoundKeyOutput[4]), .ZN(\Red_ToCheckInst_LFInst_33_LFInst_1_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_33_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_33_LFInst_2_n2 ), .B(AddRoundKeyOutput[5]), 
        .ZN(Red_SignaltoCheck[134]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_33_LFInst_2_U3  ( .A(AddRoundKeyOutput[7]), 
        .B(AddRoundKeyOutput[4]), .ZN(\Red_ToCheckInst_LFInst_33_LFInst_2_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_33_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_33_LFInst_3_n2 ), .B(AddRoundKeyOutput[5]), 
        .ZN(Red_SignaltoCheck[135]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_33_LFInst_3_U3  ( .A(AddRoundKeyOutput[6]), 
        .B(AddRoundKeyOutput[4]), .ZN(\Red_ToCheckInst_LFInst_33_LFInst_3_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_34_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_34_LFInst_0_n2 ), .B(AddRoundKeyOutput[10]), 
        .ZN(Red_SignaltoCheck[136]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_34_LFInst_0_U3  ( .A(AddRoundKeyOutput[11]), 
        .B(AddRoundKeyOutput[9]), .ZN(\Red_ToCheckInst_LFInst_34_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_34_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_34_LFInst_1_n2 ), .B(AddRoundKeyOutput[10]), 
        .ZN(Red_SignaltoCheck[137]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_34_LFInst_1_U3  ( .A(AddRoundKeyOutput[11]), 
        .B(AddRoundKeyOutput[8]), .ZN(\Red_ToCheckInst_LFInst_34_LFInst_1_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_34_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_34_LFInst_2_n2 ), .B(AddRoundKeyOutput[9]), 
        .ZN(Red_SignaltoCheck[138]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_34_LFInst_2_U3  ( .A(AddRoundKeyOutput[11]), 
        .B(AddRoundKeyOutput[8]), .ZN(\Red_ToCheckInst_LFInst_34_LFInst_2_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_34_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_34_LFInst_3_n2 ), .B(AddRoundKeyOutput[9]), 
        .ZN(Red_SignaltoCheck[139]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_34_LFInst_3_U3  ( .A(AddRoundKeyOutput[10]), 
        .B(AddRoundKeyOutput[8]), .ZN(\Red_ToCheckInst_LFInst_34_LFInst_3_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_35_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_35_LFInst_0_n2 ), .B(AddRoundKeyOutput[14]), 
        .ZN(Red_SignaltoCheck[140]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_35_LFInst_0_U3  ( .A(AddRoundKeyOutput[15]), 
        .B(AddRoundKeyOutput[13]), .ZN(\Red_ToCheckInst_LFInst_35_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_35_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_35_LFInst_1_n2 ), .B(AddRoundKeyOutput[14]), 
        .ZN(Red_SignaltoCheck[141]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_35_LFInst_1_U3  ( .A(AddRoundKeyOutput[15]), 
        .B(AddRoundKeyOutput[12]), .ZN(\Red_ToCheckInst_LFInst_35_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_35_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_35_LFInst_2_n2 ), .B(AddRoundKeyOutput[13]), 
        .ZN(Red_SignaltoCheck[142]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_35_LFInst_2_U3  ( .A(AddRoundKeyOutput[15]), 
        .B(AddRoundKeyOutput[12]), .ZN(\Red_ToCheckInst_LFInst_35_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_35_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_35_LFInst_3_n2 ), .B(AddRoundKeyOutput[13]), 
        .ZN(Red_SignaltoCheck[143]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_35_LFInst_3_U3  ( .A(AddRoundKeyOutput[14]), 
        .B(AddRoundKeyOutput[12]), .ZN(\Red_ToCheckInst_LFInst_35_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_36_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_36_LFInst_0_n2 ), .B(AddRoundKeyOutput[18]), 
        .ZN(Red_SignaltoCheck[144]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_36_LFInst_0_U3  ( .A(AddRoundKeyOutput[19]), 
        .B(AddRoundKeyOutput[17]), .ZN(\Red_ToCheckInst_LFInst_36_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_36_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_36_LFInst_1_n2 ), .B(AddRoundKeyOutput[18]), 
        .ZN(Red_SignaltoCheck[145]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_36_LFInst_1_U3  ( .A(AddRoundKeyOutput[19]), 
        .B(AddRoundKeyOutput[16]), .ZN(\Red_ToCheckInst_LFInst_36_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_36_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_36_LFInst_2_n2 ), .B(AddRoundKeyOutput[17]), 
        .ZN(Red_SignaltoCheck[146]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_36_LFInst_2_U3  ( .A(AddRoundKeyOutput[19]), 
        .B(AddRoundKeyOutput[16]), .ZN(\Red_ToCheckInst_LFInst_36_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_36_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_36_LFInst_3_n2 ), .B(AddRoundKeyOutput[17]), 
        .ZN(Red_SignaltoCheck[147]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_36_LFInst_3_U3  ( .A(AddRoundKeyOutput[18]), 
        .B(AddRoundKeyOutput[16]), .ZN(\Red_ToCheckInst_LFInst_36_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_37_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_37_LFInst_0_n2 ), .B(AddRoundKeyOutput[22]), 
        .ZN(Red_SignaltoCheck[148]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_37_LFInst_0_U3  ( .A(AddRoundKeyOutput[23]), 
        .B(AddRoundKeyOutput[21]), .ZN(\Red_ToCheckInst_LFInst_37_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_37_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_37_LFInst_1_n2 ), .B(AddRoundKeyOutput[22]), 
        .ZN(Red_SignaltoCheck[149]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_37_LFInst_1_U3  ( .A(AddRoundKeyOutput[23]), 
        .B(AddRoundKeyOutput[20]), .ZN(\Red_ToCheckInst_LFInst_37_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_37_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_37_LFInst_2_n2 ), .B(AddRoundKeyOutput[21]), 
        .ZN(Red_SignaltoCheck[150]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_37_LFInst_2_U3  ( .A(AddRoundKeyOutput[23]), 
        .B(AddRoundKeyOutput[20]), .ZN(\Red_ToCheckInst_LFInst_37_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_37_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_37_LFInst_3_n2 ), .B(AddRoundKeyOutput[21]), 
        .ZN(Red_SignaltoCheck[151]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_37_LFInst_3_U3  ( .A(AddRoundKeyOutput[22]), 
        .B(AddRoundKeyOutput[20]), .ZN(\Red_ToCheckInst_LFInst_37_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_38_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_38_LFInst_0_n2 ), .B(AddRoundKeyOutput[26]), 
        .ZN(Red_SignaltoCheck[152]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_38_LFInst_0_U3  ( .A(AddRoundKeyOutput[27]), 
        .B(AddRoundKeyOutput[25]), .ZN(\Red_ToCheckInst_LFInst_38_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_38_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_38_LFInst_1_n2 ), .B(AddRoundKeyOutput[26]), 
        .ZN(Red_SignaltoCheck[153]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_38_LFInst_1_U3  ( .A(AddRoundKeyOutput[27]), 
        .B(AddRoundKeyOutput[24]), .ZN(\Red_ToCheckInst_LFInst_38_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_38_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_38_LFInst_2_n2 ), .B(AddRoundKeyOutput[25]), 
        .ZN(Red_SignaltoCheck[154]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_38_LFInst_2_U3  ( .A(AddRoundKeyOutput[27]), 
        .B(AddRoundKeyOutput[24]), .ZN(\Red_ToCheckInst_LFInst_38_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_38_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_38_LFInst_3_n2 ), .B(AddRoundKeyOutput[25]), 
        .ZN(Red_SignaltoCheck[155]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_38_LFInst_3_U3  ( .A(AddRoundKeyOutput[26]), 
        .B(AddRoundKeyOutput[24]), .ZN(\Red_ToCheckInst_LFInst_38_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_39_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_39_LFInst_0_n2 ), .B(AddRoundKeyOutput[30]), 
        .ZN(Red_SignaltoCheck[156]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_39_LFInst_0_U3  ( .A(AddRoundKeyOutput[31]), 
        .B(AddRoundKeyOutput[29]), .ZN(\Red_ToCheckInst_LFInst_39_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_39_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_39_LFInst_1_n2 ), .B(AddRoundKeyOutput[30]), 
        .ZN(Red_SignaltoCheck[157]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_39_LFInst_1_U3  ( .A(AddRoundKeyOutput[31]), 
        .B(AddRoundKeyOutput[28]), .ZN(\Red_ToCheckInst_LFInst_39_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_39_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_39_LFInst_2_n2 ), .B(AddRoundKeyOutput[29]), 
        .ZN(Red_SignaltoCheck[158]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_39_LFInst_2_U3  ( .A(AddRoundKeyOutput[31]), 
        .B(AddRoundKeyOutput[28]), .ZN(\Red_ToCheckInst_LFInst_39_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_39_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_39_LFInst_3_n2 ), .B(AddRoundKeyOutput[29]), 
        .ZN(Red_SignaltoCheck[159]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_39_LFInst_3_U3  ( .A(AddRoundKeyOutput[30]), 
        .B(AddRoundKeyOutput[28]), .ZN(\Red_ToCheckInst_LFInst_39_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_40_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_40_LFInst_0_n2 ), .B(AddRoundKeyOutput[34]), 
        .ZN(Red_SignaltoCheck[160]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_40_LFInst_0_U3  ( .A(AddRoundKeyOutput[35]), 
        .B(AddRoundKeyOutput[33]), .ZN(\Red_ToCheckInst_LFInst_40_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_40_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_40_LFInst_1_n2 ), .B(AddRoundKeyOutput[34]), 
        .ZN(Red_SignaltoCheck[161]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_40_LFInst_1_U3  ( .A(AddRoundKeyOutput[35]), 
        .B(AddRoundKeyOutput[32]), .ZN(\Red_ToCheckInst_LFInst_40_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_40_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_40_LFInst_2_n2 ), .B(AddRoundKeyOutput[33]), 
        .ZN(Red_SignaltoCheck[162]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_40_LFInst_2_U3  ( .A(AddRoundKeyOutput[35]), 
        .B(AddRoundKeyOutput[32]), .ZN(\Red_ToCheckInst_LFInst_40_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_40_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_40_LFInst_3_n2 ), .B(AddRoundKeyOutput[33]), 
        .ZN(Red_SignaltoCheck[163]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_40_LFInst_3_U3  ( .A(AddRoundKeyOutput[34]), 
        .B(AddRoundKeyOutput[32]), .ZN(\Red_ToCheckInst_LFInst_40_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_41_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_41_LFInst_0_n2 ), .B(AddRoundKeyOutput[38]), 
        .ZN(Red_SignaltoCheck[164]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_41_LFInst_0_U3  ( .A(AddRoundKeyOutput[39]), 
        .B(AddRoundKeyOutput[37]), .ZN(\Red_ToCheckInst_LFInst_41_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_41_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_41_LFInst_1_n2 ), .B(AddRoundKeyOutput[38]), 
        .ZN(Red_SignaltoCheck[165]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_41_LFInst_1_U3  ( .A(AddRoundKeyOutput[39]), 
        .B(AddRoundKeyOutput[36]), .ZN(\Red_ToCheckInst_LFInst_41_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_41_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_41_LFInst_2_n2 ), .B(AddRoundKeyOutput[37]), 
        .ZN(Red_SignaltoCheck[166]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_41_LFInst_2_U3  ( .A(AddRoundKeyOutput[39]), 
        .B(AddRoundKeyOutput[36]), .ZN(\Red_ToCheckInst_LFInst_41_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_41_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_41_LFInst_3_n2 ), .B(AddRoundKeyOutput[37]), 
        .ZN(Red_SignaltoCheck[167]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_41_LFInst_3_U3  ( .A(AddRoundKeyOutput[38]), 
        .B(AddRoundKeyOutput[36]), .ZN(\Red_ToCheckInst_LFInst_41_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_42_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_42_LFInst_0_n2 ), .B(AddRoundKeyOutput[42]), 
        .ZN(Red_SignaltoCheck[168]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_42_LFInst_0_U3  ( .A(AddRoundKeyOutput[43]), 
        .B(AddRoundKeyOutput[41]), .ZN(\Red_ToCheckInst_LFInst_42_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_42_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_42_LFInst_1_n2 ), .B(AddRoundKeyOutput[42]), 
        .ZN(Red_SignaltoCheck[169]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_42_LFInst_1_U3  ( .A(AddRoundKeyOutput[43]), 
        .B(AddRoundKeyOutput[40]), .ZN(\Red_ToCheckInst_LFInst_42_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_42_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_42_LFInst_2_n2 ), .B(AddRoundKeyOutput[41]), 
        .ZN(Red_SignaltoCheck[170]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_42_LFInst_2_U3  ( .A(AddRoundKeyOutput[43]), 
        .B(AddRoundKeyOutput[40]), .ZN(\Red_ToCheckInst_LFInst_42_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_42_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_42_LFInst_3_n2 ), .B(AddRoundKeyOutput[41]), 
        .ZN(Red_SignaltoCheck[171]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_42_LFInst_3_U3  ( .A(AddRoundKeyOutput[42]), 
        .B(AddRoundKeyOutput[40]), .ZN(\Red_ToCheckInst_LFInst_42_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_43_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_43_LFInst_0_n2 ), .B(AddRoundKeyOutput[46]), 
        .ZN(Red_SignaltoCheck[172]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_43_LFInst_0_U3  ( .A(AddRoundKeyOutput[47]), 
        .B(AddRoundKeyOutput[45]), .ZN(\Red_ToCheckInst_LFInst_43_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_43_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_43_LFInst_1_n2 ), .B(AddRoundKeyOutput[46]), 
        .ZN(Red_SignaltoCheck[173]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_43_LFInst_1_U3  ( .A(AddRoundKeyOutput[47]), 
        .B(AddRoundKeyOutput[44]), .ZN(\Red_ToCheckInst_LFInst_43_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_43_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_43_LFInst_2_n2 ), .B(AddRoundKeyOutput[45]), 
        .ZN(Red_SignaltoCheck[174]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_43_LFInst_2_U3  ( .A(AddRoundKeyOutput[47]), 
        .B(AddRoundKeyOutput[44]), .ZN(\Red_ToCheckInst_LFInst_43_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_43_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_43_LFInst_3_n2 ), .B(AddRoundKeyOutput[45]), 
        .ZN(Red_SignaltoCheck[175]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_43_LFInst_3_U3  ( .A(AddRoundKeyOutput[46]), 
        .B(AddRoundKeyOutput[44]), .ZN(\Red_ToCheckInst_LFInst_43_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_44_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_44_LFInst_0_n2 ), .B(AddRoundKeyOutput[50]), 
        .ZN(Red_SignaltoCheck[176]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_44_LFInst_0_U3  ( .A(AddRoundKeyOutput[51]), 
        .B(AddRoundKeyOutput[49]), .ZN(\Red_ToCheckInst_LFInst_44_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_44_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_44_LFInst_1_n2 ), .B(AddRoundKeyOutput[50]), 
        .ZN(Red_SignaltoCheck[177]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_44_LFInst_1_U3  ( .A(AddRoundKeyOutput[51]), 
        .B(AddRoundKeyOutput[48]), .ZN(\Red_ToCheckInst_LFInst_44_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_44_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_44_LFInst_2_n2 ), .B(AddRoundKeyOutput[49]), 
        .ZN(Red_SignaltoCheck[178]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_44_LFInst_2_U3  ( .A(AddRoundKeyOutput[51]), 
        .B(AddRoundKeyOutput[48]), .ZN(\Red_ToCheckInst_LFInst_44_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_44_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_44_LFInst_3_n2 ), .B(AddRoundKeyOutput[49]), 
        .ZN(Red_SignaltoCheck[179]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_44_LFInst_3_U3  ( .A(AddRoundKeyOutput[50]), 
        .B(AddRoundKeyOutput[48]), .ZN(\Red_ToCheckInst_LFInst_44_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_45_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_45_LFInst_0_n2 ), .B(AddRoundKeyOutput[54]), 
        .ZN(Red_SignaltoCheck[180]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_45_LFInst_0_U3  ( .A(AddRoundKeyOutput[55]), 
        .B(AddRoundKeyOutput[53]), .ZN(\Red_ToCheckInst_LFInst_45_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_45_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_45_LFInst_1_n2 ), .B(AddRoundKeyOutput[54]), 
        .ZN(Red_SignaltoCheck[181]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_45_LFInst_1_U3  ( .A(AddRoundKeyOutput[55]), 
        .B(AddRoundKeyOutput[52]), .ZN(\Red_ToCheckInst_LFInst_45_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_45_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_45_LFInst_2_n2 ), .B(AddRoundKeyOutput[53]), 
        .ZN(Red_SignaltoCheck[182]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_45_LFInst_2_U3  ( .A(AddRoundKeyOutput[55]), 
        .B(AddRoundKeyOutput[52]), .ZN(\Red_ToCheckInst_LFInst_45_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_45_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_45_LFInst_3_n2 ), .B(AddRoundKeyOutput[53]), 
        .ZN(Red_SignaltoCheck[183]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_45_LFInst_3_U3  ( .A(AddRoundKeyOutput[54]), 
        .B(AddRoundKeyOutput[52]), .ZN(\Red_ToCheckInst_LFInst_45_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_46_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_46_LFInst_0_n2 ), .B(AddRoundKeyOutput[58]), 
        .ZN(Red_SignaltoCheck[184]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_46_LFInst_0_U3  ( .A(AddRoundKeyOutput[59]), 
        .B(AddRoundKeyOutput[57]), .ZN(\Red_ToCheckInst_LFInst_46_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_46_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_46_LFInst_1_n2 ), .B(AddRoundKeyOutput[58]), 
        .ZN(Red_SignaltoCheck[185]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_46_LFInst_1_U3  ( .A(AddRoundKeyOutput[59]), 
        .B(AddRoundKeyOutput[56]), .ZN(\Red_ToCheckInst_LFInst_46_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_46_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_46_LFInst_2_n2 ), .B(AddRoundKeyOutput[57]), 
        .ZN(Red_SignaltoCheck[186]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_46_LFInst_2_U3  ( .A(AddRoundKeyOutput[59]), 
        .B(AddRoundKeyOutput[56]), .ZN(\Red_ToCheckInst_LFInst_46_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_46_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_46_LFInst_3_n2 ), .B(AddRoundKeyOutput[57]), 
        .ZN(Red_SignaltoCheck[187]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_46_LFInst_3_U3  ( .A(AddRoundKeyOutput[58]), 
        .B(AddRoundKeyOutput[56]), .ZN(\Red_ToCheckInst_LFInst_46_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_47_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_47_LFInst_0_n2 ), .B(AddRoundKeyOutput[62]), 
        .ZN(Red_SignaltoCheck[188]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_47_LFInst_0_U3  ( .A(AddRoundKeyOutput[63]), 
        .B(AddRoundKeyOutput[61]), .ZN(\Red_ToCheckInst_LFInst_47_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_47_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_47_LFInst_1_n2 ), .B(AddRoundKeyOutput[62]), 
        .ZN(Red_SignaltoCheck[189]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_47_LFInst_1_U3  ( .A(AddRoundKeyOutput[63]), 
        .B(AddRoundKeyOutput[60]), .ZN(\Red_ToCheckInst_LFInst_47_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_47_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_47_LFInst_2_n2 ), .B(AddRoundKeyOutput[61]), 
        .ZN(Red_SignaltoCheck[190]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_47_LFInst_2_U3  ( .A(AddRoundKeyOutput[63]), 
        .B(AddRoundKeyOutput[60]), .ZN(\Red_ToCheckInst_LFInst_47_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_47_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_47_LFInst_3_n2 ), .B(AddRoundKeyOutput[61]), 
        .ZN(Red_SignaltoCheck[191]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_47_LFInst_3_U3  ( .A(AddRoundKeyOutput[62]), 
        .B(AddRoundKeyOutput[60]), .ZN(\Red_ToCheckInst_LFInst_47_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_48_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_48_LFInst_0_n2 ), .B(Output[2]), .ZN(
        Red_SignaltoCheck[192]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_48_LFInst_0_U3  ( .A(Output[3]), .B(
        Output[1]), .ZN(\Red_ToCheckInst_LFInst_48_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_48_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_48_LFInst_1_n2 ), .B(Output[2]), .ZN(
        Red_SignaltoCheck[193]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_48_LFInst_1_U3  ( .A(Output[3]), .B(
        Output[0]), .ZN(\Red_ToCheckInst_LFInst_48_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_48_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_48_LFInst_2_n2 ), .B(Output[1]), .ZN(
        Red_SignaltoCheck[194]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_48_LFInst_2_U3  ( .A(Output[3]), .B(
        Output[0]), .ZN(\Red_ToCheckInst_LFInst_48_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_48_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_48_LFInst_3_n2 ), .B(Output[1]), .ZN(
        Red_SignaltoCheck[195]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_48_LFInst_3_U3  ( .A(Output[2]), .B(
        Output[0]), .ZN(\Red_ToCheckInst_LFInst_48_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_49_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_49_LFInst_0_n2 ), .B(Output[6]), .ZN(
        Red_SignaltoCheck[196]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_49_LFInst_0_U3  ( .A(Output[7]), .B(
        Output[5]), .ZN(\Red_ToCheckInst_LFInst_49_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_49_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_49_LFInst_1_n2 ), .B(Output[6]), .ZN(
        Red_SignaltoCheck[197]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_49_LFInst_1_U3  ( .A(Output[7]), .B(
        Output[4]), .ZN(\Red_ToCheckInst_LFInst_49_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_49_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_49_LFInst_2_n2 ), .B(Output[5]), .ZN(
        Red_SignaltoCheck[198]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_49_LFInst_2_U3  ( .A(Output[7]), .B(
        Output[4]), .ZN(\Red_ToCheckInst_LFInst_49_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_49_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_49_LFInst_3_n2 ), .B(Output[5]), .ZN(
        Red_SignaltoCheck[199]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_49_LFInst_3_U3  ( .A(Output[6]), .B(
        Output[4]), .ZN(\Red_ToCheckInst_LFInst_49_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_50_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_50_LFInst_0_n2 ), .B(Output[10]), .ZN(
        Red_SignaltoCheck[200]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_50_LFInst_0_U3  ( .A(Output[11]), .B(
        Output[9]), .ZN(\Red_ToCheckInst_LFInst_50_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_50_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_50_LFInst_1_n2 ), .B(Output[10]), .ZN(
        Red_SignaltoCheck[201]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_50_LFInst_1_U3  ( .A(Output[11]), .B(
        Output[8]), .ZN(\Red_ToCheckInst_LFInst_50_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_50_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_50_LFInst_2_n2 ), .B(Output[9]), .ZN(
        Red_SignaltoCheck[202]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_50_LFInst_2_U3  ( .A(Output[11]), .B(
        Output[8]), .ZN(\Red_ToCheckInst_LFInst_50_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_50_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_50_LFInst_3_n2 ), .B(Output[9]), .ZN(
        Red_SignaltoCheck[203]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_50_LFInst_3_U3  ( .A(Output[10]), .B(
        Output[8]), .ZN(\Red_ToCheckInst_LFInst_50_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_51_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_51_LFInst_0_n2 ), .B(Output[14]), .ZN(
        Red_SignaltoCheck[204]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_51_LFInst_0_U3  ( .A(Output[15]), .B(
        Output[13]), .ZN(\Red_ToCheckInst_LFInst_51_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_51_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_51_LFInst_1_n2 ), .B(Output[14]), .ZN(
        Red_SignaltoCheck[205]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_51_LFInst_1_U3  ( .A(Output[15]), .B(
        Output[12]), .ZN(\Red_ToCheckInst_LFInst_51_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_51_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_51_LFInst_2_n2 ), .B(Output[13]), .ZN(
        Red_SignaltoCheck[206]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_51_LFInst_2_U3  ( .A(Output[15]), .B(
        Output[12]), .ZN(\Red_ToCheckInst_LFInst_51_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_51_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_51_LFInst_3_n2 ), .B(Output[13]), .ZN(
        Red_SignaltoCheck[207]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_51_LFInst_3_U3  ( .A(Output[14]), .B(
        Output[12]), .ZN(\Red_ToCheckInst_LFInst_51_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_52_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_52_LFInst_0_n2 ), .B(Output[18]), .ZN(
        Red_SignaltoCheck[208]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_52_LFInst_0_U3  ( .A(Output[19]), .B(
        Output[17]), .ZN(\Red_ToCheckInst_LFInst_52_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_52_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_52_LFInst_1_n2 ), .B(Output[18]), .ZN(
        Red_SignaltoCheck[209]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_52_LFInst_1_U3  ( .A(Output[19]), .B(
        Output[16]), .ZN(\Red_ToCheckInst_LFInst_52_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_52_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_52_LFInst_2_n2 ), .B(Output[17]), .ZN(
        Red_SignaltoCheck[210]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_52_LFInst_2_U3  ( .A(Output[19]), .B(
        Output[16]), .ZN(\Red_ToCheckInst_LFInst_52_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_52_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_52_LFInst_3_n2 ), .B(Output[17]), .ZN(
        Red_SignaltoCheck[211]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_52_LFInst_3_U3  ( .A(Output[18]), .B(
        Output[16]), .ZN(\Red_ToCheckInst_LFInst_52_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_53_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_53_LFInst_0_n2 ), .B(Output[22]), .ZN(
        Red_SignaltoCheck[212]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_53_LFInst_0_U3  ( .A(Output[23]), .B(
        Output[21]), .ZN(\Red_ToCheckInst_LFInst_53_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_53_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_53_LFInst_1_n2 ), .B(Output[22]), .ZN(
        Red_SignaltoCheck[213]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_53_LFInst_1_U3  ( .A(Output[23]), .B(
        Output[20]), .ZN(\Red_ToCheckInst_LFInst_53_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_53_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_53_LFInst_2_n2 ), .B(Output[21]), .ZN(
        Red_SignaltoCheck[214]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_53_LFInst_2_U3  ( .A(Output[23]), .B(
        Output[20]), .ZN(\Red_ToCheckInst_LFInst_53_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_53_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_53_LFInst_3_n2 ), .B(Output[21]), .ZN(
        Red_SignaltoCheck[215]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_53_LFInst_3_U3  ( .A(Output[22]), .B(
        Output[20]), .ZN(\Red_ToCheckInst_LFInst_53_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_54_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_54_LFInst_0_n2 ), .B(Output[26]), .ZN(
        Red_SignaltoCheck[216]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_54_LFInst_0_U3  ( .A(Output[27]), .B(
        Output[25]), .ZN(\Red_ToCheckInst_LFInst_54_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_54_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_54_LFInst_1_n2 ), .B(Output[26]), .ZN(
        Red_SignaltoCheck[217]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_54_LFInst_1_U3  ( .A(Output[27]), .B(
        Output[24]), .ZN(\Red_ToCheckInst_LFInst_54_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_54_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_54_LFInst_2_n2 ), .B(Output[25]), .ZN(
        Red_SignaltoCheck[218]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_54_LFInst_2_U3  ( .A(Output[27]), .B(
        Output[24]), .ZN(\Red_ToCheckInst_LFInst_54_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_54_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_54_LFInst_3_n2 ), .B(Output[25]), .ZN(
        Red_SignaltoCheck[219]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_54_LFInst_3_U3  ( .A(Output[26]), .B(
        Output[24]), .ZN(\Red_ToCheckInst_LFInst_54_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_55_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_55_LFInst_0_n2 ), .B(Output[30]), .ZN(
        Red_SignaltoCheck[220]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_55_LFInst_0_U3  ( .A(Output[31]), .B(
        Output[29]), .ZN(\Red_ToCheckInst_LFInst_55_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_55_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_55_LFInst_1_n2 ), .B(Output[30]), .ZN(
        Red_SignaltoCheck[221]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_55_LFInst_1_U3  ( .A(Output[31]), .B(
        Output[28]), .ZN(\Red_ToCheckInst_LFInst_55_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_55_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_55_LFInst_2_n2 ), .B(Output[29]), .ZN(
        Red_SignaltoCheck[222]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_55_LFInst_2_U3  ( .A(Output[31]), .B(
        Output[28]), .ZN(\Red_ToCheckInst_LFInst_55_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_55_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_55_LFInst_3_n2 ), .B(Output[29]), .ZN(
        Red_SignaltoCheck[223]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_55_LFInst_3_U3  ( .A(Output[30]), .B(
        Output[28]), .ZN(\Red_ToCheckInst_LFInst_55_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_56_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_56_LFInst_0_n2 ), .B(Output[34]), .ZN(
        Red_SignaltoCheck[224]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_56_LFInst_0_U3  ( .A(Output[35]), .B(
        Output[33]), .ZN(\Red_ToCheckInst_LFInst_56_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_56_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_56_LFInst_1_n2 ), .B(Output[34]), .ZN(
        Red_SignaltoCheck[225]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_56_LFInst_1_U3  ( .A(Output[35]), .B(
        Output[32]), .ZN(\Red_ToCheckInst_LFInst_56_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_56_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_56_LFInst_2_n2 ), .B(Output[33]), .ZN(
        Red_SignaltoCheck[226]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_56_LFInst_2_U3  ( .A(Output[35]), .B(
        Output[32]), .ZN(\Red_ToCheckInst_LFInst_56_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_56_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_56_LFInst_3_n2 ), .B(Output[33]), .ZN(
        Red_SignaltoCheck[227]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_56_LFInst_3_U3  ( .A(Output[34]), .B(
        Output[32]), .ZN(\Red_ToCheckInst_LFInst_56_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_57_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_57_LFInst_0_n2 ), .B(Output[38]), .ZN(
        Red_SignaltoCheck[228]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_57_LFInst_0_U3  ( .A(Output[39]), .B(
        Output[37]), .ZN(\Red_ToCheckInst_LFInst_57_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_57_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_57_LFInst_1_n2 ), .B(Output[38]), .ZN(
        Red_SignaltoCheck[229]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_57_LFInst_1_U3  ( .A(Output[39]), .B(
        Output[36]), .ZN(\Red_ToCheckInst_LFInst_57_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_57_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_57_LFInst_2_n2 ), .B(Output[37]), .ZN(
        Red_SignaltoCheck[230]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_57_LFInst_2_U3  ( .A(Output[39]), .B(
        Output[36]), .ZN(\Red_ToCheckInst_LFInst_57_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_57_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_57_LFInst_3_n2 ), .B(Output[37]), .ZN(
        Red_SignaltoCheck[231]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_57_LFInst_3_U3  ( .A(Output[38]), .B(
        Output[36]), .ZN(\Red_ToCheckInst_LFInst_57_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_58_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_58_LFInst_0_n2 ), .B(Output[42]), .ZN(
        Red_SignaltoCheck[232]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_58_LFInst_0_U3  ( .A(Output[43]), .B(
        Output[41]), .ZN(\Red_ToCheckInst_LFInst_58_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_58_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_58_LFInst_1_n2 ), .B(Output[42]), .ZN(
        Red_SignaltoCheck[233]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_58_LFInst_1_U3  ( .A(Output[43]), .B(
        Output[40]), .ZN(\Red_ToCheckInst_LFInst_58_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_58_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_58_LFInst_2_n2 ), .B(Output[41]), .ZN(
        Red_SignaltoCheck[234]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_58_LFInst_2_U3  ( .A(Output[43]), .B(
        Output[40]), .ZN(\Red_ToCheckInst_LFInst_58_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_58_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_58_LFInst_3_n2 ), .B(Output[41]), .ZN(
        Red_SignaltoCheck[235]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_58_LFInst_3_U3  ( .A(Output[42]), .B(
        Output[40]), .ZN(\Red_ToCheckInst_LFInst_58_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_59_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_59_LFInst_0_n2 ), .B(Output[46]), .ZN(
        Red_SignaltoCheck[236]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_59_LFInst_0_U3  ( .A(Output[47]), .B(
        Output[45]), .ZN(\Red_ToCheckInst_LFInst_59_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_59_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_59_LFInst_1_n2 ), .B(Output[46]), .ZN(
        Red_SignaltoCheck[237]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_59_LFInst_1_U3  ( .A(Output[47]), .B(
        Output[44]), .ZN(\Red_ToCheckInst_LFInst_59_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_59_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_59_LFInst_2_n2 ), .B(Output[45]), .ZN(
        Red_SignaltoCheck[238]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_59_LFInst_2_U3  ( .A(Output[47]), .B(
        Output[44]), .ZN(\Red_ToCheckInst_LFInst_59_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_59_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_59_LFInst_3_n2 ), .B(Output[45]), .ZN(
        Red_SignaltoCheck[239]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_59_LFInst_3_U3  ( .A(Output[46]), .B(
        Output[44]), .ZN(\Red_ToCheckInst_LFInst_59_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_60_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_60_LFInst_0_n2 ), .B(Output[50]), .ZN(
        Red_SignaltoCheck[240]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_60_LFInst_0_U3  ( .A(Output[51]), .B(
        Output[49]), .ZN(\Red_ToCheckInst_LFInst_60_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_60_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_60_LFInst_1_n2 ), .B(Output[50]), .ZN(
        Red_SignaltoCheck[241]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_60_LFInst_1_U3  ( .A(Output[51]), .B(
        Output[48]), .ZN(\Red_ToCheckInst_LFInst_60_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_60_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_60_LFInst_2_n2 ), .B(Output[49]), .ZN(
        Red_SignaltoCheck[242]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_60_LFInst_2_U3  ( .A(Output[51]), .B(
        Output[48]), .ZN(\Red_ToCheckInst_LFInst_60_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_60_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_60_LFInst_3_n2 ), .B(Output[49]), .ZN(
        Red_SignaltoCheck[243]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_60_LFInst_3_U3  ( .A(Output[50]), .B(
        Output[48]), .ZN(\Red_ToCheckInst_LFInst_60_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_61_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_61_LFInst_0_n2 ), .B(Output[54]), .ZN(
        Red_SignaltoCheck[244]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_61_LFInst_0_U3  ( .A(Output[55]), .B(
        Output[53]), .ZN(\Red_ToCheckInst_LFInst_61_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_61_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_61_LFInst_1_n2 ), .B(Output[54]), .ZN(
        Red_SignaltoCheck[245]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_61_LFInst_1_U3  ( .A(Output[55]), .B(
        Output[52]), .ZN(\Red_ToCheckInst_LFInst_61_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_61_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_61_LFInst_2_n2 ), .B(Output[53]), .ZN(
        Red_SignaltoCheck[246]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_61_LFInst_2_U3  ( .A(Output[55]), .B(
        Output[52]), .ZN(\Red_ToCheckInst_LFInst_61_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_61_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_61_LFInst_3_n2 ), .B(Output[53]), .ZN(
        Red_SignaltoCheck[247]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_61_LFInst_3_U3  ( .A(Output[54]), .B(
        Output[52]), .ZN(\Red_ToCheckInst_LFInst_61_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_62_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_62_LFInst_0_n2 ), .B(Output[58]), .ZN(
        Red_SignaltoCheck[248]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_62_LFInst_0_U3  ( .A(Output[59]), .B(
        Output[57]), .ZN(\Red_ToCheckInst_LFInst_62_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_62_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_62_LFInst_1_n2 ), .B(Output[58]), .ZN(
        Red_SignaltoCheck[249]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_62_LFInst_1_U3  ( .A(Output[59]), .B(
        Output[56]), .ZN(\Red_ToCheckInst_LFInst_62_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_62_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_62_LFInst_2_n2 ), .B(Output[57]), .ZN(
        Red_SignaltoCheck[250]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_62_LFInst_2_U3  ( .A(Output[59]), .B(
        Output[56]), .ZN(\Red_ToCheckInst_LFInst_62_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_62_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_62_LFInst_3_n2 ), .B(Output[57]), .ZN(
        Red_SignaltoCheck[251]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_62_LFInst_3_U3  ( .A(Output[58]), .B(
        Output[56]), .ZN(\Red_ToCheckInst_LFInst_62_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_63_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_63_LFInst_0_n2 ), .B(Output[62]), .ZN(
        Red_SignaltoCheck[252]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_63_LFInst_0_U3  ( .A(Output[63]), .B(
        Output[61]), .ZN(\Red_ToCheckInst_LFInst_63_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_63_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_63_LFInst_1_n2 ), .B(Output[62]), .ZN(
        Red_SignaltoCheck[253]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_63_LFInst_1_U3  ( .A(Output[63]), .B(
        Output[60]), .ZN(\Red_ToCheckInst_LFInst_63_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_63_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_63_LFInst_2_n2 ), .B(Output[61]), .ZN(
        Red_SignaltoCheck[254]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_63_LFInst_2_U3  ( .A(Output[63]), .B(
        Output[60]), .ZN(\Red_ToCheckInst_LFInst_63_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_63_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_63_LFInst_3_n2 ), .B(Output[61]), .ZN(
        Red_SignaltoCheck[255]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_63_LFInst_3_U3  ( .A(Output[62]), .B(
        Output[60]), .ZN(\Red_ToCheckInst_LFInst_63_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_64_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_64_LFInst_0_n2 ), .B(PermutationOutput3[62]), 
        .ZN(Red_SignaltoCheck[256]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_64_LFInst_0_U3  ( .A(PermutationOutput3[63]), .B(PermutationOutput3[61]), .ZN(\Red_ToCheckInst_LFInst_64_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_64_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_64_LFInst_1_n2 ), .B(PermutationOutput3[62]), 
        .ZN(Red_SignaltoCheck[257]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_64_LFInst_1_U3  ( .A(PermutationOutput3[63]), .B(PermutationOutput3[60]), .ZN(\Red_ToCheckInst_LFInst_64_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_64_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_64_LFInst_2_n2 ), .B(PermutationOutput3[61]), 
        .ZN(Red_SignaltoCheck[258]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_64_LFInst_2_U3  ( .A(PermutationOutput3[63]), .B(PermutationOutput3[60]), .ZN(\Red_ToCheckInst_LFInst_64_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_64_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_64_LFInst_3_n2 ), .B(PermutationOutput3[61]), 
        .ZN(Red_SignaltoCheck[259]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_64_LFInst_3_U3  ( .A(PermutationOutput3[62]), .B(PermutationOutput3[60]), .ZN(\Red_ToCheckInst_LFInst_64_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_65_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_65_LFInst_0_n2 ), .B(PermutationOutput3[50]), 
        .ZN(Red_SignaltoCheck[260]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_65_LFInst_0_U3  ( .A(PermutationOutput3[51]), .B(PermutationOutput3[49]), .ZN(\Red_ToCheckInst_LFInst_65_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_65_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_65_LFInst_1_n2 ), .B(PermutationOutput3[50]), 
        .ZN(Red_SignaltoCheck[261]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_65_LFInst_1_U3  ( .A(PermutationOutput3[51]), .B(PermutationOutput3[48]), .ZN(\Red_ToCheckInst_LFInst_65_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_65_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_65_LFInst_2_n2 ), .B(PermutationOutput3[49]), 
        .ZN(Red_SignaltoCheck[262]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_65_LFInst_2_U3  ( .A(PermutationOutput3[51]), .B(PermutationOutput3[48]), .ZN(\Red_ToCheckInst_LFInst_65_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_65_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_65_LFInst_3_n2 ), .B(PermutationOutput3[49]), 
        .ZN(Red_SignaltoCheck[263]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_65_LFInst_3_U3  ( .A(PermutationOutput3[50]), .B(PermutationOutput3[48]), .ZN(\Red_ToCheckInst_LFInst_65_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_66_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_66_LFInst_0_n2 ), .B(PermutationOutput3[54]), 
        .ZN(Red_SignaltoCheck[264]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_66_LFInst_0_U3  ( .A(PermutationOutput3[55]), .B(PermutationOutput3[53]), .ZN(\Red_ToCheckInst_LFInst_66_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_66_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_66_LFInst_1_n2 ), .B(PermutationOutput3[54]), 
        .ZN(Red_SignaltoCheck[265]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_66_LFInst_1_U3  ( .A(PermutationOutput3[55]), .B(PermutationOutput3[52]), .ZN(\Red_ToCheckInst_LFInst_66_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_66_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_66_LFInst_2_n2 ), .B(PermutationOutput3[53]), 
        .ZN(Red_SignaltoCheck[266]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_66_LFInst_2_U3  ( .A(PermutationOutput3[55]), .B(PermutationOutput3[52]), .ZN(\Red_ToCheckInst_LFInst_66_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_66_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_66_LFInst_3_n2 ), .B(PermutationOutput3[53]), 
        .ZN(Red_SignaltoCheck[267]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_66_LFInst_3_U3  ( .A(PermutationOutput3[54]), .B(PermutationOutput3[52]), .ZN(\Red_ToCheckInst_LFInst_66_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_67_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_67_LFInst_0_n2 ), .B(PermutationOutput3[58]), 
        .ZN(Red_SignaltoCheck[268]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_67_LFInst_0_U3  ( .A(PermutationOutput3[59]), .B(PermutationOutput3[57]), .ZN(\Red_ToCheckInst_LFInst_67_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_67_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_67_LFInst_1_n2 ), .B(PermutationOutput3[58]), 
        .ZN(Red_SignaltoCheck[269]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_67_LFInst_1_U3  ( .A(PermutationOutput3[59]), .B(PermutationOutput3[56]), .ZN(\Red_ToCheckInst_LFInst_67_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_67_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_67_LFInst_2_n2 ), .B(PermutationOutput3[57]), 
        .ZN(Red_SignaltoCheck[270]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_67_LFInst_2_U3  ( .A(PermutationOutput3[59]), .B(PermutationOutput3[56]), .ZN(\Red_ToCheckInst_LFInst_67_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_67_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_67_LFInst_3_n2 ), .B(PermutationOutput3[57]), 
        .ZN(Red_SignaltoCheck[271]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_67_LFInst_3_U3  ( .A(PermutationOutput3[58]), .B(PermutationOutput3[56]), .ZN(\Red_ToCheckInst_LFInst_67_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_68_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_68_LFInst_0_n2 ), .B(PermutationOutput3[34]), 
        .ZN(Red_SignaltoCheck[272]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_68_LFInst_0_U3  ( .A(PermutationOutput3[35]), .B(PermutationOutput3[33]), .ZN(\Red_ToCheckInst_LFInst_68_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_68_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_68_LFInst_1_n2 ), .B(PermutationOutput3[34]), 
        .ZN(Red_SignaltoCheck[273]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_68_LFInst_1_U3  ( .A(PermutationOutput3[35]), .B(PermutationOutput3[32]), .ZN(\Red_ToCheckInst_LFInst_68_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_68_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_68_LFInst_2_n2 ), .B(PermutationOutput3[33]), 
        .ZN(Red_SignaltoCheck[274]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_68_LFInst_2_U3  ( .A(PermutationOutput3[35]), .B(PermutationOutput3[32]), .ZN(\Red_ToCheckInst_LFInst_68_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_68_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_68_LFInst_3_n2 ), .B(PermutationOutput3[33]), 
        .ZN(Red_SignaltoCheck[275]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_68_LFInst_3_U3  ( .A(PermutationOutput3[34]), .B(PermutationOutput3[32]), .ZN(\Red_ToCheckInst_LFInst_68_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_69_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_69_LFInst_0_n2 ), .B(PermutationOutput3[46]), 
        .ZN(Red_SignaltoCheck[276]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_69_LFInst_0_U3  ( .A(PermutationOutput3[47]), .B(PermutationOutput3[45]), .ZN(\Red_ToCheckInst_LFInst_69_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_69_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_69_LFInst_1_n2 ), .B(PermutationOutput3[46]), 
        .ZN(Red_SignaltoCheck[277]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_69_LFInst_1_U3  ( .A(PermutationOutput3[47]), .B(PermutationOutput3[44]), .ZN(\Red_ToCheckInst_LFInst_69_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_69_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_69_LFInst_2_n2 ), .B(PermutationOutput3[45]), 
        .ZN(Red_SignaltoCheck[278]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_69_LFInst_2_U3  ( .A(PermutationOutput3[47]), .B(PermutationOutput3[44]), .ZN(\Red_ToCheckInst_LFInst_69_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_69_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_69_LFInst_3_n2 ), .B(PermutationOutput3[45]), 
        .ZN(Red_SignaltoCheck[279]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_69_LFInst_3_U3  ( .A(PermutationOutput3[46]), .B(PermutationOutput3[44]), .ZN(\Red_ToCheckInst_LFInst_69_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_70_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_70_LFInst_0_n2 ), .B(PermutationOutput3[42]), 
        .ZN(Red_SignaltoCheck[280]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_70_LFInst_0_U3  ( .A(PermutationOutput3[43]), .B(PermutationOutput3[41]), .ZN(\Red_ToCheckInst_LFInst_70_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_70_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_70_LFInst_1_n2 ), .B(PermutationOutput3[42]), 
        .ZN(Red_SignaltoCheck[281]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_70_LFInst_1_U3  ( .A(PermutationOutput3[43]), .B(PermutationOutput3[40]), .ZN(\Red_ToCheckInst_LFInst_70_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_70_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_70_LFInst_2_n2 ), .B(PermutationOutput3[41]), 
        .ZN(Red_SignaltoCheck[282]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_70_LFInst_2_U3  ( .A(PermutationOutput3[43]), .B(PermutationOutput3[40]), .ZN(\Red_ToCheckInst_LFInst_70_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_70_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_70_LFInst_3_n2 ), .B(PermutationOutput3[41]), 
        .ZN(Red_SignaltoCheck[283]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_70_LFInst_3_U3  ( .A(PermutationOutput3[42]), .B(PermutationOutput3[40]), .ZN(\Red_ToCheckInst_LFInst_70_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_71_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_71_LFInst_0_n2 ), .B(PermutationOutput3[38]), 
        .ZN(Red_SignaltoCheck[284]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_71_LFInst_0_U3  ( .A(PermutationOutput3[39]), .B(PermutationOutput3[37]), .ZN(\Red_ToCheckInst_LFInst_71_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_71_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_71_LFInst_1_n2 ), .B(PermutationOutput3[38]), 
        .ZN(Red_SignaltoCheck[285]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_71_LFInst_1_U3  ( .A(PermutationOutput3[39]), .B(PermutationOutput3[36]), .ZN(\Red_ToCheckInst_LFInst_71_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_71_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_71_LFInst_2_n2 ), .B(PermutationOutput3[37]), 
        .ZN(Red_SignaltoCheck[286]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_71_LFInst_2_U3  ( .A(PermutationOutput3[39]), .B(PermutationOutput3[36]), .ZN(\Red_ToCheckInst_LFInst_71_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_71_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_71_LFInst_3_n2 ), .B(PermutationOutput3[37]), 
        .ZN(Red_SignaltoCheck[287]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_71_LFInst_3_U3  ( .A(PermutationOutput3[38]), .B(PermutationOutput3[36]), .ZN(\Red_ToCheckInst_LFInst_71_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_72_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_72_LFInst_0_n2 ), .B(PermutationOutput3[18]), 
        .ZN(Red_SignaltoCheck[288]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_72_LFInst_0_U3  ( .A(PermutationOutput3[19]), .B(PermutationOutput3[17]), .ZN(\Red_ToCheckInst_LFInst_72_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_72_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_72_LFInst_1_n2 ), .B(PermutationOutput3[18]), 
        .ZN(Red_SignaltoCheck[289]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_72_LFInst_1_U3  ( .A(PermutationOutput3[19]), .B(PermutationOutput3[16]), .ZN(\Red_ToCheckInst_LFInst_72_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_72_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_72_LFInst_2_n2 ), .B(PermutationOutput3[17]), 
        .ZN(Red_SignaltoCheck[290]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_72_LFInst_2_U3  ( .A(PermutationOutput3[19]), .B(PermutationOutput3[16]), .ZN(\Red_ToCheckInst_LFInst_72_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_72_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_72_LFInst_3_n2 ), .B(PermutationOutput3[17]), 
        .ZN(Red_SignaltoCheck[291]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_72_LFInst_3_U3  ( .A(PermutationOutput3[18]), .B(PermutationOutput3[16]), .ZN(\Red_ToCheckInst_LFInst_72_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_73_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_73_LFInst_0_n2 ), .B(PermutationOutput3[30]), 
        .ZN(Red_SignaltoCheck[292]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_73_LFInst_0_U3  ( .A(PermutationOutput3[31]), .B(PermutationOutput3[29]), .ZN(\Red_ToCheckInst_LFInst_73_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_73_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_73_LFInst_1_n2 ), .B(PermutationOutput3[30]), 
        .ZN(Red_SignaltoCheck[293]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_73_LFInst_1_U3  ( .A(PermutationOutput3[31]), .B(PermutationOutput3[28]), .ZN(\Red_ToCheckInst_LFInst_73_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_73_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_73_LFInst_2_n2 ), .B(PermutationOutput3[29]), 
        .ZN(Red_SignaltoCheck[294]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_73_LFInst_2_U3  ( .A(PermutationOutput3[31]), .B(PermutationOutput3[28]), .ZN(\Red_ToCheckInst_LFInst_73_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_73_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_73_LFInst_3_n2 ), .B(PermutationOutput3[29]), 
        .ZN(Red_SignaltoCheck[295]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_73_LFInst_3_U3  ( .A(PermutationOutput3[30]), .B(PermutationOutput3[28]), .ZN(\Red_ToCheckInst_LFInst_73_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_74_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_74_LFInst_0_n2 ), .B(PermutationOutput3[26]), 
        .ZN(Red_SignaltoCheck[296]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_74_LFInst_0_U3  ( .A(PermutationOutput3[27]), .B(PermutationOutput3[25]), .ZN(\Red_ToCheckInst_LFInst_74_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_74_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_74_LFInst_1_n2 ), .B(PermutationOutput3[26]), 
        .ZN(Red_SignaltoCheck[297]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_74_LFInst_1_U3  ( .A(PermutationOutput3[27]), .B(PermutationOutput3[24]), .ZN(\Red_ToCheckInst_LFInst_74_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_74_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_74_LFInst_2_n2 ), .B(PermutationOutput3[25]), 
        .ZN(Red_SignaltoCheck[298]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_74_LFInst_2_U3  ( .A(PermutationOutput3[27]), .B(PermutationOutput3[24]), .ZN(\Red_ToCheckInst_LFInst_74_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_74_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_74_LFInst_3_n2 ), .B(PermutationOutput3[25]), 
        .ZN(Red_SignaltoCheck[299]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_74_LFInst_3_U3  ( .A(PermutationOutput3[26]), .B(PermutationOutput3[24]), .ZN(\Red_ToCheckInst_LFInst_74_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_75_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_75_LFInst_0_n2 ), .B(PermutationOutput3[22]), 
        .ZN(Red_SignaltoCheck[300]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_75_LFInst_0_U3  ( .A(PermutationOutput3[23]), .B(PermutationOutput3[21]), .ZN(\Red_ToCheckInst_LFInst_75_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_75_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_75_LFInst_1_n2 ), .B(PermutationOutput3[22]), 
        .ZN(Red_SignaltoCheck[301]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_75_LFInst_1_U3  ( .A(PermutationOutput3[23]), .B(PermutationOutput3[20]), .ZN(\Red_ToCheckInst_LFInst_75_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_75_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_75_LFInst_2_n2 ), .B(PermutationOutput3[21]), 
        .ZN(Red_SignaltoCheck[302]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_75_LFInst_2_U3  ( .A(PermutationOutput3[23]), .B(PermutationOutput3[20]), .ZN(\Red_ToCheckInst_LFInst_75_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_75_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_75_LFInst_3_n2 ), .B(PermutationOutput3[21]), 
        .ZN(Red_SignaltoCheck[303]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_75_LFInst_3_U3  ( .A(PermutationOutput3[22]), .B(PermutationOutput3[20]), .ZN(\Red_ToCheckInst_LFInst_75_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_76_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_76_LFInst_0_n2 ), .B(PermutationOutput3[6]), 
        .ZN(Red_SignaltoCheck[304]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_76_LFInst_0_U3  ( .A(PermutationOutput3[7]), 
        .B(PermutationOutput3[5]), .ZN(\Red_ToCheckInst_LFInst_76_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_76_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_76_LFInst_1_n2 ), .B(PermutationOutput3[6]), 
        .ZN(Red_SignaltoCheck[305]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_76_LFInst_1_U3  ( .A(PermutationOutput3[7]), 
        .B(PermutationOutput3[4]), .ZN(\Red_ToCheckInst_LFInst_76_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_76_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_76_LFInst_2_n2 ), .B(PermutationOutput3[5]), 
        .ZN(Red_SignaltoCheck[306]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_76_LFInst_2_U3  ( .A(PermutationOutput3[7]), 
        .B(PermutationOutput3[4]), .ZN(\Red_ToCheckInst_LFInst_76_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_76_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_76_LFInst_3_n2 ), .B(PermutationOutput3[5]), 
        .ZN(Red_SignaltoCheck[307]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_76_LFInst_3_U3  ( .A(PermutationOutput3[6]), 
        .B(PermutationOutput3[4]), .ZN(\Red_ToCheckInst_LFInst_76_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_77_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_77_LFInst_0_n2 ), .B(PermutationOutput3[10]), 
        .ZN(Red_SignaltoCheck[308]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_77_LFInst_0_U3  ( .A(PermutationOutput3[11]), .B(PermutationOutput3[9]), .ZN(\Red_ToCheckInst_LFInst_77_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_77_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_77_LFInst_1_n2 ), .B(PermutationOutput3[10]), 
        .ZN(Red_SignaltoCheck[309]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_77_LFInst_1_U3  ( .A(PermutationOutput3[11]), .B(PermutationOutput3[8]), .ZN(\Red_ToCheckInst_LFInst_77_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_77_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_77_LFInst_2_n2 ), .B(PermutationOutput3[9]), 
        .ZN(Red_SignaltoCheck[310]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_77_LFInst_2_U3  ( .A(PermutationOutput3[11]), .B(PermutationOutput3[8]), .ZN(\Red_ToCheckInst_LFInst_77_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_77_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_77_LFInst_3_n2 ), .B(PermutationOutput3[9]), 
        .ZN(Red_SignaltoCheck[311]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_77_LFInst_3_U3  ( .A(PermutationOutput3[10]), .B(PermutationOutput3[8]), .ZN(\Red_ToCheckInst_LFInst_77_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_78_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_78_LFInst_0_n2 ), .B(PermutationOutput3[14]), 
        .ZN(Red_SignaltoCheck[312]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_78_LFInst_0_U3  ( .A(PermutationOutput3[15]), .B(PermutationOutput3[13]), .ZN(\Red_ToCheckInst_LFInst_78_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_78_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_78_LFInst_1_n2 ), .B(PermutationOutput3[14]), 
        .ZN(Red_SignaltoCheck[313]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_78_LFInst_1_U3  ( .A(PermutationOutput3[15]), .B(PermutationOutput3[12]), .ZN(\Red_ToCheckInst_LFInst_78_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_78_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_78_LFInst_2_n2 ), .B(PermutationOutput3[13]), 
        .ZN(Red_SignaltoCheck[314]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_78_LFInst_2_U3  ( .A(PermutationOutput3[15]), .B(PermutationOutput3[12]), .ZN(\Red_ToCheckInst_LFInst_78_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_78_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_78_LFInst_3_n2 ), .B(PermutationOutput3[13]), 
        .ZN(Red_SignaltoCheck[315]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_78_LFInst_3_U3  ( .A(PermutationOutput3[14]), .B(PermutationOutput3[12]), .ZN(\Red_ToCheckInst_LFInst_78_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_79_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_79_LFInst_0_n2 ), .B(PermutationOutput3[2]), 
        .ZN(Red_SignaltoCheck[316]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_79_LFInst_0_U3  ( .A(PermutationOutput3[3]), 
        .B(PermutationOutput3[1]), .ZN(\Red_ToCheckInst_LFInst_79_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_79_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_79_LFInst_1_n2 ), .B(PermutationOutput3[2]), 
        .ZN(Red_SignaltoCheck[317]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_79_LFInst_1_U3  ( .A(PermutationOutput3[3]), 
        .B(PermutationOutput3[0]), .ZN(\Red_ToCheckInst_LFInst_79_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_79_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_79_LFInst_2_n2 ), .B(PermutationOutput3[1]), 
        .ZN(Red_SignaltoCheck[318]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_79_LFInst_2_U3  ( .A(PermutationOutput3[3]), 
        .B(PermutationOutput3[0]), .ZN(\Red_ToCheckInst_LFInst_79_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_79_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_79_LFInst_3_n2 ), .B(PermutationOutput3[1]), 
        .ZN(Red_SignaltoCheck[319]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_79_LFInst_3_U3  ( .A(PermutationOutput3[2]), 
        .B(PermutationOutput3[0]), .ZN(\Red_ToCheckInst_LFInst_79_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_80_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_80_LFInst_0_n2 ), .B(PermutationOutput2[62]), 
        .ZN(Red_SignaltoCheck[320]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_80_LFInst_0_U3  ( .A(PermutationOutput2[63]), .B(PermutationOutput2[61]), .ZN(\Red_ToCheckInst_LFInst_80_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_80_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_80_LFInst_1_n2 ), .B(PermutationOutput2[62]), 
        .ZN(Red_SignaltoCheck[321]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_80_LFInst_1_U3  ( .A(PermutationOutput2[63]), .B(PermutationOutput2[60]), .ZN(\Red_ToCheckInst_LFInst_80_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_80_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_80_LFInst_2_n2 ), .B(PermutationOutput2[61]), 
        .ZN(Red_SignaltoCheck[322]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_80_LFInst_2_U3  ( .A(PermutationOutput2[63]), .B(PermutationOutput2[60]), .ZN(\Red_ToCheckInst_LFInst_80_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_80_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_80_LFInst_3_n2 ), .B(PermutationOutput2[61]), 
        .ZN(Red_SignaltoCheck[323]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_80_LFInst_3_U3  ( .A(PermutationOutput2[62]), .B(PermutationOutput2[60]), .ZN(\Red_ToCheckInst_LFInst_80_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_81_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_81_LFInst_0_n2 ), .B(PermutationOutput2[50]), 
        .ZN(Red_SignaltoCheck[324]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_81_LFInst_0_U3  ( .A(PermutationOutput2[51]), .B(PermutationOutput2[49]), .ZN(\Red_ToCheckInst_LFInst_81_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_81_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_81_LFInst_1_n2 ), .B(PermutationOutput2[50]), 
        .ZN(Red_SignaltoCheck[325]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_81_LFInst_1_U3  ( .A(PermutationOutput2[51]), .B(PermutationOutput2[48]), .ZN(\Red_ToCheckInst_LFInst_81_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_81_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_81_LFInst_2_n2 ), .B(PermutationOutput2[49]), 
        .ZN(Red_SignaltoCheck[326]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_81_LFInst_2_U3  ( .A(PermutationOutput2[51]), .B(PermutationOutput2[48]), .ZN(\Red_ToCheckInst_LFInst_81_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_81_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_81_LFInst_3_n2 ), .B(PermutationOutput2[49]), 
        .ZN(Red_SignaltoCheck[327]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_81_LFInst_3_U3  ( .A(PermutationOutput2[50]), .B(PermutationOutput2[48]), .ZN(\Red_ToCheckInst_LFInst_81_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_82_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_82_LFInst_0_n2 ), .B(PermutationOutput2[54]), 
        .ZN(Red_SignaltoCheck[328]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_82_LFInst_0_U3  ( .A(PermutationOutput2[55]), .B(PermutationOutput2[53]), .ZN(\Red_ToCheckInst_LFInst_82_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_82_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_82_LFInst_1_n2 ), .B(PermutationOutput2[54]), 
        .ZN(Red_SignaltoCheck[329]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_82_LFInst_1_U3  ( .A(PermutationOutput2[55]), .B(PermutationOutput2[52]), .ZN(\Red_ToCheckInst_LFInst_82_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_82_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_82_LFInst_2_n2 ), .B(PermutationOutput2[53]), 
        .ZN(Red_SignaltoCheck[330]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_82_LFInst_2_U3  ( .A(PermutationOutput2[55]), .B(PermutationOutput2[52]), .ZN(\Red_ToCheckInst_LFInst_82_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_82_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_82_LFInst_3_n2 ), .B(PermutationOutput2[53]), 
        .ZN(Red_SignaltoCheck[331]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_82_LFInst_3_U3  ( .A(PermutationOutput2[54]), .B(PermutationOutput2[52]), .ZN(\Red_ToCheckInst_LFInst_82_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_83_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_83_LFInst_0_n2 ), .B(PermutationOutput2[58]), 
        .ZN(Red_SignaltoCheck[332]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_83_LFInst_0_U3  ( .A(PermutationOutput2[59]), .B(PermutationOutput2[57]), .ZN(\Red_ToCheckInst_LFInst_83_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_83_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_83_LFInst_1_n2 ), .B(PermutationOutput2[58]), 
        .ZN(Red_SignaltoCheck[333]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_83_LFInst_1_U3  ( .A(PermutationOutput2[59]), .B(PermutationOutput2[56]), .ZN(\Red_ToCheckInst_LFInst_83_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_83_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_83_LFInst_2_n2 ), .B(PermutationOutput2[57]), 
        .ZN(Red_SignaltoCheck[334]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_83_LFInst_2_U3  ( .A(PermutationOutput2[59]), .B(PermutationOutput2[56]), .ZN(\Red_ToCheckInst_LFInst_83_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_83_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_83_LFInst_3_n2 ), .B(PermutationOutput2[57]), 
        .ZN(Red_SignaltoCheck[335]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_83_LFInst_3_U3  ( .A(PermutationOutput2[58]), .B(PermutationOutput2[56]), .ZN(\Red_ToCheckInst_LFInst_83_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_84_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_84_LFInst_0_n2 ), .B(PermutationOutput2[34]), 
        .ZN(Red_SignaltoCheck[336]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_84_LFInst_0_U3  ( .A(PermutationOutput2[35]), .B(PermutationOutput2[33]), .ZN(\Red_ToCheckInst_LFInst_84_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_84_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_84_LFInst_1_n2 ), .B(PermutationOutput2[34]), 
        .ZN(Red_SignaltoCheck[337]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_84_LFInst_1_U3  ( .A(PermutationOutput2[35]), .B(PermutationOutput2[32]), .ZN(\Red_ToCheckInst_LFInst_84_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_84_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_84_LFInst_2_n2 ), .B(PermutationOutput2[33]), 
        .ZN(Red_SignaltoCheck[338]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_84_LFInst_2_U3  ( .A(PermutationOutput2[35]), .B(PermutationOutput2[32]), .ZN(\Red_ToCheckInst_LFInst_84_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_84_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_84_LFInst_3_n2 ), .B(PermutationOutput2[33]), 
        .ZN(Red_SignaltoCheck[339]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_84_LFInst_3_U3  ( .A(PermutationOutput2[34]), .B(PermutationOutput2[32]), .ZN(\Red_ToCheckInst_LFInst_84_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_85_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_85_LFInst_0_n2 ), .B(PermutationOutput2[46]), 
        .ZN(Red_SignaltoCheck[340]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_85_LFInst_0_U3  ( .A(PermutationOutput2[47]), .B(PermutationOutput2[45]), .ZN(\Red_ToCheckInst_LFInst_85_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_85_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_85_LFInst_1_n2 ), .B(PermutationOutput2[46]), 
        .ZN(Red_SignaltoCheck[341]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_85_LFInst_1_U3  ( .A(PermutationOutput2[47]), .B(PermutationOutput2[44]), .ZN(\Red_ToCheckInst_LFInst_85_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_85_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_85_LFInst_2_n2 ), .B(PermutationOutput2[45]), 
        .ZN(Red_SignaltoCheck[342]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_85_LFInst_2_U3  ( .A(PermutationOutput2[47]), .B(PermutationOutput2[44]), .ZN(\Red_ToCheckInst_LFInst_85_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_85_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_85_LFInst_3_n2 ), .B(PermutationOutput2[45]), 
        .ZN(Red_SignaltoCheck[343]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_85_LFInst_3_U3  ( .A(PermutationOutput2[46]), .B(PermutationOutput2[44]), .ZN(\Red_ToCheckInst_LFInst_85_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_86_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_86_LFInst_0_n2 ), .B(PermutationOutput2[42]), 
        .ZN(Red_SignaltoCheck[344]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_86_LFInst_0_U3  ( .A(PermutationOutput2[43]), .B(PermutationOutput2[41]), .ZN(\Red_ToCheckInst_LFInst_86_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_86_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_86_LFInst_1_n2 ), .B(PermutationOutput2[42]), 
        .ZN(Red_SignaltoCheck[345]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_86_LFInst_1_U3  ( .A(PermutationOutput2[43]), .B(PermutationOutput2[40]), .ZN(\Red_ToCheckInst_LFInst_86_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_86_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_86_LFInst_2_n2 ), .B(PermutationOutput2[41]), 
        .ZN(Red_SignaltoCheck[346]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_86_LFInst_2_U3  ( .A(PermutationOutput2[43]), .B(PermutationOutput2[40]), .ZN(\Red_ToCheckInst_LFInst_86_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_86_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_86_LFInst_3_n2 ), .B(PermutationOutput2[41]), 
        .ZN(Red_SignaltoCheck[347]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_86_LFInst_3_U3  ( .A(PermutationOutput2[42]), .B(PermutationOutput2[40]), .ZN(\Red_ToCheckInst_LFInst_86_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_87_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_87_LFInst_0_n2 ), .B(PermutationOutput2[38]), 
        .ZN(Red_SignaltoCheck[348]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_87_LFInst_0_U3  ( .A(PermutationOutput2[39]), .B(PermutationOutput2[37]), .ZN(\Red_ToCheckInst_LFInst_87_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_87_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_87_LFInst_1_n2 ), .B(PermutationOutput2[38]), 
        .ZN(Red_SignaltoCheck[349]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_87_LFInst_1_U3  ( .A(PermutationOutput2[39]), .B(PermutationOutput2[36]), .ZN(\Red_ToCheckInst_LFInst_87_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_87_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_87_LFInst_2_n2 ), .B(PermutationOutput2[37]), 
        .ZN(Red_SignaltoCheck[350]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_87_LFInst_2_U3  ( .A(PermutationOutput2[39]), .B(PermutationOutput2[36]), .ZN(\Red_ToCheckInst_LFInst_87_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_87_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_87_LFInst_3_n2 ), .B(PermutationOutput2[37]), 
        .ZN(Red_SignaltoCheck[351]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_87_LFInst_3_U3  ( .A(PermutationOutput2[38]), .B(PermutationOutput2[36]), .ZN(\Red_ToCheckInst_LFInst_87_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_88_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_88_LFInst_0_n2 ), .B(PermutationOutput2[18]), 
        .ZN(Red_SignaltoCheck[352]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_88_LFInst_0_U3  ( .A(PermutationOutput2[19]), .B(PermutationOutput2[17]), .ZN(\Red_ToCheckInst_LFInst_88_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_88_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_88_LFInst_1_n2 ), .B(PermutationOutput2[18]), 
        .ZN(Red_SignaltoCheck[353]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_88_LFInst_1_U3  ( .A(PermutationOutput2[19]), .B(PermutationOutput2[16]), .ZN(\Red_ToCheckInst_LFInst_88_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_88_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_88_LFInst_2_n2 ), .B(PermutationOutput2[17]), 
        .ZN(Red_SignaltoCheck[354]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_88_LFInst_2_U3  ( .A(PermutationOutput2[19]), .B(PermutationOutput2[16]), .ZN(\Red_ToCheckInst_LFInst_88_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_88_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_88_LFInst_3_n2 ), .B(PermutationOutput2[17]), 
        .ZN(Red_SignaltoCheck[355]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_88_LFInst_3_U3  ( .A(PermutationOutput2[18]), .B(PermutationOutput2[16]), .ZN(\Red_ToCheckInst_LFInst_88_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_89_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_89_LFInst_0_n2 ), .B(PermutationOutput2[30]), 
        .ZN(Red_SignaltoCheck[356]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_89_LFInst_0_U3  ( .A(PermutationOutput2[31]), .B(PermutationOutput2[29]), .ZN(\Red_ToCheckInst_LFInst_89_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_89_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_89_LFInst_1_n2 ), .B(PermutationOutput2[30]), 
        .ZN(Red_SignaltoCheck[357]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_89_LFInst_1_U3  ( .A(PermutationOutput2[31]), .B(PermutationOutput2[28]), .ZN(\Red_ToCheckInst_LFInst_89_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_89_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_89_LFInst_2_n2 ), .B(PermutationOutput2[29]), 
        .ZN(Red_SignaltoCheck[358]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_89_LFInst_2_U3  ( .A(PermutationOutput2[31]), .B(PermutationOutput2[28]), .ZN(\Red_ToCheckInst_LFInst_89_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_89_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_89_LFInst_3_n2 ), .B(PermutationOutput2[29]), 
        .ZN(Red_SignaltoCheck[359]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_89_LFInst_3_U3  ( .A(PermutationOutput2[30]), .B(PermutationOutput2[28]), .ZN(\Red_ToCheckInst_LFInst_89_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_90_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_90_LFInst_0_n2 ), .B(PermutationOutput2[26]), 
        .ZN(Red_SignaltoCheck[360]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_90_LFInst_0_U3  ( .A(PermutationOutput2[27]), .B(PermutationOutput2[25]), .ZN(\Red_ToCheckInst_LFInst_90_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_90_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_90_LFInst_1_n2 ), .B(PermutationOutput2[26]), 
        .ZN(Red_SignaltoCheck[361]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_90_LFInst_1_U3  ( .A(PermutationOutput2[27]), .B(PermutationOutput2[24]), .ZN(\Red_ToCheckInst_LFInst_90_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_90_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_90_LFInst_2_n2 ), .B(PermutationOutput2[25]), 
        .ZN(Red_SignaltoCheck[362]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_90_LFInst_2_U3  ( .A(PermutationOutput2[27]), .B(PermutationOutput2[24]), .ZN(\Red_ToCheckInst_LFInst_90_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_90_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_90_LFInst_3_n2 ), .B(PermutationOutput2[25]), 
        .ZN(Red_SignaltoCheck[363]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_90_LFInst_3_U3  ( .A(PermutationOutput2[26]), .B(PermutationOutput2[24]), .ZN(\Red_ToCheckInst_LFInst_90_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_91_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_91_LFInst_0_n2 ), .B(PermutationOutput2[22]), 
        .ZN(Red_SignaltoCheck[364]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_91_LFInst_0_U3  ( .A(PermutationOutput2[23]), .B(PermutationOutput2[21]), .ZN(\Red_ToCheckInst_LFInst_91_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_91_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_91_LFInst_1_n2 ), .B(PermutationOutput2[22]), 
        .ZN(Red_SignaltoCheck[365]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_91_LFInst_1_U3  ( .A(PermutationOutput2[23]), .B(PermutationOutput2[20]), .ZN(\Red_ToCheckInst_LFInst_91_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_91_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_91_LFInst_2_n2 ), .B(PermutationOutput2[21]), 
        .ZN(Red_SignaltoCheck[366]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_91_LFInst_2_U3  ( .A(PermutationOutput2[23]), .B(PermutationOutput2[20]), .ZN(\Red_ToCheckInst_LFInst_91_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_91_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_91_LFInst_3_n2 ), .B(PermutationOutput2[21]), 
        .ZN(Red_SignaltoCheck[367]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_91_LFInst_3_U3  ( .A(PermutationOutput2[22]), .B(PermutationOutput2[20]), .ZN(\Red_ToCheckInst_LFInst_91_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_92_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_92_LFInst_0_n2 ), .B(PermutationOutput2[6]), 
        .ZN(Red_SignaltoCheck[368]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_92_LFInst_0_U3  ( .A(PermutationOutput2[7]), 
        .B(PermutationOutput2[5]), .ZN(\Red_ToCheckInst_LFInst_92_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_92_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_92_LFInst_1_n2 ), .B(PermutationOutput2[6]), 
        .ZN(Red_SignaltoCheck[369]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_92_LFInst_1_U3  ( .A(PermutationOutput2[7]), 
        .B(PermutationOutput2[4]), .ZN(\Red_ToCheckInst_LFInst_92_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_92_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_92_LFInst_2_n2 ), .B(PermutationOutput2[5]), 
        .ZN(Red_SignaltoCheck[370]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_92_LFInst_2_U3  ( .A(PermutationOutput2[7]), 
        .B(PermutationOutput2[4]), .ZN(\Red_ToCheckInst_LFInst_92_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_92_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_92_LFInst_3_n2 ), .B(PermutationOutput2[5]), 
        .ZN(Red_SignaltoCheck[371]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_92_LFInst_3_U3  ( .A(PermutationOutput2[6]), 
        .B(PermutationOutput2[4]), .ZN(\Red_ToCheckInst_LFInst_92_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_93_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_93_LFInst_0_n2 ), .B(PermutationOutput2[10]), 
        .ZN(Red_SignaltoCheck[372]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_93_LFInst_0_U3  ( .A(PermutationOutput2[11]), .B(PermutationOutput2[9]), .ZN(\Red_ToCheckInst_LFInst_93_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_93_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_93_LFInst_1_n2 ), .B(PermutationOutput2[10]), 
        .ZN(Red_SignaltoCheck[373]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_93_LFInst_1_U3  ( .A(PermutationOutput2[11]), .B(PermutationOutput2[8]), .ZN(\Red_ToCheckInst_LFInst_93_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_93_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_93_LFInst_2_n2 ), .B(PermutationOutput2[9]), 
        .ZN(Red_SignaltoCheck[374]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_93_LFInst_2_U3  ( .A(PermutationOutput2[11]), .B(PermutationOutput2[8]), .ZN(\Red_ToCheckInst_LFInst_93_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_93_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_93_LFInst_3_n2 ), .B(PermutationOutput2[9]), 
        .ZN(Red_SignaltoCheck[375]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_93_LFInst_3_U3  ( .A(PermutationOutput2[10]), .B(PermutationOutput2[8]), .ZN(\Red_ToCheckInst_LFInst_93_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_94_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_94_LFInst_0_n2 ), .B(PermutationOutput2[14]), 
        .ZN(Red_SignaltoCheck[376]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_94_LFInst_0_U3  ( .A(PermutationOutput2[15]), .B(PermutationOutput2[13]), .ZN(\Red_ToCheckInst_LFInst_94_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_94_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_94_LFInst_1_n2 ), .B(PermutationOutput2[14]), 
        .ZN(Red_SignaltoCheck[377]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_94_LFInst_1_U3  ( .A(PermutationOutput2[15]), .B(PermutationOutput2[12]), .ZN(\Red_ToCheckInst_LFInst_94_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_94_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_94_LFInst_2_n2 ), .B(PermutationOutput2[13]), 
        .ZN(Red_SignaltoCheck[378]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_94_LFInst_2_U3  ( .A(PermutationOutput2[15]), .B(PermutationOutput2[12]), .ZN(\Red_ToCheckInst_LFInst_94_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_94_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_94_LFInst_3_n2 ), .B(PermutationOutput2[13]), 
        .ZN(Red_SignaltoCheck[379]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_94_LFInst_3_U3  ( .A(PermutationOutput2[14]), .B(PermutationOutput2[12]), .ZN(\Red_ToCheckInst_LFInst_94_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_95_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_95_LFInst_0_n2 ), .B(PermutationOutput2[2]), 
        .ZN(Red_SignaltoCheck[380]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_95_LFInst_0_U3  ( .A(PermutationOutput2[3]), 
        .B(PermutationOutput2[1]), .ZN(\Red_ToCheckInst_LFInst_95_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_95_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_95_LFInst_1_n2 ), .B(PermutationOutput2[2]), 
        .ZN(Red_SignaltoCheck[381]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_95_LFInst_1_U3  ( .A(PermutationOutput2[3]), 
        .B(PermutationOutput2[0]), .ZN(\Red_ToCheckInst_LFInst_95_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_95_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_95_LFInst_2_n2 ), .B(PermutationOutput2[1]), 
        .ZN(Red_SignaltoCheck[382]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_95_LFInst_2_U3  ( .A(PermutationOutput2[3]), 
        .B(PermutationOutput2[0]), .ZN(\Red_ToCheckInst_LFInst_95_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_95_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_95_LFInst_3_n2 ), .B(PermutationOutput2[1]), 
        .ZN(Red_SignaltoCheck[383]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_95_LFInst_3_U3  ( .A(PermutationOutput2[2]), 
        .B(PermutationOutput2[0]), .ZN(\Red_ToCheckInst_LFInst_95_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_96_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_96_LFInst_0_n2 ), .B(PermutationOutput[62]), 
        .ZN(Red_SignaltoCheck[384]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_96_LFInst_0_U3  ( .A(PermutationOutput[63]), 
        .B(PermutationOutput[61]), .ZN(\Red_ToCheckInst_LFInst_96_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_96_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_96_LFInst_1_n2 ), .B(PermutationOutput[62]), 
        .ZN(Red_SignaltoCheck[385]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_96_LFInst_1_U3  ( .A(PermutationOutput[63]), 
        .B(PermutationOutput[60]), .ZN(\Red_ToCheckInst_LFInst_96_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_96_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_96_LFInst_2_n2 ), .B(PermutationOutput[61]), 
        .ZN(Red_SignaltoCheck[386]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_96_LFInst_2_U3  ( .A(PermutationOutput[63]), 
        .B(PermutationOutput[60]), .ZN(\Red_ToCheckInst_LFInst_96_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_96_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_96_LFInst_3_n2 ), .B(PermutationOutput[61]), 
        .ZN(Red_SignaltoCheck[387]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_96_LFInst_3_U3  ( .A(PermutationOutput[62]), 
        .B(PermutationOutput[60]), .ZN(\Red_ToCheckInst_LFInst_96_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_97_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_97_LFInst_0_n2 ), .B(PermutationOutput[50]), 
        .ZN(Red_SignaltoCheck[388]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_97_LFInst_0_U3  ( .A(PermutationOutput[51]), 
        .B(PermutationOutput[49]), .ZN(\Red_ToCheckInst_LFInst_97_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_97_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_97_LFInst_1_n2 ), .B(PermutationOutput[50]), 
        .ZN(Red_SignaltoCheck[389]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_97_LFInst_1_U3  ( .A(PermutationOutput[51]), 
        .B(PermutationOutput[48]), .ZN(\Red_ToCheckInst_LFInst_97_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_97_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_97_LFInst_2_n2 ), .B(PermutationOutput[49]), 
        .ZN(Red_SignaltoCheck[390]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_97_LFInst_2_U3  ( .A(PermutationOutput[51]), 
        .B(PermutationOutput[48]), .ZN(\Red_ToCheckInst_LFInst_97_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_97_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_97_LFInst_3_n2 ), .B(PermutationOutput[49]), 
        .ZN(Red_SignaltoCheck[391]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_97_LFInst_3_U3  ( .A(PermutationOutput[50]), 
        .B(PermutationOutput[48]), .ZN(\Red_ToCheckInst_LFInst_97_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_98_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_98_LFInst_0_n2 ), .B(PermutationOutput[54]), 
        .ZN(Red_SignaltoCheck[392]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_98_LFInst_0_U3  ( .A(PermutationOutput[55]), 
        .B(PermutationOutput[53]), .ZN(\Red_ToCheckInst_LFInst_98_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_98_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_98_LFInst_1_n2 ), .B(PermutationOutput[54]), 
        .ZN(Red_SignaltoCheck[393]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_98_LFInst_1_U3  ( .A(PermutationOutput[55]), 
        .B(PermutationOutput[52]), .ZN(\Red_ToCheckInst_LFInst_98_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_98_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_98_LFInst_2_n2 ), .B(PermutationOutput[53]), 
        .ZN(Red_SignaltoCheck[394]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_98_LFInst_2_U3  ( .A(PermutationOutput[55]), 
        .B(PermutationOutput[52]), .ZN(\Red_ToCheckInst_LFInst_98_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_98_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_98_LFInst_3_n2 ), .B(PermutationOutput[53]), 
        .ZN(Red_SignaltoCheck[395]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_98_LFInst_3_U3  ( .A(PermutationOutput[54]), 
        .B(PermutationOutput[52]), .ZN(\Red_ToCheckInst_LFInst_98_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_99_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_99_LFInst_0_n2 ), .B(PermutationOutput[58]), 
        .ZN(Red_SignaltoCheck[396]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_99_LFInst_0_U3  ( .A(PermutationOutput[59]), 
        .B(PermutationOutput[57]), .ZN(\Red_ToCheckInst_LFInst_99_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_99_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_99_LFInst_1_n2 ), .B(PermutationOutput[58]), 
        .ZN(Red_SignaltoCheck[397]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_99_LFInst_1_U3  ( .A(PermutationOutput[59]), 
        .B(PermutationOutput[56]), .ZN(\Red_ToCheckInst_LFInst_99_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_99_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_99_LFInst_2_n2 ), .B(PermutationOutput[57]), 
        .ZN(Red_SignaltoCheck[398]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_99_LFInst_2_U3  ( .A(PermutationOutput[59]), 
        .B(PermutationOutput[56]), .ZN(\Red_ToCheckInst_LFInst_99_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_99_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_99_LFInst_3_n2 ), .B(PermutationOutput[57]), 
        .ZN(Red_SignaltoCheck[399]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_99_LFInst_3_U3  ( .A(PermutationOutput[58]), 
        .B(PermutationOutput[56]), .ZN(\Red_ToCheckInst_LFInst_99_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_100_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_100_LFInst_0_n2 ), .B(PermutationOutput[34]), 
        .ZN(Red_SignaltoCheck[400]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_100_LFInst_0_U3  ( .A(PermutationOutput[35]), .B(PermutationOutput[33]), .ZN(\Red_ToCheckInst_LFInst_100_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_100_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_100_LFInst_1_n2 ), .B(PermutationOutput[34]), 
        .ZN(Red_SignaltoCheck[401]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_100_LFInst_1_U3  ( .A(PermutationOutput[35]), .B(PermutationOutput[32]), .ZN(\Red_ToCheckInst_LFInst_100_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_100_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_100_LFInst_2_n2 ), .B(PermutationOutput[33]), 
        .ZN(Red_SignaltoCheck[402]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_100_LFInst_2_U3  ( .A(PermutationOutput[35]), .B(PermutationOutput[32]), .ZN(\Red_ToCheckInst_LFInst_100_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_100_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_100_LFInst_3_n2 ), .B(PermutationOutput[33]), 
        .ZN(Red_SignaltoCheck[403]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_100_LFInst_3_U3  ( .A(PermutationOutput[34]), .B(PermutationOutput[32]), .ZN(\Red_ToCheckInst_LFInst_100_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_101_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_101_LFInst_0_n2 ), .B(PermutationOutput[46]), 
        .ZN(Red_SignaltoCheck[404]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_101_LFInst_0_U3  ( .A(PermutationOutput[47]), .B(PermutationOutput[45]), .ZN(\Red_ToCheckInst_LFInst_101_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_101_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_101_LFInst_1_n2 ), .B(PermutationOutput[46]), 
        .ZN(Red_SignaltoCheck[405]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_101_LFInst_1_U3  ( .A(PermutationOutput[47]), .B(PermutationOutput[44]), .ZN(\Red_ToCheckInst_LFInst_101_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_101_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_101_LFInst_2_n2 ), .B(PermutationOutput[45]), 
        .ZN(Red_SignaltoCheck[406]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_101_LFInst_2_U3  ( .A(PermutationOutput[47]), .B(PermutationOutput[44]), .ZN(\Red_ToCheckInst_LFInst_101_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_101_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_101_LFInst_3_n2 ), .B(PermutationOutput[45]), 
        .ZN(Red_SignaltoCheck[407]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_101_LFInst_3_U3  ( .A(PermutationOutput[46]), .B(PermutationOutput[44]), .ZN(\Red_ToCheckInst_LFInst_101_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_102_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_102_LFInst_0_n2 ), .B(PermutationOutput[42]), 
        .ZN(Red_SignaltoCheck[408]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_102_LFInst_0_U3  ( .A(PermutationOutput[43]), .B(PermutationOutput[41]), .ZN(\Red_ToCheckInst_LFInst_102_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_102_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_102_LFInst_1_n2 ), .B(PermutationOutput[42]), 
        .ZN(Red_SignaltoCheck[409]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_102_LFInst_1_U3  ( .A(PermutationOutput[43]), .B(PermutationOutput[40]), .ZN(\Red_ToCheckInst_LFInst_102_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_102_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_102_LFInst_2_n2 ), .B(PermutationOutput[41]), 
        .ZN(Red_SignaltoCheck[410]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_102_LFInst_2_U3  ( .A(PermutationOutput[43]), .B(PermutationOutput[40]), .ZN(\Red_ToCheckInst_LFInst_102_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_102_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_102_LFInst_3_n2 ), .B(PermutationOutput[41]), 
        .ZN(Red_SignaltoCheck[411]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_102_LFInst_3_U3  ( .A(PermutationOutput[42]), .B(PermutationOutput[40]), .ZN(\Red_ToCheckInst_LFInst_102_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_103_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_103_LFInst_0_n2 ), .B(PermutationOutput[38]), 
        .ZN(Red_SignaltoCheck[412]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_103_LFInst_0_U3  ( .A(PermutationOutput[39]), .B(PermutationOutput[37]), .ZN(\Red_ToCheckInst_LFInst_103_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_103_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_103_LFInst_1_n2 ), .B(PermutationOutput[38]), 
        .ZN(Red_SignaltoCheck[413]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_103_LFInst_1_U3  ( .A(PermutationOutput[39]), .B(PermutationOutput[36]), .ZN(\Red_ToCheckInst_LFInst_103_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_103_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_103_LFInst_2_n2 ), .B(PermutationOutput[37]), 
        .ZN(Red_SignaltoCheck[414]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_103_LFInst_2_U3  ( .A(PermutationOutput[39]), .B(PermutationOutput[36]), .ZN(\Red_ToCheckInst_LFInst_103_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_103_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_103_LFInst_3_n2 ), .B(PermutationOutput[37]), 
        .ZN(Red_SignaltoCheck[415]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_103_LFInst_3_U3  ( .A(PermutationOutput[38]), .B(PermutationOutput[36]), .ZN(\Red_ToCheckInst_LFInst_103_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_104_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_104_LFInst_0_n2 ), .B(PermutationOutput[18]), 
        .ZN(Red_SignaltoCheck[416]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_104_LFInst_0_U3  ( .A(PermutationOutput[19]), .B(PermutationOutput[17]), .ZN(\Red_ToCheckInst_LFInst_104_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_104_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_104_LFInst_1_n2 ), .B(PermutationOutput[18]), 
        .ZN(Red_SignaltoCheck[417]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_104_LFInst_1_U3  ( .A(PermutationOutput[19]), .B(PermutationOutput[16]), .ZN(\Red_ToCheckInst_LFInst_104_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_104_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_104_LFInst_2_n2 ), .B(PermutationOutput[17]), 
        .ZN(Red_SignaltoCheck[418]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_104_LFInst_2_U3  ( .A(PermutationOutput[19]), .B(PermutationOutput[16]), .ZN(\Red_ToCheckInst_LFInst_104_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_104_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_104_LFInst_3_n2 ), .B(PermutationOutput[17]), 
        .ZN(Red_SignaltoCheck[419]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_104_LFInst_3_U3  ( .A(PermutationOutput[18]), .B(PermutationOutput[16]), .ZN(\Red_ToCheckInst_LFInst_104_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_105_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_105_LFInst_0_n2 ), .B(PermutationOutput[30]), 
        .ZN(Red_SignaltoCheck[420]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_105_LFInst_0_U3  ( .A(PermutationOutput[31]), .B(PermutationOutput[29]), .ZN(\Red_ToCheckInst_LFInst_105_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_105_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_105_LFInst_1_n2 ), .B(PermutationOutput[30]), 
        .ZN(Red_SignaltoCheck[421]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_105_LFInst_1_U3  ( .A(PermutationOutput[31]), .B(PermutationOutput[28]), .ZN(\Red_ToCheckInst_LFInst_105_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_105_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_105_LFInst_2_n2 ), .B(PermutationOutput[29]), 
        .ZN(Red_SignaltoCheck[422]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_105_LFInst_2_U3  ( .A(PermutationOutput[31]), .B(PermutationOutput[28]), .ZN(\Red_ToCheckInst_LFInst_105_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_105_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_105_LFInst_3_n2 ), .B(PermutationOutput[29]), 
        .ZN(Red_SignaltoCheck[423]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_105_LFInst_3_U3  ( .A(PermutationOutput[30]), .B(PermutationOutput[28]), .ZN(\Red_ToCheckInst_LFInst_105_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_106_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_106_LFInst_0_n2 ), .B(PermutationOutput[26]), 
        .ZN(Red_SignaltoCheck[424]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_106_LFInst_0_U3  ( .A(PermutationOutput[27]), .B(PermutationOutput[25]), .ZN(\Red_ToCheckInst_LFInst_106_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_106_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_106_LFInst_1_n2 ), .B(PermutationOutput[26]), 
        .ZN(Red_SignaltoCheck[425]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_106_LFInst_1_U3  ( .A(PermutationOutput[27]), .B(PermutationOutput[24]), .ZN(\Red_ToCheckInst_LFInst_106_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_106_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_106_LFInst_2_n2 ), .B(PermutationOutput[25]), 
        .ZN(Red_SignaltoCheck[426]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_106_LFInst_2_U3  ( .A(PermutationOutput[27]), .B(PermutationOutput[24]), .ZN(\Red_ToCheckInst_LFInst_106_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_106_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_106_LFInst_3_n2 ), .B(PermutationOutput[25]), 
        .ZN(Red_SignaltoCheck[427]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_106_LFInst_3_U3  ( .A(PermutationOutput[26]), .B(PermutationOutput[24]), .ZN(\Red_ToCheckInst_LFInst_106_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_107_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_107_LFInst_0_n2 ), .B(PermutationOutput[22]), 
        .ZN(Red_SignaltoCheck[428]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_107_LFInst_0_U3  ( .A(PermutationOutput[23]), .B(PermutationOutput[21]), .ZN(\Red_ToCheckInst_LFInst_107_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_107_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_107_LFInst_1_n2 ), .B(PermutationOutput[22]), 
        .ZN(Red_SignaltoCheck[429]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_107_LFInst_1_U3  ( .A(PermutationOutput[23]), .B(PermutationOutput[20]), .ZN(\Red_ToCheckInst_LFInst_107_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_107_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_107_LFInst_2_n2 ), .B(PermutationOutput[21]), 
        .ZN(Red_SignaltoCheck[430]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_107_LFInst_2_U3  ( .A(PermutationOutput[23]), .B(PermutationOutput[20]), .ZN(\Red_ToCheckInst_LFInst_107_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_107_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_107_LFInst_3_n2 ), .B(PermutationOutput[21]), 
        .ZN(Red_SignaltoCheck[431]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_107_LFInst_3_U3  ( .A(PermutationOutput[22]), .B(PermutationOutput[20]), .ZN(\Red_ToCheckInst_LFInst_107_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_108_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_108_LFInst_0_n2 ), .B(PermutationOutput[6]), 
        .ZN(Red_SignaltoCheck[432]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_108_LFInst_0_U3  ( .A(PermutationOutput[7]), 
        .B(PermutationOutput[5]), .ZN(\Red_ToCheckInst_LFInst_108_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_108_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_108_LFInst_1_n2 ), .B(PermutationOutput[6]), 
        .ZN(Red_SignaltoCheck[433]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_108_LFInst_1_U3  ( .A(PermutationOutput[7]), 
        .B(PermutationOutput[4]), .ZN(\Red_ToCheckInst_LFInst_108_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_108_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_108_LFInst_2_n2 ), .B(PermutationOutput[5]), 
        .ZN(Red_SignaltoCheck[434]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_108_LFInst_2_U3  ( .A(PermutationOutput[7]), 
        .B(PermutationOutput[4]), .ZN(\Red_ToCheckInst_LFInst_108_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_108_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_108_LFInst_3_n2 ), .B(PermutationOutput[5]), 
        .ZN(Red_SignaltoCheck[435]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_108_LFInst_3_U3  ( .A(PermutationOutput[6]), 
        .B(PermutationOutput[4]), .ZN(\Red_ToCheckInst_LFInst_108_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_109_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_109_LFInst_0_n2 ), .B(PermutationOutput[10]), 
        .ZN(Red_SignaltoCheck[436]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_109_LFInst_0_U3  ( .A(PermutationOutput[11]), .B(PermutationOutput[9]), .ZN(\Red_ToCheckInst_LFInst_109_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_109_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_109_LFInst_1_n2 ), .B(PermutationOutput[10]), 
        .ZN(Red_SignaltoCheck[437]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_109_LFInst_1_U3  ( .A(PermutationOutput[11]), .B(PermutationOutput[8]), .ZN(\Red_ToCheckInst_LFInst_109_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_109_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_109_LFInst_2_n2 ), .B(PermutationOutput[9]), 
        .ZN(Red_SignaltoCheck[438]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_109_LFInst_2_U3  ( .A(PermutationOutput[11]), .B(PermutationOutput[8]), .ZN(\Red_ToCheckInst_LFInst_109_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_109_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_109_LFInst_3_n2 ), .B(PermutationOutput[9]), 
        .ZN(Red_SignaltoCheck[439]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_109_LFInst_3_U3  ( .A(PermutationOutput[10]), .B(PermutationOutput[8]), .ZN(\Red_ToCheckInst_LFInst_109_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_110_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_110_LFInst_0_n2 ), .B(PermutationOutput[14]), 
        .ZN(Red_SignaltoCheck[440]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_110_LFInst_0_U3  ( .A(PermutationOutput[15]), .B(PermutationOutput[13]), .ZN(\Red_ToCheckInst_LFInst_110_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_110_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_110_LFInst_1_n2 ), .B(PermutationOutput[14]), 
        .ZN(Red_SignaltoCheck[441]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_110_LFInst_1_U3  ( .A(PermutationOutput[15]), .B(PermutationOutput[12]), .ZN(\Red_ToCheckInst_LFInst_110_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_110_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_110_LFInst_2_n2 ), .B(PermutationOutput[13]), 
        .ZN(Red_SignaltoCheck[442]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_110_LFInst_2_U3  ( .A(PermutationOutput[15]), .B(PermutationOutput[12]), .ZN(\Red_ToCheckInst_LFInst_110_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_110_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_110_LFInst_3_n2 ), .B(PermutationOutput[13]), 
        .ZN(Red_SignaltoCheck[443]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_110_LFInst_3_U3  ( .A(PermutationOutput[14]), .B(PermutationOutput[12]), .ZN(\Red_ToCheckInst_LFInst_110_LFInst_3_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_111_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_111_LFInst_0_n2 ), .B(PermutationOutput[2]), 
        .ZN(Red_SignaltoCheck[444]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_111_LFInst_0_U3  ( .A(PermutationOutput[3]), 
        .B(PermutationOutput[1]), .ZN(\Red_ToCheckInst_LFInst_111_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_111_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_111_LFInst_1_n2 ), .B(PermutationOutput[2]), 
        .ZN(Red_SignaltoCheck[445]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_111_LFInst_1_U3  ( .A(PermutationOutput[3]), 
        .B(PermutationOutput[0]), .ZN(\Red_ToCheckInst_LFInst_111_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_111_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_111_LFInst_2_n2 ), .B(PermutationOutput[1]), 
        .ZN(Red_SignaltoCheck[446]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_111_LFInst_2_U3  ( .A(PermutationOutput[3]), 
        .B(PermutationOutput[0]), .ZN(\Red_ToCheckInst_LFInst_111_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_111_LFInst_3_U4  ( .A(
        \Red_ToCheckInst_LFInst_111_LFInst_3_n2 ), .B(PermutationOutput[1]), 
        .ZN(Red_SignaltoCheck[447]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_111_LFInst_3_U3  ( .A(PermutationOutput[2]), 
        .B(PermutationOutput[0]), .ZN(\Red_ToCheckInst_LFInst_111_LFInst_3_n2 ) );
  NOR2_X1 \Check1_CheckInst_0_U223  ( .A1(\Check1_CheckInst_0_n222 ), .A2(
        \Check1_CheckInst_0_n221 ), .ZN(Error[0]) );
  NAND2_X1 \Check1_CheckInst_0_U222  ( .A1(\Check1_CheckInst_0_n220 ), .A2(
        \Check1_CheckInst_0_n219 ), .ZN(\Check1_CheckInst_0_n221 ) );
  NOR2_X1 \Check1_CheckInst_0_U221  ( .A1(\Check1_CheckInst_0_n218 ), .A2(
        \Check1_CheckInst_0_n217 ), .ZN(\Check1_CheckInst_0_n219 ) );
  NAND2_X1 \Check1_CheckInst_0_U220  ( .A1(\Check1_CheckInst_0_n216 ), .A2(
        \Check1_CheckInst_0_n215 ), .ZN(\Check1_CheckInst_0_n217 ) );
  NOR2_X1 \Check1_CheckInst_0_U219  ( .A1(\Check1_CheckInst_0_n214 ), .A2(
        \Check1_CheckInst_0_n213 ), .ZN(\Check1_CheckInst_0_n215 ) );
  NAND2_X1 \Check1_CheckInst_0_U218  ( .A1(\Check1_CheckInst_0_n212 ), .A2(
        \Check1_CheckInst_0_n211 ), .ZN(\Check1_CheckInst_0_n213 ) );
  NOR2_X1 \Check1_CheckInst_0_U217  ( .A1(\Check1_CheckInst_0_n210 ), .A2(
        \Check1_CheckInst_0_n209 ), .ZN(\Check1_CheckInst_0_n211 ) );
  NAND2_X1 \Check1_CheckInst_0_U216  ( .A1(\Check1_CheckInst_0_n208 ), .A2(
        \Check1_CheckInst_0_n207 ), .ZN(\Check1_CheckInst_0_n209 ) );
  NOR2_X1 \Check1_CheckInst_0_U215  ( .A1(\Check1_CheckInst_0_n206 ), .A2(
        \Check1_CheckInst_0_n205 ), .ZN(\Check1_CheckInst_0_n207 ) );
  NAND2_X1 \Check1_CheckInst_0_U214  ( .A1(\Check1_CheckInst_0_n204 ), .A2(
        \Check1_CheckInst_0_n203 ), .ZN(\Check1_CheckInst_0_n205 ) );
  XNOR2_X1 \Check1_CheckInst_0_U213  ( .A(Red_Feedback3[36]), .B(
        Red_SignaltoCheck[228]), .ZN(\Check1_CheckInst_0_n203 ) );
  XNOR2_X1 \Check1_CheckInst_0_U212  ( .A(Red_Feedback3[44]), .B(
        Red_SignaltoCheck[236]), .ZN(\Check1_CheckInst_0_n204 ) );
  NAND2_X1 \Check1_CheckInst_0_U211  ( .A1(\Check1_CheckInst_0_n202 ), .A2(
        \Check1_CheckInst_0_n201 ), .ZN(\Check1_CheckInst_0_n206 ) );
  XNOR2_X1 \Check1_CheckInst_0_U210  ( .A(Red_Feedback3[28]), .B(
        Red_SignaltoCheck[220]), .ZN(\Check1_CheckInst_0_n201 ) );
  XNOR2_X1 \Check1_CheckInst_0_U209  ( .A(Red_Feedback3[40]), .B(
        Red_SignaltoCheck[232]), .ZN(\Check1_CheckInst_0_n202 ) );
  NOR2_X1 \Check1_CheckInst_0_U208  ( .A1(\Check1_CheckInst_0_n200 ), .A2(
        \Check1_CheckInst_0_n199 ), .ZN(\Check1_CheckInst_0_n208 ) );
  XOR2_X1 \Check1_CheckInst_0_U207  ( .A(Red_StateRegOutput3[12]), .B(
        Red_SignaltoCheck[268]), .Z(\Check1_CheckInst_0_n199 ) );
  XOR2_X1 \Check1_CheckInst_0_U206  ( .A(Red_Feedback3[32]), .B(
        Red_SignaltoCheck[224]), .Z(\Check1_CheckInst_0_n200 ) );
  NAND2_X1 \Check1_CheckInst_0_U205  ( .A1(\Check1_CheckInst_0_n198 ), .A2(
        \Check1_CheckInst_0_n197 ), .ZN(\Check1_CheckInst_0_n210 ) );
  XNOR2_X1 \Check1_CheckInst_0_U204  ( .A(Red_StateRegOutput3[8]), .B(
        Red_SignaltoCheck[264]), .ZN(\Check1_CheckInst_0_n197 ) );
  XNOR2_X1 \Check1_CheckInst_0_U203  ( .A(Red_StateRegOutput3[16]), .B(
        Red_SignaltoCheck[272]), .ZN(\Check1_CheckInst_0_n198 ) );
  NOR2_X1 \Check1_CheckInst_0_U202  ( .A1(\Check1_CheckInst_0_n196 ), .A2(
        \Check1_CheckInst_0_n195 ), .ZN(\Check1_CheckInst_0_n212 ) );
  NAND2_X1 \Check1_CheckInst_0_U201  ( .A1(\Check1_CheckInst_0_n194 ), .A2(
        \Check1_CheckInst_0_n193 ), .ZN(\Check1_CheckInst_0_n195 ) );
  NOR2_X1 \Check1_CheckInst_0_U200  ( .A1(\Check1_CheckInst_0_n192 ), .A2(
        \Check1_CheckInst_0_n191 ), .ZN(\Check1_CheckInst_0_n193 ) );
  NAND2_X1 \Check1_CheckInst_0_U199  ( .A1(\Check1_CheckInst_0_n190 ), .A2(
        \Check1_CheckInst_0_n189 ), .ZN(\Check1_CheckInst_0_n191 ) );
  XNOR2_X1 \Check1_CheckInst_0_U198  ( .A(Red_StateRegOutput3[4]), .B(
        Red_SignaltoCheck[260]), .ZN(\Check1_CheckInst_0_n189 ) );
  XNOR2_X1 \Check1_CheckInst_0_U197  ( .A(Red_StateRegOutput3[0]), .B(
        Red_SignaltoCheck[256]), .ZN(\Check1_CheckInst_0_n190 ) );
  NAND2_X1 \Check1_CheckInst_0_U196  ( .A1(\Check1_CheckInst_0_n188 ), .A2(
        \Check1_CheckInst_0_n187 ), .ZN(\Check1_CheckInst_0_n192 ) );
  XNOR2_X1 \Check1_CheckInst_0_U195  ( .A(Red_Feedback3[60]), .B(
        Red_SignaltoCheck[252]), .ZN(\Check1_CheckInst_0_n187 ) );
  XNOR2_X1 \Check1_CheckInst_0_U194  ( .A(Red_Feedback3[56]), .B(
        Red_SignaltoCheck[248]), .ZN(\Check1_CheckInst_0_n188 ) );
  NOR2_X1 \Check1_CheckInst_0_U193  ( .A1(\Check1_CheckInst_0_n186 ), .A2(
        \Check1_CheckInst_0_n185 ), .ZN(\Check1_CheckInst_0_n194 ) );
  XOR2_X1 \Check1_CheckInst_0_U192  ( .A(Red_StateRegOutput[28]), .B(
        Red_SignaltoCheck[412]), .Z(\Check1_CheckInst_0_n185 ) );
  XOR2_X1 \Check1_CheckInst_0_U191  ( .A(Red_StateRegOutput[24]), .B(
        Red_SignaltoCheck[408]), .Z(\Check1_CheckInst_0_n186 ) );
  NAND2_X1 \Check1_CheckInst_0_U190  ( .A1(\Check1_CheckInst_0_n184 ), .A2(
        \Check1_CheckInst_0_n183 ), .ZN(\Check1_CheckInst_0_n196 ) );
  XNOR2_X1 \Check1_CheckInst_0_U189  ( .A(Red_StateRegOutput[12]), .B(
        Red_SignaltoCheck[396]), .ZN(\Check1_CheckInst_0_n183 ) );
  XNOR2_X1 \Check1_CheckInst_0_U188  ( .A(Red_StateRegOutput[20]), .B(
        Red_SignaltoCheck[404]), .ZN(\Check1_CheckInst_0_n184 ) );
  NAND2_X1 \Check1_CheckInst_0_U187  ( .A1(\Check1_CheckInst_0_n182 ), .A2(
        \Check1_CheckInst_0_n181 ), .ZN(\Check1_CheckInst_0_n214 ) );
  NOR2_X1 \Check1_CheckInst_0_U186  ( .A1(\Check1_CheckInst_0_n180 ), .A2(
        \Check1_CheckInst_0_n179 ), .ZN(\Check1_CheckInst_0_n181 ) );
  NAND2_X1 \Check1_CheckInst_0_U185  ( .A1(\Check1_CheckInst_0_n178 ), .A2(
        \Check1_CheckInst_0_n177 ), .ZN(\Check1_CheckInst_0_n179 ) );
  NOR2_X1 \Check1_CheckInst_0_U184  ( .A1(\Check1_CheckInst_0_n176 ), .A2(
        \Check1_CheckInst_0_n175 ), .ZN(\Check1_CheckInst_0_n177 ) );
  XOR2_X1 \Check1_CheckInst_0_U183  ( .A(Red_StateRegOutput[4]), .B(
        Red_SignaltoCheck[388]), .Z(\Check1_CheckInst_0_n175 ) );
  XOR2_X1 \Check1_CheckInst_0_U182  ( .A(Red_StateRegOutput[16]), .B(
        Red_SignaltoCheck[400]), .Z(\Check1_CheckInst_0_n176 ) );
  NOR2_X1 \Check1_CheckInst_0_U181  ( .A1(\Check1_CheckInst_0_n174 ), .A2(
        \Check1_CheckInst_0_n173 ), .ZN(\Check1_CheckInst_0_n178 ) );
  XOR2_X1 \Check1_CheckInst_0_U180  ( .A(Red_StateRegOutput[52]), .B(
        Red_SignaltoCheck[436]), .Z(\Check1_CheckInst_0_n173 ) );
  XOR2_X1 \Check1_CheckInst_0_U179  ( .A(Red_StateRegOutput[8]), .B(
        Red_SignaltoCheck[392]), .Z(\Check1_CheckInst_0_n174 ) );
  NAND2_X1 \Check1_CheckInst_0_U178  ( .A1(\Check1_CheckInst_0_n172 ), .A2(
        \Check1_CheckInst_0_n171 ), .ZN(\Check1_CheckInst_0_n180 ) );
  XNOR2_X1 \Check1_CheckInst_0_U177  ( .A(Red_StateRegOutput[48]), .B(
        Red_SignaltoCheck[432]), .ZN(\Check1_CheckInst_0_n171 ) );
  XNOR2_X1 \Check1_CheckInst_0_U176  ( .A(Red_StateRegOutput[56]), .B(
        Red_SignaltoCheck[440]), .ZN(\Check1_CheckInst_0_n172 ) );
  NOR2_X1 \Check1_CheckInst_0_U175  ( .A1(\Check1_CheckInst_0_n170 ), .A2(
        \Check1_CheckInst_0_n169 ), .ZN(\Check1_CheckInst_0_n182 ) );
  XOR2_X1 \Check1_CheckInst_0_U174  ( .A(Red_StateRegOutput[44]), .B(
        Red_SignaltoCheck[428]), .Z(\Check1_CheckInst_0_n169 ) );
  XOR2_X1 \Check1_CheckInst_0_U173  ( .A(Red_StateRegOutput[40]), .B(
        Red_SignaltoCheck[424]), .Z(\Check1_CheckInst_0_n170 ) );
  NOR2_X1 \Check1_CheckInst_0_U172  ( .A1(\Check1_CheckInst_0_n168 ), .A2(
        \Check1_CheckInst_0_n167 ), .ZN(\Check1_CheckInst_0_n216 ) );
  NAND2_X1 \Check1_CheckInst_0_U171  ( .A1(\Check1_CheckInst_0_n166 ), .A2(
        \Check1_CheckInst_0_n165 ), .ZN(\Check1_CheckInst_0_n167 ) );
  NOR2_X1 \Check1_CheckInst_0_U170  ( .A1(\Check1_CheckInst_0_n164 ), .A2(
        \Check1_CheckInst_0_n163 ), .ZN(\Check1_CheckInst_0_n165 ) );
  NAND2_X1 \Check1_CheckInst_0_U169  ( .A1(\Check1_CheckInst_0_n162 ), .A2(
        \Check1_CheckInst_0_n161 ), .ZN(\Check1_CheckInst_0_n163 ) );
  XNOR2_X1 \Check1_CheckInst_0_U168  ( .A(Red_StateRegOutput[36]), .B(
        Red_SignaltoCheck[420]), .ZN(\Check1_CheckInst_0_n161 ) );
  XNOR2_X1 \Check1_CheckInst_0_U167  ( .A(Red_StateRegOutput[32]), .B(
        Red_SignaltoCheck[416]), .ZN(\Check1_CheckInst_0_n162 ) );
  NAND2_X1 \Check1_CheckInst_0_U166  ( .A1(\Check1_CheckInst_0_n160 ), .A2(
        \Check1_CheckInst_0_n159 ), .ZN(\Check1_CheckInst_0_n164 ) );
  XNOR2_X1 \Check1_CheckInst_0_U165  ( .A(Red_StateRegOutput2[36]), .B(
        Red_SignaltoCheck[356]), .ZN(\Check1_CheckInst_0_n159 ) );
  XNOR2_X1 \Check1_CheckInst_0_U164  ( .A(Red_StateRegOutput2[32]), .B(
        Red_SignaltoCheck[352]), .ZN(\Check1_CheckInst_0_n160 ) );
  NOR2_X1 \Check1_CheckInst_0_U163  ( .A1(\Check1_CheckInst_0_n158 ), .A2(
        \Check1_CheckInst_0_n157 ), .ZN(\Check1_CheckInst_0_n166 ) );
  XOR2_X1 \Check1_CheckInst_0_U162  ( .A(Red_StateRegOutput2[20]), .B(
        Red_SignaltoCheck[340]), .Z(\Check1_CheckInst_0_n157 ) );
  XOR2_X1 \Check1_CheckInst_0_U161  ( .A(Red_StateRegOutput2[28]), .B(
        Red_SignaltoCheck[348]), .Z(\Check1_CheckInst_0_n158 ) );
  NAND2_X1 \Check1_CheckInst_0_U160  ( .A1(\Check1_CheckInst_0_n156 ), .A2(
        \Check1_CheckInst_0_n155 ), .ZN(\Check1_CheckInst_0_n168 ) );
  XNOR2_X1 \Check1_CheckInst_0_U159  ( .A(Red_StateRegOutput2[12]), .B(
        Red_SignaltoCheck[332]), .ZN(\Check1_CheckInst_0_n155 ) );
  XNOR2_X1 \Check1_CheckInst_0_U158  ( .A(Red_StateRegOutput2[24]), .B(
        Red_SignaltoCheck[344]), .ZN(\Check1_CheckInst_0_n156 ) );
  NAND2_X1 \Check1_CheckInst_0_U157  ( .A1(\Check1_CheckInst_0_n154 ), .A2(
        \Check1_CheckInst_0_n153 ), .ZN(\Check1_CheckInst_0_n218 ) );
  NOR2_X1 \Check1_CheckInst_0_U156  ( .A1(\Check1_CheckInst_0_n152 ), .A2(
        \Check1_CheckInst_0_n151 ), .ZN(\Check1_CheckInst_0_n153 ) );
  NAND2_X1 \Check1_CheckInst_0_U155  ( .A1(\Check1_CheckInst_0_n150 ), .A2(
        \Check1_CheckInst_0_n149 ), .ZN(\Check1_CheckInst_0_n151 ) );
  NOR2_X1 \Check1_CheckInst_0_U154  ( .A1(\Check1_CheckInst_0_n148 ), .A2(
        \Check1_CheckInst_0_n147 ), .ZN(\Check1_CheckInst_0_n149 ) );
  NAND2_X1 \Check1_CheckInst_0_U153  ( .A1(\Check1_CheckInst_0_n146 ), .A2(
        \Check1_CheckInst_0_n145 ), .ZN(\Check1_CheckInst_0_n147 ) );
  NOR2_X1 \Check1_CheckInst_0_U152  ( .A1(\Check1_CheckInst_0_n144 ), .A2(
        \Check1_CheckInst_0_n143 ), .ZN(\Check1_CheckInst_0_n145 ) );
  NAND2_X1 \Check1_CheckInst_0_U151  ( .A1(\Check1_CheckInst_0_n142 ), .A2(
        \Check1_CheckInst_0_n141 ), .ZN(\Check1_CheckInst_0_n143 ) );
  XNOR2_X1 \Check1_CheckInst_0_U150  ( .A(Red_StateRegOutput2[60]), .B(
        Red_SignaltoCheck[380]), .ZN(\Check1_CheckInst_0_n141 ) );
  XNOR2_X1 \Check1_CheckInst_0_U149  ( .A(Red_StateRegOutput2[16]), .B(
        Red_SignaltoCheck[336]), .ZN(\Check1_CheckInst_0_n142 ) );
  NAND2_X1 \Check1_CheckInst_0_U148  ( .A1(\Check1_CheckInst_0_n140 ), .A2(
        \Check1_CheckInst_0_n139 ), .ZN(\Check1_CheckInst_0_n144 ) );
  XNOR2_X1 \Check1_CheckInst_0_U147  ( .A(Red_StateRegOutput2[56]), .B(
        Red_SignaltoCheck[376]), .ZN(\Check1_CheckInst_0_n139 ) );
  XNOR2_X1 \Check1_CheckInst_0_U146  ( .A(Red_StateRegOutput[0]), .B(
        Red_SignaltoCheck[384]), .ZN(\Check1_CheckInst_0_n140 ) );
  NOR2_X1 \Check1_CheckInst_0_U145  ( .A1(\Check1_CheckInst_0_n138 ), .A2(
        \Check1_CheckInst_0_n137 ), .ZN(\Check1_CheckInst_0_n146 ) );
  XOR2_X1 \Check1_CheckInst_0_U144  ( .A(Red_StateRegOutput2[52]), .B(
        Red_SignaltoCheck[372]), .Z(\Check1_CheckInst_0_n137 ) );
  XOR2_X1 \Check1_CheckInst_0_U143  ( .A(Red_StateRegOutput2[48]), .B(
        Red_SignaltoCheck[368]), .Z(\Check1_CheckInst_0_n138 ) );
  NAND2_X1 \Check1_CheckInst_0_U142  ( .A1(\Check1_CheckInst_0_n136 ), .A2(
        \Check1_CheckInst_0_n135 ), .ZN(\Check1_CheckInst_0_n148 ) );
  XNOR2_X1 \Check1_CheckInst_0_U141  ( .A(Red_StateRegOutput2[44]), .B(
        Red_SignaltoCheck[364]), .ZN(\Check1_CheckInst_0_n135 ) );
  XNOR2_X1 \Check1_CheckInst_0_U140  ( .A(Red_StateRegOutput2[40]), .B(
        Red_SignaltoCheck[360]), .ZN(\Check1_CheckInst_0_n136 ) );
  NOR2_X1 \Check1_CheckInst_0_U139  ( .A1(\Check1_CheckInst_0_n134 ), .A2(
        \Check1_CheckInst_0_n133 ), .ZN(\Check1_CheckInst_0_n150 ) );
  NAND2_X1 \Check1_CheckInst_0_U138  ( .A1(\Check1_CheckInst_0_n132 ), .A2(
        \Check1_CheckInst_0_n131 ), .ZN(\Check1_CheckInst_0_n133 ) );
  NOR2_X1 \Check1_CheckInst_0_U137  ( .A1(\Check1_CheckInst_0_n130 ), .A2(
        \Check1_CheckInst_0_n129 ), .ZN(\Check1_CheckInst_0_n131 ) );
  NAND2_X1 \Check1_CheckInst_0_U136  ( .A1(\Check1_CheckInst_0_n128 ), .A2(
        \Check1_CheckInst_0_n127 ), .ZN(\Check1_CheckInst_0_n129 ) );
  XNOR2_X1 \Check1_CheckInst_0_U135  ( .A(Red_AddRoundKeyOutput2[12]), .B(
        Red_SignaltoCheck[76]), .ZN(\Check1_CheckInst_0_n127 ) );
  XNOR2_X1 \Check1_CheckInst_0_U134  ( .A(Red_AddRoundKeyOutput2[8]), .B(
        Red_SignaltoCheck[72]), .ZN(\Check1_CheckInst_0_n128 ) );
  NAND2_X1 \Check1_CheckInst_0_U133  ( .A1(\Check1_CheckInst_0_n126 ), .A2(
        \Check1_CheckInst_0_n125 ), .ZN(\Check1_CheckInst_0_n130 ) );
  XNOR2_X1 \Check1_CheckInst_0_U132  ( .A(Red_AddRoundKeyOutput3[60]), .B(
        Red_SignaltoCheck[60]), .ZN(\Check1_CheckInst_0_n125 ) );
  XNOR2_X1 \Check1_CheckInst_0_U131  ( .A(Red_AddRoundKeyOutput2[4]), .B(
        Red_SignaltoCheck[68]), .ZN(\Check1_CheckInst_0_n126 ) );
  NOR2_X1 \Check1_CheckInst_0_U130  ( .A1(\Check1_CheckInst_0_n124 ), .A2(
        \Check1_CheckInst_0_n123 ), .ZN(\Check1_CheckInst_0_n132 ) );
  XOR2_X1 \Check1_CheckInst_0_U129  ( .A(Red_AddRoundKeyOutput3[52]), .B(
        Red_SignaltoCheck[52]), .Z(\Check1_CheckInst_0_n123 ) );
  XOR2_X1 \Check1_CheckInst_0_U128  ( .A(Red_AddRoundKeyOutput2[0]), .B(
        Red_SignaltoCheck[64]), .Z(\Check1_CheckInst_0_n124 ) );
  NAND2_X1 \Check1_CheckInst_0_U127  ( .A1(\Check1_CheckInst_0_n122 ), .A2(
        \Check1_CheckInst_0_n121 ), .ZN(\Check1_CheckInst_0_n134 ) );
  XNOR2_X1 \Check1_CheckInst_0_U126  ( .A(Red_AddRoundKeyOutput2[36]), .B(
        Red_SignaltoCheck[100]), .ZN(\Check1_CheckInst_0_n121 ) );
  XNOR2_X1 \Check1_CheckInst_0_U125  ( .A(Red_AddRoundKeyOutput3[56]), .B(
        Red_SignaltoCheck[56]), .ZN(\Check1_CheckInst_0_n122 ) );
  NAND2_X1 \Check1_CheckInst_0_U124  ( .A1(\Check1_CheckInst_0_n120 ), .A2(
        \Check1_CheckInst_0_n119 ), .ZN(\Check1_CheckInst_0_n152 ) );
  NOR2_X1 \Check1_CheckInst_0_U123  ( .A1(\Check1_CheckInst_0_n118 ), .A2(
        \Check1_CheckInst_0_n117 ), .ZN(\Check1_CheckInst_0_n119 ) );
  NAND2_X1 \Check1_CheckInst_0_U122  ( .A1(\Check1_CheckInst_0_n116 ), .A2(
        \Check1_CheckInst_0_n115 ), .ZN(\Check1_CheckInst_0_n117 ) );
  NOR2_X1 \Check1_CheckInst_0_U121  ( .A1(\Check1_CheckInst_0_n114 ), .A2(
        \Check1_CheckInst_0_n113 ), .ZN(\Check1_CheckInst_0_n115 ) );
  XOR2_X1 \Check1_CheckInst_0_U120  ( .A(Red_AddRoundKeyOutput2[32]), .B(
        Red_SignaltoCheck[96]), .Z(\Check1_CheckInst_0_n113 ) );
  XOR2_X1 \Check1_CheckInst_0_U119  ( .A(Red_AddRoundKeyOutput2[40]), .B(
        Red_SignaltoCheck[104]), .Z(\Check1_CheckInst_0_n114 ) );
  NOR2_X1 \Check1_CheckInst_0_U118  ( .A1(\Check1_CheckInst_0_n112 ), .A2(
        \Check1_CheckInst_0_n111 ), .ZN(\Check1_CheckInst_0_n116 ) );
  XOR2_X1 \Check1_CheckInst_0_U117  ( .A(Red_AddRoundKeyOutput2[28]), .B(
        Red_SignaltoCheck[92]), .Z(\Check1_CheckInst_0_n111 ) );
  XOR2_X1 \Check1_CheckInst_0_U116  ( .A(Red_AddRoundKeyOutput2[24]), .B(
        Red_SignaltoCheck[88]), .Z(\Check1_CheckInst_0_n112 ) );
  NAND2_X1 \Check1_CheckInst_0_U115  ( .A1(\Check1_CheckInst_0_n110 ), .A2(
        \Check1_CheckInst_0_n109 ), .ZN(\Check1_CheckInst_0_n118 ) );
  XNOR2_X1 \Check1_CheckInst_0_U114  ( .A(Red_AddRoundKeyOutput2[20]), .B(
        Red_SignaltoCheck[84]), .ZN(\Check1_CheckInst_0_n109 ) );
  XNOR2_X1 \Check1_CheckInst_0_U113  ( .A(Red_AddRoundKeyOutput2[16]), .B(
        Red_SignaltoCheck[80]), .ZN(\Check1_CheckInst_0_n110 ) );
  NOR2_X1 \Check1_CheckInst_0_U112  ( .A1(\Check1_CheckInst_0_n108 ), .A2(
        \Check1_CheckInst_0_n107 ), .ZN(\Check1_CheckInst_0_n120 ) );
  XOR2_X1 \Check1_CheckInst_0_U111  ( .A(Red_AddRoundKeyOutput3[24]), .B(
        Red_SignaltoCheck[24]), .Z(\Check1_CheckInst_0_n107 ) );
  XOR2_X1 \Check1_CheckInst_0_U110  ( .A(Red_AddRoundKeyOutput3[36]), .B(
        Red_SignaltoCheck[36]), .Z(\Check1_CheckInst_0_n108 ) );
  NOR2_X1 \Check1_CheckInst_0_U109  ( .A1(\Check1_CheckInst_0_n106 ), .A2(
        \Check1_CheckInst_0_n105 ), .ZN(\Check1_CheckInst_0_n154 ) );
  NAND2_X1 \Check1_CheckInst_0_U108  ( .A1(\Check1_CheckInst_0_n104 ), .A2(
        \Check1_CheckInst_0_n103 ), .ZN(\Check1_CheckInst_0_n105 ) );
  NOR2_X1 \Check1_CheckInst_0_U107  ( .A1(\Check1_CheckInst_0_n102 ), .A2(
        \Check1_CheckInst_0_n101 ), .ZN(\Check1_CheckInst_0_n103 ) );
  NAND2_X1 \Check1_CheckInst_0_U106  ( .A1(\Check1_CheckInst_0_n100 ), .A2(
        \Check1_CheckInst_0_n99 ), .ZN(\Check1_CheckInst_0_n101 ) );
  XNOR2_X1 \Check1_CheckInst_0_U105  ( .A(Red_AddRoundKeyOutput3[28]), .B(
        Red_SignaltoCheck[28]), .ZN(\Check1_CheckInst_0_n99 ) );
  XNOR2_X1 \Check1_CheckInst_0_U104  ( .A(Red_AddRoundKeyOutput3[32]), .B(
        Red_SignaltoCheck[32]), .ZN(\Check1_CheckInst_0_n100 ) );
  NAND2_X1 \Check1_CheckInst_0_U103  ( .A1(\Check1_CheckInst_0_n98 ), .A2(
        \Check1_CheckInst_0_n97 ), .ZN(\Check1_CheckInst_0_n102 ) );
  XNOR2_X1 \Check1_CheckInst_0_U102  ( .A(Red_AddRoundKeyOutput3[44]), .B(
        Red_SignaltoCheck[44]), .ZN(\Check1_CheckInst_0_n97 ) );
  XNOR2_X1 \Check1_CheckInst_0_U101  ( .A(Red_AddRoundKeyOutput3[40]), .B(
        Red_SignaltoCheck[40]), .ZN(\Check1_CheckInst_0_n98 ) );
  NOR2_X1 \Check1_CheckInst_0_U100  ( .A1(\Check1_CheckInst_0_n96 ), .A2(
        \Check1_CheckInst_0_n95 ), .ZN(\Check1_CheckInst_0_n104 ) );
  XOR2_X1 \Check1_CheckInst_0_U99  ( .A(Red_AddRoundKeyOutput3[8]), .B(
        Red_SignaltoCheck[8]), .Z(\Check1_CheckInst_0_n95 ) );
  XOR2_X1 \Check1_CheckInst_0_U98  ( .A(Red_AddRoundKeyOutput3[48]), .B(
        Red_SignaltoCheck[48]), .Z(\Check1_CheckInst_0_n96 ) );
  NAND2_X1 \Check1_CheckInst_0_U97  ( .A1(\Check1_CheckInst_0_n94 ), .A2(
        \Check1_CheckInst_0_n93 ), .ZN(\Check1_CheckInst_0_n106 ) );
  XNOR2_X1 \Check1_CheckInst_0_U96  ( .A(Red_StateRegOutput[60]), .B(
        Red_SignaltoCheck[444]), .ZN(\Check1_CheckInst_0_n93 ) );
  XNOR2_X1 \Check1_CheckInst_0_U95  ( .A(Red_SignaltoCheck[0]), .B(
        Red_AddRoundKeyOutput3[0]), .ZN(\Check1_CheckInst_0_n94 ) );
  NOR2_X1 \Check1_CheckInst_0_U94  ( .A1(\Check1_CheckInst_0_n92 ), .A2(
        \Check1_CheckInst_0_n91 ), .ZN(\Check1_CheckInst_0_n220 ) );
  NAND2_X1 \Check1_CheckInst_0_U93  ( .A1(\Check1_CheckInst_0_n90 ), .A2(
        \Check1_CheckInst_0_n89 ), .ZN(\Check1_CheckInst_0_n91 ) );
  NOR2_X1 \Check1_CheckInst_0_U92  ( .A1(\Check1_CheckInst_0_n88 ), .A2(
        \Check1_CheckInst_0_n87 ), .ZN(\Check1_CheckInst_0_n89 ) );
  NAND2_X1 \Check1_CheckInst_0_U91  ( .A1(\Check1_CheckInst_0_n86 ), .A2(
        \Check1_CheckInst_0_n85 ), .ZN(\Check1_CheckInst_0_n87 ) );
  NOR2_X1 \Check1_CheckInst_0_U90  ( .A1(\Check1_CheckInst_0_n84 ), .A2(
        \Check1_CheckInst_0_n83 ), .ZN(\Check1_CheckInst_0_n85 ) );
  NAND2_X1 \Check1_CheckInst_0_U89  ( .A1(\Check1_CheckInst_0_n82 ), .A2(
        \Check1_CheckInst_0_n81 ), .ZN(\Check1_CheckInst_0_n83 ) );
  NOR2_X1 \Check1_CheckInst_0_U88  ( .A1(\Check1_CheckInst_0_n80 ), .A2(
        \Check1_CheckInst_0_n79 ), .ZN(\Check1_CheckInst_0_n81 ) );
  XOR2_X1 \Check1_CheckInst_0_U87  ( .A(Red_AddRoundKeyOutput3[12]), .B(
        Red_SignaltoCheck[12]), .Z(\Check1_CheckInst_0_n79 ) );
  XOR2_X1 \Check1_CheckInst_0_U86  ( .A(Red_SignaltoCheck[4]), .B(
        Red_AddRoundKeyOutput3[4]), .Z(\Check1_CheckInst_0_n80 ) );
  NOR2_X1 \Check1_CheckInst_0_U85  ( .A1(\Check1_CheckInst_0_n78 ), .A2(
        \Check1_CheckInst_0_n77 ), .ZN(\Check1_CheckInst_0_n82 ) );
  XOR2_X1 \Check1_CheckInst_0_U84  ( .A(Red_AddRoundKeyOutput3[20]), .B(
        Red_SignaltoCheck[20]), .Z(\Check1_CheckInst_0_n77 ) );
  XOR2_X1 \Check1_CheckInst_0_U83  ( .A(Red_AddRoundKeyOutput3[16]), .B(
        Red_SignaltoCheck[16]), .Z(\Check1_CheckInst_0_n78 ) );
  NAND2_X1 \Check1_CheckInst_0_U82  ( .A1(\Check1_CheckInst_0_n76 ), .A2(
        \Check1_CheckInst_0_n75 ), .ZN(\Check1_CheckInst_0_n84 ) );
  XNOR2_X1 \Check1_CheckInst_0_U81  ( .A(Red_AddRoundKeyOutput[60]), .B(
        Red_SignaltoCheck[188]), .ZN(\Check1_CheckInst_0_n75 ) );
  XNOR2_X1 \Check1_CheckInst_0_U80  ( .A(Red_AddRoundKeyOutput[56]), .B(
        Red_SignaltoCheck[184]), .ZN(\Check1_CheckInst_0_n76 ) );
  NOR2_X1 \Check1_CheckInst_0_U79  ( .A1(\Check1_CheckInst_0_n74 ), .A2(
        \Check1_CheckInst_0_n73 ), .ZN(\Check1_CheckInst_0_n86 ) );
  XOR2_X1 \Check1_CheckInst_0_U78  ( .A(Red_AddRoundKeyOutput[44]), .B(
        Red_SignaltoCheck[172]), .Z(\Check1_CheckInst_0_n73 ) );
  XOR2_X1 \Check1_CheckInst_0_U77  ( .A(Red_AddRoundKeyOutput[52]), .B(
        Red_SignaltoCheck[180]), .Z(\Check1_CheckInst_0_n74 ) );
  NAND2_X1 \Check1_CheckInst_0_U76  ( .A1(\Check1_CheckInst_0_n72 ), .A2(
        \Check1_CheckInst_0_n71 ), .ZN(\Check1_CheckInst_0_n88 ) );
  NOR2_X1 \Check1_CheckInst_0_U75  ( .A1(\Check1_CheckInst_0_n70 ), .A2(
        \Check1_CheckInst_0_n69 ), .ZN(\Check1_CheckInst_0_n71 ) );
  NAND2_X1 \Check1_CheckInst_0_U74  ( .A1(\Check1_CheckInst_0_n68 ), .A2(
        \Check1_CheckInst_0_n67 ), .ZN(\Check1_CheckInst_0_n69 ) );
  NOR2_X1 \Check1_CheckInst_0_U73  ( .A1(\Check1_CheckInst_0_n66 ), .A2(
        \Check1_CheckInst_0_n65 ), .ZN(\Check1_CheckInst_0_n67 ) );
  XOR2_X1 \Check1_CheckInst_0_U72  ( .A(Red_AddRoundKeyOutput[36]), .B(
        Red_SignaltoCheck[164]), .Z(\Check1_CheckInst_0_n65 ) );
  XOR2_X1 \Check1_CheckInst_0_U71  ( .A(Red_AddRoundKeyOutput[48]), .B(
        Red_SignaltoCheck[176]), .Z(\Check1_CheckInst_0_n66 ) );
  NOR2_X1 \Check1_CheckInst_0_U70  ( .A1(\Check1_CheckInst_0_n64 ), .A2(
        \Check1_CheckInst_0_n63 ), .ZN(\Check1_CheckInst_0_n68 ) );
  XOR2_X1 \Check1_CheckInst_0_U69  ( .A(Red_Feedback3[20]), .B(
        Red_SignaltoCheck[212]), .Z(\Check1_CheckInst_0_n63 ) );
  XOR2_X1 \Check1_CheckInst_0_U68  ( .A(Red_AddRoundKeyOutput[40]), .B(
        Red_SignaltoCheck[168]), .Z(\Check1_CheckInst_0_n64 ) );
  NAND2_X1 \Check1_CheckInst_0_U67  ( .A1(\Check1_CheckInst_0_n62 ), .A2(
        \Check1_CheckInst_0_n61 ), .ZN(\Check1_CheckInst_0_n70 ) );
  XNOR2_X1 \Check1_CheckInst_0_U66  ( .A(Red_Feedback3[16]), .B(
        Red_SignaltoCheck[208]), .ZN(\Check1_CheckInst_0_n61 ) );
  XNOR2_X1 \Check1_CheckInst_0_U65  ( .A(Red_Feedback3[24]), .B(
        Red_SignaltoCheck[216]), .ZN(\Check1_CheckInst_0_n62 ) );
  NOR2_X1 \Check1_CheckInst_0_U64  ( .A1(\Check1_CheckInst_0_n60 ), .A2(
        \Check1_CheckInst_0_n59 ), .ZN(\Check1_CheckInst_0_n72 ) );
  XOR2_X1 \Check1_CheckInst_0_U63  ( .A(Red_Feedback3[12]), .B(
        Red_SignaltoCheck[204]), .Z(\Check1_CheckInst_0_n59 ) );
  XOR2_X1 \Check1_CheckInst_0_U62  ( .A(Red_Feedback3[8]), .B(
        Red_SignaltoCheck[200]), .Z(\Check1_CheckInst_0_n60 ) );
  NOR2_X1 \Check1_CheckInst_0_U61  ( .A1(\Check1_CheckInst_0_n58 ), .A2(
        \Check1_CheckInst_0_n57 ), .ZN(\Check1_CheckInst_0_n90 ) );
  NAND2_X1 \Check1_CheckInst_0_U60  ( .A1(\Check1_CheckInst_0_n56 ), .A2(
        \Check1_CheckInst_0_n55 ), .ZN(\Check1_CheckInst_0_n57 ) );
  NOR2_X1 \Check1_CheckInst_0_U59  ( .A1(\Check1_CheckInst_0_n54 ), .A2(
        \Check1_CheckInst_0_n53 ), .ZN(\Check1_CheckInst_0_n55 ) );
  NAND2_X1 \Check1_CheckInst_0_U58  ( .A1(\Check1_CheckInst_0_n52 ), .A2(
        \Check1_CheckInst_0_n51 ), .ZN(\Check1_CheckInst_0_n53 ) );
  XNOR2_X1 \Check1_CheckInst_0_U57  ( .A(Red_Feedback3[4]), .B(
        Red_SignaltoCheck[196]), .ZN(\Check1_CheckInst_0_n51 ) );
  XNOR2_X1 \Check1_CheckInst_0_U56  ( .A(Red_Feedback3[0]), .B(
        Red_SignaltoCheck[192]), .ZN(\Check1_CheckInst_0_n52 ) );
  NAND2_X1 \Check1_CheckInst_0_U55  ( .A1(\Check1_CheckInst_0_n50 ), .A2(
        \Check1_CheckInst_0_n49 ), .ZN(\Check1_CheckInst_0_n54 ) );
  XNOR2_X1 \Check1_CheckInst_0_U54  ( .A(Red_AddRoundKeyOutput[4]), .B(
        Red_SignaltoCheck[132]), .ZN(\Check1_CheckInst_0_n49 ) );
  XNOR2_X1 \Check1_CheckInst_0_U53  ( .A(Red_AddRoundKeyOutput[0]), .B(
        Red_SignaltoCheck[128]), .ZN(\Check1_CheckInst_0_n50 ) );
  NOR2_X1 \Check1_CheckInst_0_U52  ( .A1(\Check1_CheckInst_0_n48 ), .A2(
        \Check1_CheckInst_0_n47 ), .ZN(\Check1_CheckInst_0_n56 ) );
  XOR2_X1 \Check1_CheckInst_0_U51  ( .A(Red_AddRoundKeyOutput2[52]), .B(
        Red_SignaltoCheck[116]), .Z(\Check1_CheckInst_0_n47 ) );
  XOR2_X1 \Check1_CheckInst_0_U50  ( .A(Red_AddRoundKeyOutput2[60]), .B(
        Red_SignaltoCheck[124]), .Z(\Check1_CheckInst_0_n48 ) );
  NAND2_X1 \Check1_CheckInst_0_U49  ( .A1(\Check1_CheckInst_0_n46 ), .A2(
        \Check1_CheckInst_0_n45 ), .ZN(\Check1_CheckInst_0_n58 ) );
  XNOR2_X1 \Check1_CheckInst_0_U48  ( .A(Red_AddRoundKeyOutput2[44]), .B(
        Red_SignaltoCheck[108]), .ZN(\Check1_CheckInst_0_n45 ) );
  XNOR2_X1 \Check1_CheckInst_0_U47  ( .A(Red_AddRoundKeyOutput2[56]), .B(
        Red_SignaltoCheck[120]), .ZN(\Check1_CheckInst_0_n46 ) );
  NAND2_X1 \Check1_CheckInst_0_U46  ( .A1(\Check1_CheckInst_0_n44 ), .A2(
        \Check1_CheckInst_0_n43 ), .ZN(\Check1_CheckInst_0_n92 ) );
  NOR2_X1 \Check1_CheckInst_0_U45  ( .A1(\Check1_CheckInst_0_n42 ), .A2(
        \Check1_CheckInst_0_n41 ), .ZN(\Check1_CheckInst_0_n43 ) );
  NAND2_X1 \Check1_CheckInst_0_U44  ( .A1(\Check1_CheckInst_0_n40 ), .A2(
        \Check1_CheckInst_0_n39 ), .ZN(\Check1_CheckInst_0_n41 ) );
  NOR2_X1 \Check1_CheckInst_0_U43  ( .A1(\Check1_CheckInst_0_n38 ), .A2(
        \Check1_CheckInst_0_n37 ), .ZN(\Check1_CheckInst_0_n39 ) );
  XOR2_X1 \Check1_CheckInst_0_U42  ( .A(Red_AddRoundKeyOutput[28]), .B(
        Red_SignaltoCheck[156]), .Z(\Check1_CheckInst_0_n37 ) );
  XOR2_X1 \Check1_CheckInst_0_U41  ( .A(Red_AddRoundKeyOutput2[48]), .B(
        Red_SignaltoCheck[112]), .Z(\Check1_CheckInst_0_n38 ) );
  NOR2_X1 \Check1_CheckInst_0_U40  ( .A1(\Check1_CheckInst_0_n36 ), .A2(
        \Check1_CheckInst_0_n35 ), .ZN(\Check1_CheckInst_0_n40 ) );
  XOR2_X1 \Check1_CheckInst_0_U39  ( .A(Red_AddRoundKeyOutput[24]), .B(
        Red_SignaltoCheck[152]), .Z(\Check1_CheckInst_0_n35 ) );
  XOR2_X1 \Check1_CheckInst_0_U38  ( .A(Red_AddRoundKeyOutput[32]), .B(
        Red_SignaltoCheck[160]), .Z(\Check1_CheckInst_0_n36 ) );
  NAND2_X1 \Check1_CheckInst_0_U37  ( .A1(\Check1_CheckInst_0_n34 ), .A2(
        \Check1_CheckInst_0_n33 ), .ZN(\Check1_CheckInst_0_n42 ) );
  XNOR2_X1 \Check1_CheckInst_0_U36  ( .A(Red_AddRoundKeyOutput[20]), .B(
        Red_SignaltoCheck[148]), .ZN(\Check1_CheckInst_0_n33 ) );
  XNOR2_X1 \Check1_CheckInst_0_U35  ( .A(Red_AddRoundKeyOutput[16]), .B(
        Red_SignaltoCheck[144]), .ZN(\Check1_CheckInst_0_n34 ) );
  NOR2_X1 \Check1_CheckInst_0_U34  ( .A1(\Check1_CheckInst_0_n32 ), .A2(
        \Check1_CheckInst_0_n31 ), .ZN(\Check1_CheckInst_0_n44 ) );
  XOR2_X1 \Check1_CheckInst_0_U33  ( .A(Red_AddRoundKeyOutput[12]), .B(
        Red_SignaltoCheck[140]), .Z(\Check1_CheckInst_0_n31 ) );
  XOR2_X1 \Check1_CheckInst_0_U32  ( .A(Red_AddRoundKeyOutput[8]), .B(
        Red_SignaltoCheck[136]), .Z(\Check1_CheckInst_0_n32 ) );
  NAND2_X1 \Check1_CheckInst_0_U31  ( .A1(\Check1_CheckInst_0_n30 ), .A2(
        \Check1_CheckInst_0_n29 ), .ZN(\Check1_CheckInst_0_n222 ) );
  NOR2_X1 \Check1_CheckInst_0_U30  ( .A1(\Check1_CheckInst_0_n28 ), .A2(
        \Check1_CheckInst_0_n27 ), .ZN(\Check1_CheckInst_0_n29 ) );
  NAND2_X1 \Check1_CheckInst_0_U29  ( .A1(\Check1_CheckInst_0_n26 ), .A2(
        \Check1_CheckInst_0_n25 ), .ZN(\Check1_CheckInst_0_n27 ) );
  NOR2_X1 \Check1_CheckInst_0_U28  ( .A1(\Check1_CheckInst_0_n24 ), .A2(
        \Check1_CheckInst_0_n23 ), .ZN(\Check1_CheckInst_0_n25 ) );
  NAND2_X1 \Check1_CheckInst_0_U27  ( .A1(\Check1_CheckInst_0_n22 ), .A2(
        \Check1_CheckInst_0_n21 ), .ZN(\Check1_CheckInst_0_n23 ) );
  XNOR2_X1 \Check1_CheckInst_0_U26  ( .A(Red_StateRegOutput3[28]), .B(
        Red_SignaltoCheck[284]), .ZN(\Check1_CheckInst_0_n21 ) );
  XNOR2_X1 \Check1_CheckInst_0_U25  ( .A(Red_StateRegOutput3[36]), .B(
        Red_SignaltoCheck[292]), .ZN(\Check1_CheckInst_0_n22 ) );
  NAND2_X1 \Check1_CheckInst_0_U24  ( .A1(\Check1_CheckInst_0_n20 ), .A2(
        \Check1_CheckInst_0_n19 ), .ZN(\Check1_CheckInst_0_n24 ) );
  XNOR2_X1 \Check1_CheckInst_0_U23  ( .A(Red_StateRegOutput3[44]), .B(
        Red_SignaltoCheck[300]), .ZN(\Check1_CheckInst_0_n19 ) );
  XNOR2_X1 \Check1_CheckInst_0_U22  ( .A(Red_StateRegOutput3[40]), .B(
        Red_SignaltoCheck[296]), .ZN(\Check1_CheckInst_0_n20 ) );
  NOR2_X1 \Check1_CheckInst_0_U21  ( .A1(\Check1_CheckInst_0_n18 ), .A2(
        \Check1_CheckInst_0_n17 ), .ZN(\Check1_CheckInst_0_n26 ) );
  NAND2_X1 \Check1_CheckInst_0_U20  ( .A1(\Check1_CheckInst_0_n16 ), .A2(
        \Check1_CheckInst_0_n15 ), .ZN(\Check1_CheckInst_0_n17 ) );
  XNOR2_X1 \Check1_CheckInst_0_U19  ( .A(Red_StateRegOutput2[4]), .B(
        Red_SignaltoCheck[324]), .ZN(\Check1_CheckInst_0_n15 ) );
  XNOR2_X1 \Check1_CheckInst_0_U18  ( .A(Red_StateRegOutput3[24]), .B(
        Red_SignaltoCheck[280]), .ZN(\Check1_CheckInst_0_n16 ) );
  NAND2_X1 \Check1_CheckInst_0_U17  ( .A1(\Check1_CheckInst_0_n14 ), .A2(
        \Check1_CheckInst_0_n13 ), .ZN(\Check1_CheckInst_0_n18 ) );
  XNOR2_X1 \Check1_CheckInst_0_U16  ( .A(Red_StateRegOutput3[20]), .B(
        Red_SignaltoCheck[276]), .ZN(\Check1_CheckInst_0_n13 ) );
  XNOR2_X1 \Check1_CheckInst_0_U15  ( .A(Red_StateRegOutput3[32]), .B(
        Red_SignaltoCheck[288]), .ZN(\Check1_CheckInst_0_n14 ) );
  NAND2_X1 \Check1_CheckInst_0_U14  ( .A1(\Check1_CheckInst_0_n12 ), .A2(
        \Check1_CheckInst_0_n11 ), .ZN(\Check1_CheckInst_0_n28 ) );
  NOR2_X1 \Check1_CheckInst_0_U13  ( .A1(\Check1_CheckInst_0_n10 ), .A2(
        \Check1_CheckInst_0_n9 ), .ZN(\Check1_CheckInst_0_n11 ) );
  XOR2_X1 \Check1_CheckInst_0_U12  ( .A(Red_StateRegOutput3[60]), .B(
        Red_SignaltoCheck[316]), .Z(\Check1_CheckInst_0_n9 ) );
  XOR2_X1 \Check1_CheckInst_0_U11  ( .A(Red_StateRegOutput3[56]), .B(
        Red_SignaltoCheck[312]), .Z(\Check1_CheckInst_0_n10 ) );
  NOR2_X1 \Check1_CheckInst_0_U10  ( .A1(\Check1_CheckInst_0_n8 ), .A2(
        \Check1_CheckInst_0_n7 ), .ZN(\Check1_CheckInst_0_n12 ) );
  XOR2_X1 \Check1_CheckInst_0_U9  ( .A(Red_StateRegOutput2[0]), .B(
        Red_SignaltoCheck[320]), .Z(\Check1_CheckInst_0_n7 ) );
  XOR2_X1 \Check1_CheckInst_0_U8  ( .A(Red_StateRegOutput2[8]), .B(
        Red_SignaltoCheck[328]), .Z(\Check1_CheckInst_0_n8 ) );
  NOR2_X1 \Check1_CheckInst_0_U7  ( .A1(\Check1_CheckInst_0_n6 ), .A2(
        \Check1_CheckInst_0_n5 ), .ZN(\Check1_CheckInst_0_n30 ) );
  NAND2_X1 \Check1_CheckInst_0_U6  ( .A1(\Check1_CheckInst_0_n4 ), .A2(
        \Check1_CheckInst_0_n3 ), .ZN(\Check1_CheckInst_0_n5 ) );
  XNOR2_X1 \Check1_CheckInst_0_U5  ( .A(Red_Feedback3[52]), .B(
        Red_SignaltoCheck[244]), .ZN(\Check1_CheckInst_0_n3 ) );
  XNOR2_X1 \Check1_CheckInst_0_U4  ( .A(Red_Feedback3[48]), .B(
        Red_SignaltoCheck[240]), .ZN(\Check1_CheckInst_0_n4 ) );
  NAND2_X1 \Check1_CheckInst_0_U3  ( .A1(\Check1_CheckInst_0_n2 ), .A2(
        \Check1_CheckInst_0_n1 ), .ZN(\Check1_CheckInst_0_n6 ) );
  XNOR2_X1 \Check1_CheckInst_0_U2  ( .A(Red_StateRegOutput3[52]), .B(
        Red_SignaltoCheck[308]), .ZN(\Check1_CheckInst_0_n1 ) );
  XNOR2_X1 \Check1_CheckInst_0_U1  ( .A(Red_StateRegOutput3[48]), .B(
        Red_SignaltoCheck[304]), .ZN(\Check1_CheckInst_0_n2 ) );
  NOR2_X1 \Check1_CheckInst_1_U223  ( .A1(\Check1_CheckInst_1_n224 ), .A2(
        \Check1_CheckInst_1_n223 ), .ZN(Error[1]) );
  NAND2_X1 \Check1_CheckInst_1_U222  ( .A1(\Check1_CheckInst_1_n222 ), .A2(
        \Check1_CheckInst_1_n221 ), .ZN(\Check1_CheckInst_1_n223 ) );
  NOR2_X1 \Check1_CheckInst_1_U221  ( .A1(\Check1_CheckInst_1_n220 ), .A2(
        \Check1_CheckInst_1_n219 ), .ZN(\Check1_CheckInst_1_n221 ) );
  NAND2_X1 \Check1_CheckInst_1_U220  ( .A1(\Check1_CheckInst_1_n218 ), .A2(
        \Check1_CheckInst_1_n217 ), .ZN(\Check1_CheckInst_1_n219 ) );
  NOR2_X1 \Check1_CheckInst_1_U219  ( .A1(\Check1_CheckInst_1_n216 ), .A2(
        \Check1_CheckInst_1_n215 ), .ZN(\Check1_CheckInst_1_n217 ) );
  NAND2_X1 \Check1_CheckInst_1_U218  ( .A1(\Check1_CheckInst_1_n214 ), .A2(
        \Check1_CheckInst_1_n213 ), .ZN(\Check1_CheckInst_1_n215 ) );
  NOR2_X1 \Check1_CheckInst_1_U217  ( .A1(\Check1_CheckInst_1_n212 ), .A2(
        \Check1_CheckInst_1_n211 ), .ZN(\Check1_CheckInst_1_n213 ) );
  NAND2_X1 \Check1_CheckInst_1_U216  ( .A1(\Check1_CheckInst_1_n210 ), .A2(
        \Check1_CheckInst_1_n209 ), .ZN(\Check1_CheckInst_1_n211 ) );
  NOR2_X1 \Check1_CheckInst_1_U215  ( .A1(\Check1_CheckInst_1_n208 ), .A2(
        \Check1_CheckInst_1_n207 ), .ZN(\Check1_CheckInst_1_n209 ) );
  NAND2_X1 \Check1_CheckInst_1_U214  ( .A1(\Check1_CheckInst_1_n206 ), .A2(
        \Check1_CheckInst_1_n205 ), .ZN(\Check1_CheckInst_1_n207 ) );
  XNOR2_X1 \Check1_CheckInst_1_U213  ( .A(Red_Feedback3[37]), .B(
        Red_SignaltoCheck[229]), .ZN(\Check1_CheckInst_1_n205 ) );
  XNOR2_X1 \Check1_CheckInst_1_U212  ( .A(Red_Feedback3[45]), .B(
        Red_SignaltoCheck[237]), .ZN(\Check1_CheckInst_1_n206 ) );
  NAND2_X1 \Check1_CheckInst_1_U211  ( .A1(\Check1_CheckInst_1_n204 ), .A2(
        \Check1_CheckInst_1_n203 ), .ZN(\Check1_CheckInst_1_n208 ) );
  XNOR2_X1 \Check1_CheckInst_1_U210  ( .A(Red_Feedback3[29]), .B(
        Red_SignaltoCheck[221]), .ZN(\Check1_CheckInst_1_n203 ) );
  XNOR2_X1 \Check1_CheckInst_1_U209  ( .A(Red_Feedback3[41]), .B(
        Red_SignaltoCheck[233]), .ZN(\Check1_CheckInst_1_n204 ) );
  NOR2_X1 \Check1_CheckInst_1_U208  ( .A1(\Check1_CheckInst_1_n202 ), .A2(
        \Check1_CheckInst_1_n201 ), .ZN(\Check1_CheckInst_1_n210 ) );
  XOR2_X1 \Check1_CheckInst_1_U207  ( .A(Red_StateRegOutput3[13]), .B(
        Red_SignaltoCheck[269]), .Z(\Check1_CheckInst_1_n201 ) );
  XOR2_X1 \Check1_CheckInst_1_U206  ( .A(Red_Feedback3[33]), .B(
        Red_SignaltoCheck[225]), .Z(\Check1_CheckInst_1_n202 ) );
  NAND2_X1 \Check1_CheckInst_1_U205  ( .A1(\Check1_CheckInst_1_n200 ), .A2(
        \Check1_CheckInst_1_n199 ), .ZN(\Check1_CheckInst_1_n212 ) );
  XNOR2_X1 \Check1_CheckInst_1_U204  ( .A(Red_StateRegOutput3[9]), .B(
        Red_SignaltoCheck[265]), .ZN(\Check1_CheckInst_1_n199 ) );
  XNOR2_X1 \Check1_CheckInst_1_U203  ( .A(Red_StateRegOutput3[17]), .B(
        Red_SignaltoCheck[273]), .ZN(\Check1_CheckInst_1_n200 ) );
  NOR2_X1 \Check1_CheckInst_1_U202  ( .A1(\Check1_CheckInst_1_n198 ), .A2(
        \Check1_CheckInst_1_n197 ), .ZN(\Check1_CheckInst_1_n214 ) );
  NAND2_X1 \Check1_CheckInst_1_U201  ( .A1(\Check1_CheckInst_1_n196 ), .A2(
        \Check1_CheckInst_1_n195 ), .ZN(\Check1_CheckInst_1_n197 ) );
  NOR2_X1 \Check1_CheckInst_1_U200  ( .A1(\Check1_CheckInst_1_n194 ), .A2(
        \Check1_CheckInst_1_n193 ), .ZN(\Check1_CheckInst_1_n195 ) );
  NAND2_X1 \Check1_CheckInst_1_U199  ( .A1(\Check1_CheckInst_1_n192 ), .A2(
        \Check1_CheckInst_1_n191 ), .ZN(\Check1_CheckInst_1_n193 ) );
  XNOR2_X1 \Check1_CheckInst_1_U198  ( .A(Red_StateRegOutput3[5]), .B(
        Red_SignaltoCheck[261]), .ZN(\Check1_CheckInst_1_n191 ) );
  XNOR2_X1 \Check1_CheckInst_1_U197  ( .A(Red_StateRegOutput3[1]), .B(
        Red_SignaltoCheck[257]), .ZN(\Check1_CheckInst_1_n192 ) );
  NAND2_X1 \Check1_CheckInst_1_U196  ( .A1(\Check1_CheckInst_1_n190 ), .A2(
        \Check1_CheckInst_1_n189 ), .ZN(\Check1_CheckInst_1_n194 ) );
  XNOR2_X1 \Check1_CheckInst_1_U195  ( .A(Red_Feedback3[61]), .B(
        Red_SignaltoCheck[253]), .ZN(\Check1_CheckInst_1_n189 ) );
  XNOR2_X1 \Check1_CheckInst_1_U194  ( .A(Red_Feedback3[57]), .B(
        Red_SignaltoCheck[249]), .ZN(\Check1_CheckInst_1_n190 ) );
  NOR2_X1 \Check1_CheckInst_1_U193  ( .A1(\Check1_CheckInst_1_n188 ), .A2(
        \Check1_CheckInst_1_n187 ), .ZN(\Check1_CheckInst_1_n196 ) );
  XOR2_X1 \Check1_CheckInst_1_U192  ( .A(Red_StateRegOutput[29]), .B(
        Red_SignaltoCheck[413]), .Z(\Check1_CheckInst_1_n187 ) );
  XOR2_X1 \Check1_CheckInst_1_U191  ( .A(Red_StateRegOutput[25]), .B(
        Red_SignaltoCheck[409]), .Z(\Check1_CheckInst_1_n188 ) );
  NAND2_X1 \Check1_CheckInst_1_U190  ( .A1(\Check1_CheckInst_1_n186 ), .A2(
        \Check1_CheckInst_1_n185 ), .ZN(\Check1_CheckInst_1_n198 ) );
  XNOR2_X1 \Check1_CheckInst_1_U189  ( .A(Red_StateRegOutput[13]), .B(
        Red_SignaltoCheck[397]), .ZN(\Check1_CheckInst_1_n185 ) );
  XNOR2_X1 \Check1_CheckInst_1_U188  ( .A(Red_StateRegOutput[21]), .B(
        Red_SignaltoCheck[405]), .ZN(\Check1_CheckInst_1_n186 ) );
  NAND2_X1 \Check1_CheckInst_1_U187  ( .A1(\Check1_CheckInst_1_n184 ), .A2(
        \Check1_CheckInst_1_n183 ), .ZN(\Check1_CheckInst_1_n216 ) );
  NOR2_X1 \Check1_CheckInst_1_U186  ( .A1(\Check1_CheckInst_1_n182 ), .A2(
        \Check1_CheckInst_1_n181 ), .ZN(\Check1_CheckInst_1_n183 ) );
  NAND2_X1 \Check1_CheckInst_1_U185  ( .A1(\Check1_CheckInst_1_n180 ), .A2(
        \Check1_CheckInst_1_n179 ), .ZN(\Check1_CheckInst_1_n181 ) );
  NOR2_X1 \Check1_CheckInst_1_U184  ( .A1(\Check1_CheckInst_1_n178 ), .A2(
        \Check1_CheckInst_1_n177 ), .ZN(\Check1_CheckInst_1_n179 ) );
  XOR2_X1 \Check1_CheckInst_1_U183  ( .A(Red_StateRegOutput[5]), .B(
        Red_SignaltoCheck[389]), .Z(\Check1_CheckInst_1_n177 ) );
  XOR2_X1 \Check1_CheckInst_1_U182  ( .A(Red_StateRegOutput[17]), .B(
        Red_SignaltoCheck[401]), .Z(\Check1_CheckInst_1_n178 ) );
  NOR2_X1 \Check1_CheckInst_1_U181  ( .A1(\Check1_CheckInst_1_n176 ), .A2(
        \Check1_CheckInst_1_n175 ), .ZN(\Check1_CheckInst_1_n180 ) );
  XOR2_X1 \Check1_CheckInst_1_U180  ( .A(Red_StateRegOutput[53]), .B(
        Red_SignaltoCheck[437]), .Z(\Check1_CheckInst_1_n175 ) );
  XOR2_X1 \Check1_CheckInst_1_U179  ( .A(Red_StateRegOutput[9]), .B(
        Red_SignaltoCheck[393]), .Z(\Check1_CheckInst_1_n176 ) );
  NAND2_X1 \Check1_CheckInst_1_U178  ( .A1(\Check1_CheckInst_1_n174 ), .A2(
        \Check1_CheckInst_1_n173 ), .ZN(\Check1_CheckInst_1_n182 ) );
  XNOR2_X1 \Check1_CheckInst_1_U177  ( .A(Red_StateRegOutput[49]), .B(
        Red_SignaltoCheck[433]), .ZN(\Check1_CheckInst_1_n173 ) );
  XNOR2_X1 \Check1_CheckInst_1_U176  ( .A(Red_StateRegOutput[57]), .B(
        Red_SignaltoCheck[441]), .ZN(\Check1_CheckInst_1_n174 ) );
  NOR2_X1 \Check1_CheckInst_1_U175  ( .A1(\Check1_CheckInst_1_n172 ), .A2(
        \Check1_CheckInst_1_n171 ), .ZN(\Check1_CheckInst_1_n184 ) );
  XOR2_X1 \Check1_CheckInst_1_U174  ( .A(Red_StateRegOutput[45]), .B(
        Red_SignaltoCheck[429]), .Z(\Check1_CheckInst_1_n171 ) );
  XOR2_X1 \Check1_CheckInst_1_U173  ( .A(Red_StateRegOutput[41]), .B(
        Red_SignaltoCheck[425]), .Z(\Check1_CheckInst_1_n172 ) );
  NOR2_X1 \Check1_CheckInst_1_U172  ( .A1(\Check1_CheckInst_1_n170 ), .A2(
        \Check1_CheckInst_1_n169 ), .ZN(\Check1_CheckInst_1_n218 ) );
  NAND2_X1 \Check1_CheckInst_1_U171  ( .A1(\Check1_CheckInst_1_n168 ), .A2(
        \Check1_CheckInst_1_n167 ), .ZN(\Check1_CheckInst_1_n169 ) );
  NOR2_X1 \Check1_CheckInst_1_U170  ( .A1(\Check1_CheckInst_1_n166 ), .A2(
        \Check1_CheckInst_1_n165 ), .ZN(\Check1_CheckInst_1_n167 ) );
  NAND2_X1 \Check1_CheckInst_1_U169  ( .A1(\Check1_CheckInst_1_n164 ), .A2(
        \Check1_CheckInst_1_n163 ), .ZN(\Check1_CheckInst_1_n165 ) );
  XNOR2_X1 \Check1_CheckInst_1_U168  ( .A(Red_StateRegOutput[37]), .B(
        Red_SignaltoCheck[421]), .ZN(\Check1_CheckInst_1_n163 ) );
  XNOR2_X1 \Check1_CheckInst_1_U167  ( .A(Red_StateRegOutput[33]), .B(
        Red_SignaltoCheck[417]), .ZN(\Check1_CheckInst_1_n164 ) );
  NAND2_X1 \Check1_CheckInst_1_U166  ( .A1(\Check1_CheckInst_1_n162 ), .A2(
        \Check1_CheckInst_1_n161 ), .ZN(\Check1_CheckInst_1_n166 ) );
  XNOR2_X1 \Check1_CheckInst_1_U165  ( .A(Red_StateRegOutput2[37]), .B(
        Red_SignaltoCheck[357]), .ZN(\Check1_CheckInst_1_n161 ) );
  XNOR2_X1 \Check1_CheckInst_1_U164  ( .A(Red_StateRegOutput2[33]), .B(
        Red_SignaltoCheck[353]), .ZN(\Check1_CheckInst_1_n162 ) );
  NOR2_X1 \Check1_CheckInst_1_U163  ( .A1(\Check1_CheckInst_1_n160 ), .A2(
        \Check1_CheckInst_1_n159 ), .ZN(\Check1_CheckInst_1_n168 ) );
  XOR2_X1 \Check1_CheckInst_1_U162  ( .A(Red_StateRegOutput2[21]), .B(
        Red_SignaltoCheck[341]), .Z(\Check1_CheckInst_1_n159 ) );
  XOR2_X1 \Check1_CheckInst_1_U161  ( .A(Red_StateRegOutput2[29]), .B(
        Red_SignaltoCheck[349]), .Z(\Check1_CheckInst_1_n160 ) );
  NAND2_X1 \Check1_CheckInst_1_U160  ( .A1(\Check1_CheckInst_1_n158 ), .A2(
        \Check1_CheckInst_1_n157 ), .ZN(\Check1_CheckInst_1_n170 ) );
  XNOR2_X1 \Check1_CheckInst_1_U159  ( .A(Red_StateRegOutput2[13]), .B(
        Red_SignaltoCheck[333]), .ZN(\Check1_CheckInst_1_n157 ) );
  XNOR2_X1 \Check1_CheckInst_1_U158  ( .A(Red_StateRegOutput2[25]), .B(
        Red_SignaltoCheck[345]), .ZN(\Check1_CheckInst_1_n158 ) );
  NAND2_X1 \Check1_CheckInst_1_U157  ( .A1(\Check1_CheckInst_1_n156 ), .A2(
        \Check1_CheckInst_1_n155 ), .ZN(\Check1_CheckInst_1_n220 ) );
  NOR2_X1 \Check1_CheckInst_1_U156  ( .A1(\Check1_CheckInst_1_n154 ), .A2(
        \Check1_CheckInst_1_n153 ), .ZN(\Check1_CheckInst_1_n155 ) );
  NAND2_X1 \Check1_CheckInst_1_U155  ( .A1(\Check1_CheckInst_1_n152 ), .A2(
        \Check1_CheckInst_1_n151 ), .ZN(\Check1_CheckInst_1_n153 ) );
  NOR2_X1 \Check1_CheckInst_1_U154  ( .A1(\Check1_CheckInst_1_n150 ), .A2(
        \Check1_CheckInst_1_n149 ), .ZN(\Check1_CheckInst_1_n151 ) );
  NAND2_X1 \Check1_CheckInst_1_U153  ( .A1(\Check1_CheckInst_1_n148 ), .A2(
        \Check1_CheckInst_1_n147 ), .ZN(\Check1_CheckInst_1_n149 ) );
  NOR2_X1 \Check1_CheckInst_1_U152  ( .A1(\Check1_CheckInst_1_n146 ), .A2(
        \Check1_CheckInst_1_n145 ), .ZN(\Check1_CheckInst_1_n147 ) );
  NAND2_X1 \Check1_CheckInst_1_U151  ( .A1(\Check1_CheckInst_1_n144 ), .A2(
        \Check1_CheckInst_1_n143 ), .ZN(\Check1_CheckInst_1_n145 ) );
  XNOR2_X1 \Check1_CheckInst_1_U150  ( .A(Red_StateRegOutput2[61]), .B(
        Red_SignaltoCheck[381]), .ZN(\Check1_CheckInst_1_n143 ) );
  XNOR2_X1 \Check1_CheckInst_1_U149  ( .A(Red_StateRegOutput2[17]), .B(
        Red_SignaltoCheck[337]), .ZN(\Check1_CheckInst_1_n144 ) );
  NAND2_X1 \Check1_CheckInst_1_U148  ( .A1(\Check1_CheckInst_1_n142 ), .A2(
        \Check1_CheckInst_1_n141 ), .ZN(\Check1_CheckInst_1_n146 ) );
  XNOR2_X1 \Check1_CheckInst_1_U147  ( .A(Red_StateRegOutput2[57]), .B(
        Red_SignaltoCheck[377]), .ZN(\Check1_CheckInst_1_n141 ) );
  XNOR2_X1 \Check1_CheckInst_1_U146  ( .A(Red_StateRegOutput[1]), .B(
        Red_SignaltoCheck[385]), .ZN(\Check1_CheckInst_1_n142 ) );
  NOR2_X1 \Check1_CheckInst_1_U145  ( .A1(\Check1_CheckInst_1_n140 ), .A2(
        \Check1_CheckInst_1_n139 ), .ZN(\Check1_CheckInst_1_n148 ) );
  XOR2_X1 \Check1_CheckInst_1_U144  ( .A(Red_StateRegOutput2[53]), .B(
        Red_SignaltoCheck[373]), .Z(\Check1_CheckInst_1_n139 ) );
  XOR2_X1 \Check1_CheckInst_1_U143  ( .A(Red_StateRegOutput2[49]), .B(
        Red_SignaltoCheck[369]), .Z(\Check1_CheckInst_1_n140 ) );
  NAND2_X1 \Check1_CheckInst_1_U142  ( .A1(\Check1_CheckInst_1_n138 ), .A2(
        \Check1_CheckInst_1_n137 ), .ZN(\Check1_CheckInst_1_n150 ) );
  XNOR2_X1 \Check1_CheckInst_1_U141  ( .A(Red_StateRegOutput2[45]), .B(
        Red_SignaltoCheck[365]), .ZN(\Check1_CheckInst_1_n137 ) );
  XNOR2_X1 \Check1_CheckInst_1_U140  ( .A(Red_StateRegOutput2[41]), .B(
        Red_SignaltoCheck[361]), .ZN(\Check1_CheckInst_1_n138 ) );
  NOR2_X1 \Check1_CheckInst_1_U139  ( .A1(\Check1_CheckInst_1_n136 ), .A2(
        \Check1_CheckInst_1_n135 ), .ZN(\Check1_CheckInst_1_n152 ) );
  NAND2_X1 \Check1_CheckInst_1_U138  ( .A1(\Check1_CheckInst_1_n134 ), .A2(
        \Check1_CheckInst_1_n133 ), .ZN(\Check1_CheckInst_1_n135 ) );
  NOR2_X1 \Check1_CheckInst_1_U137  ( .A1(\Check1_CheckInst_1_n132 ), .A2(
        \Check1_CheckInst_1_n131 ), .ZN(\Check1_CheckInst_1_n133 ) );
  NAND2_X1 \Check1_CheckInst_1_U136  ( .A1(\Check1_CheckInst_1_n130 ), .A2(
        \Check1_CheckInst_1_n129 ), .ZN(\Check1_CheckInst_1_n131 ) );
  XNOR2_X1 \Check1_CheckInst_1_U135  ( .A(Red_AddRoundKeyOutput2[13]), .B(
        Red_SignaltoCheck[77]), .ZN(\Check1_CheckInst_1_n129 ) );
  XNOR2_X1 \Check1_CheckInst_1_U134  ( .A(Red_AddRoundKeyOutput2[9]), .B(
        Red_SignaltoCheck[73]), .ZN(\Check1_CheckInst_1_n130 ) );
  NAND2_X1 \Check1_CheckInst_1_U133  ( .A1(\Check1_CheckInst_1_n128 ), .A2(
        \Check1_CheckInst_1_n127 ), .ZN(\Check1_CheckInst_1_n132 ) );
  XNOR2_X1 \Check1_CheckInst_1_U132  ( .A(Red_AddRoundKeyOutput3[61]), .B(
        Red_SignaltoCheck[61]), .ZN(\Check1_CheckInst_1_n127 ) );
  XNOR2_X1 \Check1_CheckInst_1_U131  ( .A(Red_AddRoundKeyOutput2[5]), .B(
        Red_SignaltoCheck[69]), .ZN(\Check1_CheckInst_1_n128 ) );
  NOR2_X1 \Check1_CheckInst_1_U130  ( .A1(\Check1_CheckInst_1_n126 ), .A2(
        \Check1_CheckInst_1_n125 ), .ZN(\Check1_CheckInst_1_n134 ) );
  XOR2_X1 \Check1_CheckInst_1_U129  ( .A(Red_AddRoundKeyOutput3[53]), .B(
        Red_SignaltoCheck[53]), .Z(\Check1_CheckInst_1_n125 ) );
  XOR2_X1 \Check1_CheckInst_1_U128  ( .A(Red_AddRoundKeyOutput2[1]), .B(
        Red_SignaltoCheck[65]), .Z(\Check1_CheckInst_1_n126 ) );
  NAND2_X1 \Check1_CheckInst_1_U127  ( .A1(\Check1_CheckInst_1_n124 ), .A2(
        \Check1_CheckInst_1_n123 ), .ZN(\Check1_CheckInst_1_n136 ) );
  XNOR2_X1 \Check1_CheckInst_1_U126  ( .A(Red_AddRoundKeyOutput2[37]), .B(
        Red_SignaltoCheck[101]), .ZN(\Check1_CheckInst_1_n123 ) );
  XNOR2_X1 \Check1_CheckInst_1_U125  ( .A(Red_AddRoundKeyOutput3[57]), .B(
        Red_SignaltoCheck[57]), .ZN(\Check1_CheckInst_1_n124 ) );
  NAND2_X1 \Check1_CheckInst_1_U124  ( .A1(\Check1_CheckInst_1_n122 ), .A2(
        \Check1_CheckInst_1_n121 ), .ZN(\Check1_CheckInst_1_n154 ) );
  NOR2_X1 \Check1_CheckInst_1_U123  ( .A1(\Check1_CheckInst_1_n120 ), .A2(
        \Check1_CheckInst_1_n119 ), .ZN(\Check1_CheckInst_1_n121 ) );
  NAND2_X1 \Check1_CheckInst_1_U122  ( .A1(\Check1_CheckInst_1_n118 ), .A2(
        \Check1_CheckInst_1_n117 ), .ZN(\Check1_CheckInst_1_n119 ) );
  NOR2_X1 \Check1_CheckInst_1_U121  ( .A1(\Check1_CheckInst_1_n116 ), .A2(
        \Check1_CheckInst_1_n115 ), .ZN(\Check1_CheckInst_1_n117 ) );
  XOR2_X1 \Check1_CheckInst_1_U120  ( .A(Red_AddRoundKeyOutput2[33]), .B(
        Red_SignaltoCheck[97]), .Z(\Check1_CheckInst_1_n115 ) );
  XOR2_X1 \Check1_CheckInst_1_U119  ( .A(Red_AddRoundKeyOutput2[41]), .B(
        Red_SignaltoCheck[105]), .Z(\Check1_CheckInst_1_n116 ) );
  NOR2_X1 \Check1_CheckInst_1_U118  ( .A1(\Check1_CheckInst_1_n114 ), .A2(
        \Check1_CheckInst_1_n113 ), .ZN(\Check1_CheckInst_1_n118 ) );
  XOR2_X1 \Check1_CheckInst_1_U117  ( .A(Red_AddRoundKeyOutput2[29]), .B(
        Red_SignaltoCheck[93]), .Z(\Check1_CheckInst_1_n113 ) );
  XOR2_X1 \Check1_CheckInst_1_U116  ( .A(Red_AddRoundKeyOutput2[25]), .B(
        Red_SignaltoCheck[89]), .Z(\Check1_CheckInst_1_n114 ) );
  NAND2_X1 \Check1_CheckInst_1_U115  ( .A1(\Check1_CheckInst_1_n112 ), .A2(
        \Check1_CheckInst_1_n111 ), .ZN(\Check1_CheckInst_1_n120 ) );
  XNOR2_X1 \Check1_CheckInst_1_U114  ( .A(Red_AddRoundKeyOutput2[21]), .B(
        Red_SignaltoCheck[85]), .ZN(\Check1_CheckInst_1_n111 ) );
  XNOR2_X1 \Check1_CheckInst_1_U113  ( .A(Red_AddRoundKeyOutput2[17]), .B(
        Red_SignaltoCheck[81]), .ZN(\Check1_CheckInst_1_n112 ) );
  NOR2_X1 \Check1_CheckInst_1_U112  ( .A1(\Check1_CheckInst_1_n110 ), .A2(
        \Check1_CheckInst_1_n109 ), .ZN(\Check1_CheckInst_1_n122 ) );
  XOR2_X1 \Check1_CheckInst_1_U111  ( .A(Red_AddRoundKeyOutput3[25]), .B(
        Red_SignaltoCheck[25]), .Z(\Check1_CheckInst_1_n109 ) );
  XOR2_X1 \Check1_CheckInst_1_U110  ( .A(Red_AddRoundKeyOutput3[37]), .B(
        Red_SignaltoCheck[37]), .Z(\Check1_CheckInst_1_n110 ) );
  NOR2_X1 \Check1_CheckInst_1_U109  ( .A1(\Check1_CheckInst_1_n108 ), .A2(
        \Check1_CheckInst_1_n107 ), .ZN(\Check1_CheckInst_1_n156 ) );
  NAND2_X1 \Check1_CheckInst_1_U108  ( .A1(\Check1_CheckInst_1_n106 ), .A2(
        \Check1_CheckInst_1_n105 ), .ZN(\Check1_CheckInst_1_n107 ) );
  NOR2_X1 \Check1_CheckInst_1_U107  ( .A1(\Check1_CheckInst_1_n104 ), .A2(
        \Check1_CheckInst_1_n103 ), .ZN(\Check1_CheckInst_1_n105 ) );
  NAND2_X1 \Check1_CheckInst_1_U106  ( .A1(\Check1_CheckInst_1_n102 ), .A2(
        \Check1_CheckInst_1_n101 ), .ZN(\Check1_CheckInst_1_n103 ) );
  XNOR2_X1 \Check1_CheckInst_1_U105  ( .A(Red_AddRoundKeyOutput3[29]), .B(
        Red_SignaltoCheck[29]), .ZN(\Check1_CheckInst_1_n101 ) );
  XNOR2_X1 \Check1_CheckInst_1_U104  ( .A(Red_AddRoundKeyOutput3[33]), .B(
        Red_SignaltoCheck[33]), .ZN(\Check1_CheckInst_1_n102 ) );
  NAND2_X1 \Check1_CheckInst_1_U103  ( .A1(\Check1_CheckInst_1_n100 ), .A2(
        \Check1_CheckInst_1_n99 ), .ZN(\Check1_CheckInst_1_n104 ) );
  XNOR2_X1 \Check1_CheckInst_1_U102  ( .A(Red_AddRoundKeyOutput3[45]), .B(
        Red_SignaltoCheck[45]), .ZN(\Check1_CheckInst_1_n99 ) );
  XNOR2_X1 \Check1_CheckInst_1_U101  ( .A(Red_AddRoundKeyOutput3[41]), .B(
        Red_SignaltoCheck[41]), .ZN(\Check1_CheckInst_1_n100 ) );
  NOR2_X1 \Check1_CheckInst_1_U100  ( .A1(\Check1_CheckInst_1_n98 ), .A2(
        \Check1_CheckInst_1_n97 ), .ZN(\Check1_CheckInst_1_n106 ) );
  XOR2_X1 \Check1_CheckInst_1_U99  ( .A(Red_AddRoundKeyOutput3[9]), .B(
        Red_SignaltoCheck[9]), .Z(\Check1_CheckInst_1_n97 ) );
  XOR2_X1 \Check1_CheckInst_1_U98  ( .A(Red_AddRoundKeyOutput3[49]), .B(
        Red_SignaltoCheck[49]), .Z(\Check1_CheckInst_1_n98 ) );
  NAND2_X1 \Check1_CheckInst_1_U97  ( .A1(\Check1_CheckInst_1_n96 ), .A2(
        \Check1_CheckInst_1_n95 ), .ZN(\Check1_CheckInst_1_n108 ) );
  XNOR2_X1 \Check1_CheckInst_1_U96  ( .A(Red_StateRegOutput[61]), .B(
        Red_SignaltoCheck[445]), .ZN(\Check1_CheckInst_1_n95 ) );
  XNOR2_X1 \Check1_CheckInst_1_U95  ( .A(Red_SignaltoCheck[1]), .B(
        Red_AddRoundKeyOutput3[1]), .ZN(\Check1_CheckInst_1_n96 ) );
  NOR2_X1 \Check1_CheckInst_1_U94  ( .A1(\Check1_CheckInst_1_n94 ), .A2(
        \Check1_CheckInst_1_n93 ), .ZN(\Check1_CheckInst_1_n222 ) );
  NAND2_X1 \Check1_CheckInst_1_U93  ( .A1(\Check1_CheckInst_1_n92 ), .A2(
        \Check1_CheckInst_1_n91 ), .ZN(\Check1_CheckInst_1_n93 ) );
  NOR2_X1 \Check1_CheckInst_1_U92  ( .A1(\Check1_CheckInst_1_n90 ), .A2(
        \Check1_CheckInst_1_n89 ), .ZN(\Check1_CheckInst_1_n91 ) );
  NAND2_X1 \Check1_CheckInst_1_U91  ( .A1(\Check1_CheckInst_1_n88 ), .A2(
        \Check1_CheckInst_1_n87 ), .ZN(\Check1_CheckInst_1_n89 ) );
  NOR2_X1 \Check1_CheckInst_1_U90  ( .A1(\Check1_CheckInst_1_n86 ), .A2(
        \Check1_CheckInst_1_n85 ), .ZN(\Check1_CheckInst_1_n87 ) );
  NAND2_X1 \Check1_CheckInst_1_U89  ( .A1(\Check1_CheckInst_1_n84 ), .A2(
        \Check1_CheckInst_1_n83 ), .ZN(\Check1_CheckInst_1_n85 ) );
  NOR2_X1 \Check1_CheckInst_1_U88  ( .A1(\Check1_CheckInst_1_n82 ), .A2(
        \Check1_CheckInst_1_n81 ), .ZN(\Check1_CheckInst_1_n83 ) );
  XOR2_X1 \Check1_CheckInst_1_U87  ( .A(Red_AddRoundKeyOutput3[13]), .B(
        Red_SignaltoCheck[13]), .Z(\Check1_CheckInst_1_n81 ) );
  XOR2_X1 \Check1_CheckInst_1_U86  ( .A(Red_SignaltoCheck[5]), .B(
        Red_AddRoundKeyOutput3[5]), .Z(\Check1_CheckInst_1_n82 ) );
  NOR2_X1 \Check1_CheckInst_1_U85  ( .A1(\Check1_CheckInst_1_n80 ), .A2(
        \Check1_CheckInst_1_n79 ), .ZN(\Check1_CheckInst_1_n84 ) );
  XOR2_X1 \Check1_CheckInst_1_U84  ( .A(Red_AddRoundKeyOutput3[21]), .B(
        Red_SignaltoCheck[21]), .Z(\Check1_CheckInst_1_n79 ) );
  XOR2_X1 \Check1_CheckInst_1_U83  ( .A(Red_AddRoundKeyOutput3[17]), .B(
        Red_SignaltoCheck[17]), .Z(\Check1_CheckInst_1_n80 ) );
  NAND2_X1 \Check1_CheckInst_1_U82  ( .A1(\Check1_CheckInst_1_n78 ), .A2(
        \Check1_CheckInst_1_n77 ), .ZN(\Check1_CheckInst_1_n86 ) );
  XNOR2_X1 \Check1_CheckInst_1_U81  ( .A(Red_AddRoundKeyOutput[61]), .B(
        Red_SignaltoCheck[189]), .ZN(\Check1_CheckInst_1_n77 ) );
  XNOR2_X1 \Check1_CheckInst_1_U80  ( .A(Red_AddRoundKeyOutput[57]), .B(
        Red_SignaltoCheck[185]), .ZN(\Check1_CheckInst_1_n78 ) );
  NOR2_X1 \Check1_CheckInst_1_U79  ( .A1(\Check1_CheckInst_1_n76 ), .A2(
        \Check1_CheckInst_1_n75 ), .ZN(\Check1_CheckInst_1_n88 ) );
  XOR2_X1 \Check1_CheckInst_1_U78  ( .A(Red_AddRoundKeyOutput[45]), .B(
        Red_SignaltoCheck[173]), .Z(\Check1_CheckInst_1_n75 ) );
  XOR2_X1 \Check1_CheckInst_1_U77  ( .A(Red_AddRoundKeyOutput[53]), .B(
        Red_SignaltoCheck[181]), .Z(\Check1_CheckInst_1_n76 ) );
  NAND2_X1 \Check1_CheckInst_1_U76  ( .A1(\Check1_CheckInst_1_n74 ), .A2(
        \Check1_CheckInst_1_n73 ), .ZN(\Check1_CheckInst_1_n90 ) );
  NOR2_X1 \Check1_CheckInst_1_U75  ( .A1(\Check1_CheckInst_1_n72 ), .A2(
        \Check1_CheckInst_1_n71 ), .ZN(\Check1_CheckInst_1_n73 ) );
  NAND2_X1 \Check1_CheckInst_1_U74  ( .A1(\Check1_CheckInst_1_n70 ), .A2(
        \Check1_CheckInst_1_n69 ), .ZN(\Check1_CheckInst_1_n71 ) );
  NOR2_X1 \Check1_CheckInst_1_U73  ( .A1(\Check1_CheckInst_1_n68 ), .A2(
        \Check1_CheckInst_1_n67 ), .ZN(\Check1_CheckInst_1_n69 ) );
  XOR2_X1 \Check1_CheckInst_1_U72  ( .A(Red_AddRoundKeyOutput[37]), .B(
        Red_SignaltoCheck[165]), .Z(\Check1_CheckInst_1_n67 ) );
  XOR2_X1 \Check1_CheckInst_1_U71  ( .A(Red_AddRoundKeyOutput[49]), .B(
        Red_SignaltoCheck[177]), .Z(\Check1_CheckInst_1_n68 ) );
  NOR2_X1 \Check1_CheckInst_1_U70  ( .A1(\Check1_CheckInst_1_n66 ), .A2(
        \Check1_CheckInst_1_n65 ), .ZN(\Check1_CheckInst_1_n70 ) );
  XOR2_X1 \Check1_CheckInst_1_U69  ( .A(Red_Feedback3[21]), .B(
        Red_SignaltoCheck[213]), .Z(\Check1_CheckInst_1_n65 ) );
  XOR2_X1 \Check1_CheckInst_1_U68  ( .A(Red_AddRoundKeyOutput[41]), .B(
        Red_SignaltoCheck[169]), .Z(\Check1_CheckInst_1_n66 ) );
  NAND2_X1 \Check1_CheckInst_1_U67  ( .A1(\Check1_CheckInst_1_n64 ), .A2(
        \Check1_CheckInst_1_n63 ), .ZN(\Check1_CheckInst_1_n72 ) );
  XNOR2_X1 \Check1_CheckInst_1_U66  ( .A(Red_Feedback3[17]), .B(
        Red_SignaltoCheck[209]), .ZN(\Check1_CheckInst_1_n63 ) );
  XNOR2_X1 \Check1_CheckInst_1_U65  ( .A(Red_Feedback3[25]), .B(
        Red_SignaltoCheck[217]), .ZN(\Check1_CheckInst_1_n64 ) );
  NOR2_X1 \Check1_CheckInst_1_U64  ( .A1(\Check1_CheckInst_1_n62 ), .A2(
        \Check1_CheckInst_1_n61 ), .ZN(\Check1_CheckInst_1_n74 ) );
  XOR2_X1 \Check1_CheckInst_1_U63  ( .A(Red_Feedback3[13]), .B(
        Red_SignaltoCheck[205]), .Z(\Check1_CheckInst_1_n61 ) );
  XOR2_X1 \Check1_CheckInst_1_U62  ( .A(Red_Feedback3[9]), .B(
        Red_SignaltoCheck[201]), .Z(\Check1_CheckInst_1_n62 ) );
  NOR2_X1 \Check1_CheckInst_1_U61  ( .A1(\Check1_CheckInst_1_n60 ), .A2(
        \Check1_CheckInst_1_n59 ), .ZN(\Check1_CheckInst_1_n92 ) );
  NAND2_X1 \Check1_CheckInst_1_U60  ( .A1(\Check1_CheckInst_1_n58 ), .A2(
        \Check1_CheckInst_1_n57 ), .ZN(\Check1_CheckInst_1_n59 ) );
  NOR2_X1 \Check1_CheckInst_1_U59  ( .A1(\Check1_CheckInst_1_n56 ), .A2(
        \Check1_CheckInst_1_n55 ), .ZN(\Check1_CheckInst_1_n57 ) );
  NAND2_X1 \Check1_CheckInst_1_U58  ( .A1(\Check1_CheckInst_1_n54 ), .A2(
        \Check1_CheckInst_1_n53 ), .ZN(\Check1_CheckInst_1_n55 ) );
  XNOR2_X1 \Check1_CheckInst_1_U57  ( .A(Red_Feedback3[5]), .B(
        Red_SignaltoCheck[197]), .ZN(\Check1_CheckInst_1_n53 ) );
  XNOR2_X1 \Check1_CheckInst_1_U56  ( .A(Red_Feedback3[1]), .B(
        Red_SignaltoCheck[193]), .ZN(\Check1_CheckInst_1_n54 ) );
  NAND2_X1 \Check1_CheckInst_1_U55  ( .A1(\Check1_CheckInst_1_n52 ), .A2(
        \Check1_CheckInst_1_n51 ), .ZN(\Check1_CheckInst_1_n56 ) );
  XNOR2_X1 \Check1_CheckInst_1_U54  ( .A(Red_AddRoundKeyOutput[5]), .B(
        Red_SignaltoCheck[133]), .ZN(\Check1_CheckInst_1_n51 ) );
  XNOR2_X1 \Check1_CheckInst_1_U53  ( .A(Red_AddRoundKeyOutput[1]), .B(
        Red_SignaltoCheck[129]), .ZN(\Check1_CheckInst_1_n52 ) );
  NOR2_X1 \Check1_CheckInst_1_U52  ( .A1(\Check1_CheckInst_1_n50 ), .A2(
        \Check1_CheckInst_1_n49 ), .ZN(\Check1_CheckInst_1_n58 ) );
  XOR2_X1 \Check1_CheckInst_1_U51  ( .A(Red_AddRoundKeyOutput2[53]), .B(
        Red_SignaltoCheck[117]), .Z(\Check1_CheckInst_1_n49 ) );
  XOR2_X1 \Check1_CheckInst_1_U50  ( .A(Red_AddRoundKeyOutput2[61]), .B(
        Red_SignaltoCheck[125]), .Z(\Check1_CheckInst_1_n50 ) );
  NAND2_X1 \Check1_CheckInst_1_U49  ( .A1(\Check1_CheckInst_1_n48 ), .A2(
        \Check1_CheckInst_1_n47 ), .ZN(\Check1_CheckInst_1_n60 ) );
  XNOR2_X1 \Check1_CheckInst_1_U48  ( .A(Red_AddRoundKeyOutput2[45]), .B(
        Red_SignaltoCheck[109]), .ZN(\Check1_CheckInst_1_n47 ) );
  XNOR2_X1 \Check1_CheckInst_1_U47  ( .A(Red_AddRoundKeyOutput2[57]), .B(
        Red_SignaltoCheck[121]), .ZN(\Check1_CheckInst_1_n48 ) );
  NAND2_X1 \Check1_CheckInst_1_U46  ( .A1(\Check1_CheckInst_1_n46 ), .A2(
        \Check1_CheckInst_1_n45 ), .ZN(\Check1_CheckInst_1_n94 ) );
  NOR2_X1 \Check1_CheckInst_1_U45  ( .A1(\Check1_CheckInst_1_n44 ), .A2(
        \Check1_CheckInst_1_n43 ), .ZN(\Check1_CheckInst_1_n45 ) );
  NAND2_X1 \Check1_CheckInst_1_U44  ( .A1(\Check1_CheckInst_1_n42 ), .A2(
        \Check1_CheckInst_1_n41 ), .ZN(\Check1_CheckInst_1_n43 ) );
  NOR2_X1 \Check1_CheckInst_1_U43  ( .A1(\Check1_CheckInst_1_n40 ), .A2(
        \Check1_CheckInst_1_n39 ), .ZN(\Check1_CheckInst_1_n41 ) );
  XOR2_X1 \Check1_CheckInst_1_U42  ( .A(Red_AddRoundKeyOutput[29]), .B(
        Red_SignaltoCheck[157]), .Z(\Check1_CheckInst_1_n39 ) );
  XOR2_X1 \Check1_CheckInst_1_U41  ( .A(Red_AddRoundKeyOutput2[49]), .B(
        Red_SignaltoCheck[113]), .Z(\Check1_CheckInst_1_n40 ) );
  NOR2_X1 \Check1_CheckInst_1_U40  ( .A1(\Check1_CheckInst_1_n38 ), .A2(
        \Check1_CheckInst_1_n37 ), .ZN(\Check1_CheckInst_1_n42 ) );
  XOR2_X1 \Check1_CheckInst_1_U39  ( .A(Red_AddRoundKeyOutput[25]), .B(
        Red_SignaltoCheck[153]), .Z(\Check1_CheckInst_1_n37 ) );
  XOR2_X1 \Check1_CheckInst_1_U38  ( .A(Red_AddRoundKeyOutput[33]), .B(
        Red_SignaltoCheck[161]), .Z(\Check1_CheckInst_1_n38 ) );
  NAND2_X1 \Check1_CheckInst_1_U37  ( .A1(\Check1_CheckInst_1_n36 ), .A2(
        \Check1_CheckInst_1_n35 ), .ZN(\Check1_CheckInst_1_n44 ) );
  XNOR2_X1 \Check1_CheckInst_1_U36  ( .A(Red_AddRoundKeyOutput[21]), .B(
        Red_SignaltoCheck[149]), .ZN(\Check1_CheckInst_1_n35 ) );
  XNOR2_X1 \Check1_CheckInst_1_U35  ( .A(Red_AddRoundKeyOutput[17]), .B(
        Red_SignaltoCheck[145]), .ZN(\Check1_CheckInst_1_n36 ) );
  NOR2_X1 \Check1_CheckInst_1_U34  ( .A1(\Check1_CheckInst_1_n34 ), .A2(
        \Check1_CheckInst_1_n33 ), .ZN(\Check1_CheckInst_1_n46 ) );
  XOR2_X1 \Check1_CheckInst_1_U33  ( .A(Red_AddRoundKeyOutput[13]), .B(
        Red_SignaltoCheck[141]), .Z(\Check1_CheckInst_1_n33 ) );
  XOR2_X1 \Check1_CheckInst_1_U32  ( .A(Red_AddRoundKeyOutput[9]), .B(
        Red_SignaltoCheck[137]), .Z(\Check1_CheckInst_1_n34 ) );
  NAND2_X1 \Check1_CheckInst_1_U31  ( .A1(\Check1_CheckInst_1_n32 ), .A2(
        \Check1_CheckInst_1_n31 ), .ZN(\Check1_CheckInst_1_n224 ) );
  NOR2_X1 \Check1_CheckInst_1_U30  ( .A1(\Check1_CheckInst_1_n30 ), .A2(
        \Check1_CheckInst_1_n29 ), .ZN(\Check1_CheckInst_1_n31 ) );
  NAND2_X1 \Check1_CheckInst_1_U29  ( .A1(\Check1_CheckInst_1_n28 ), .A2(
        \Check1_CheckInst_1_n27 ), .ZN(\Check1_CheckInst_1_n29 ) );
  NOR2_X1 \Check1_CheckInst_1_U28  ( .A1(\Check1_CheckInst_1_n26 ), .A2(
        \Check1_CheckInst_1_n25 ), .ZN(\Check1_CheckInst_1_n27 ) );
  NAND2_X1 \Check1_CheckInst_1_U27  ( .A1(\Check1_CheckInst_1_n24 ), .A2(
        \Check1_CheckInst_1_n23 ), .ZN(\Check1_CheckInst_1_n25 ) );
  XNOR2_X1 \Check1_CheckInst_1_U26  ( .A(Red_StateRegOutput3[29]), .B(
        Red_SignaltoCheck[285]), .ZN(\Check1_CheckInst_1_n23 ) );
  XNOR2_X1 \Check1_CheckInst_1_U25  ( .A(Red_StateRegOutput3[37]), .B(
        Red_SignaltoCheck[293]), .ZN(\Check1_CheckInst_1_n24 ) );
  NAND2_X1 \Check1_CheckInst_1_U24  ( .A1(\Check1_CheckInst_1_n22 ), .A2(
        \Check1_CheckInst_1_n21 ), .ZN(\Check1_CheckInst_1_n26 ) );
  XNOR2_X1 \Check1_CheckInst_1_U23  ( .A(Red_StateRegOutput3[45]), .B(
        Red_SignaltoCheck[301]), .ZN(\Check1_CheckInst_1_n21 ) );
  XNOR2_X1 \Check1_CheckInst_1_U22  ( .A(Red_StateRegOutput3[41]), .B(
        Red_SignaltoCheck[297]), .ZN(\Check1_CheckInst_1_n22 ) );
  NOR2_X1 \Check1_CheckInst_1_U21  ( .A1(\Check1_CheckInst_1_n20 ), .A2(
        \Check1_CheckInst_1_n19 ), .ZN(\Check1_CheckInst_1_n28 ) );
  NAND2_X1 \Check1_CheckInst_1_U20  ( .A1(\Check1_CheckInst_1_n18 ), .A2(
        \Check1_CheckInst_1_n17 ), .ZN(\Check1_CheckInst_1_n19 ) );
  XNOR2_X1 \Check1_CheckInst_1_U19  ( .A(Red_StateRegOutput2[5]), .B(
        Red_SignaltoCheck[325]), .ZN(\Check1_CheckInst_1_n17 ) );
  XNOR2_X1 \Check1_CheckInst_1_U18  ( .A(Red_StateRegOutput3[25]), .B(
        Red_SignaltoCheck[281]), .ZN(\Check1_CheckInst_1_n18 ) );
  NAND2_X1 \Check1_CheckInst_1_U17  ( .A1(\Check1_CheckInst_1_n16 ), .A2(
        \Check1_CheckInst_1_n15 ), .ZN(\Check1_CheckInst_1_n20 ) );
  XNOR2_X1 \Check1_CheckInst_1_U16  ( .A(Red_StateRegOutput3[21]), .B(
        Red_SignaltoCheck[277]), .ZN(\Check1_CheckInst_1_n15 ) );
  XNOR2_X1 \Check1_CheckInst_1_U15  ( .A(Red_StateRegOutput3[33]), .B(
        Red_SignaltoCheck[289]), .ZN(\Check1_CheckInst_1_n16 ) );
  NAND2_X1 \Check1_CheckInst_1_U14  ( .A1(\Check1_CheckInst_1_n14 ), .A2(
        \Check1_CheckInst_1_n13 ), .ZN(\Check1_CheckInst_1_n30 ) );
  NOR2_X1 \Check1_CheckInst_1_U13  ( .A1(\Check1_CheckInst_1_n12 ), .A2(
        \Check1_CheckInst_1_n11 ), .ZN(\Check1_CheckInst_1_n13 ) );
  XOR2_X1 \Check1_CheckInst_1_U12  ( .A(Red_StateRegOutput3[61]), .B(
        Red_SignaltoCheck[317]), .Z(\Check1_CheckInst_1_n11 ) );
  XOR2_X1 \Check1_CheckInst_1_U11  ( .A(Red_StateRegOutput3[57]), .B(
        Red_SignaltoCheck[313]), .Z(\Check1_CheckInst_1_n12 ) );
  NOR2_X1 \Check1_CheckInst_1_U10  ( .A1(\Check1_CheckInst_1_n10 ), .A2(
        \Check1_CheckInst_1_n9 ), .ZN(\Check1_CheckInst_1_n14 ) );
  XOR2_X1 \Check1_CheckInst_1_U9  ( .A(Red_StateRegOutput2[1]), .B(
        Red_SignaltoCheck[321]), .Z(\Check1_CheckInst_1_n9 ) );
  XOR2_X1 \Check1_CheckInst_1_U8  ( .A(Red_StateRegOutput2[9]), .B(
        Red_SignaltoCheck[329]), .Z(\Check1_CheckInst_1_n10 ) );
  NOR2_X1 \Check1_CheckInst_1_U7  ( .A1(\Check1_CheckInst_1_n8 ), .A2(
        \Check1_CheckInst_1_n7 ), .ZN(\Check1_CheckInst_1_n32 ) );
  NAND2_X1 \Check1_CheckInst_1_U6  ( .A1(\Check1_CheckInst_1_n6 ), .A2(
        \Check1_CheckInst_1_n5 ), .ZN(\Check1_CheckInst_1_n7 ) );
  XNOR2_X1 \Check1_CheckInst_1_U5  ( .A(Red_Feedback3[53]), .B(
        Red_SignaltoCheck[245]), .ZN(\Check1_CheckInst_1_n5 ) );
  XNOR2_X1 \Check1_CheckInst_1_U4  ( .A(Red_Feedback3[49]), .B(
        Red_SignaltoCheck[241]), .ZN(\Check1_CheckInst_1_n6 ) );
  NAND2_X1 \Check1_CheckInst_1_U3  ( .A1(\Check1_CheckInst_1_n4 ), .A2(
        \Check1_CheckInst_1_n3 ), .ZN(\Check1_CheckInst_1_n8 ) );
  XNOR2_X1 \Check1_CheckInst_1_U2  ( .A(Red_StateRegOutput3[53]), .B(
        Red_SignaltoCheck[309]), .ZN(\Check1_CheckInst_1_n3 ) );
  XNOR2_X1 \Check1_CheckInst_1_U1  ( .A(Red_StateRegOutput3[49]), .B(
        Red_SignaltoCheck[305]), .ZN(\Check1_CheckInst_1_n4 ) );
  NOR2_X1 \Check1_CheckInst_2_U223  ( .A1(\Check1_CheckInst_2_n224 ), .A2(
        \Check1_CheckInst_2_n223 ), .ZN(Error[2]) );
  NAND2_X1 \Check1_CheckInst_2_U222  ( .A1(\Check1_CheckInst_2_n222 ), .A2(
        \Check1_CheckInst_2_n221 ), .ZN(\Check1_CheckInst_2_n223 ) );
  NOR2_X1 \Check1_CheckInst_2_U221  ( .A1(\Check1_CheckInst_2_n220 ), .A2(
        \Check1_CheckInst_2_n219 ), .ZN(\Check1_CheckInst_2_n221 ) );
  NAND2_X1 \Check1_CheckInst_2_U220  ( .A1(\Check1_CheckInst_2_n218 ), .A2(
        \Check1_CheckInst_2_n217 ), .ZN(\Check1_CheckInst_2_n219 ) );
  NOR2_X1 \Check1_CheckInst_2_U219  ( .A1(\Check1_CheckInst_2_n216 ), .A2(
        \Check1_CheckInst_2_n215 ), .ZN(\Check1_CheckInst_2_n217 ) );
  NAND2_X1 \Check1_CheckInst_2_U218  ( .A1(\Check1_CheckInst_2_n214 ), .A2(
        \Check1_CheckInst_2_n213 ), .ZN(\Check1_CheckInst_2_n215 ) );
  NOR2_X1 \Check1_CheckInst_2_U217  ( .A1(\Check1_CheckInst_2_n212 ), .A2(
        \Check1_CheckInst_2_n211 ), .ZN(\Check1_CheckInst_2_n213 ) );
  NAND2_X1 \Check1_CheckInst_2_U216  ( .A1(\Check1_CheckInst_2_n210 ), .A2(
        \Check1_CheckInst_2_n209 ), .ZN(\Check1_CheckInst_2_n211 ) );
  NOR2_X1 \Check1_CheckInst_2_U215  ( .A1(\Check1_CheckInst_2_n208 ), .A2(
        \Check1_CheckInst_2_n207 ), .ZN(\Check1_CheckInst_2_n209 ) );
  NAND2_X1 \Check1_CheckInst_2_U214  ( .A1(\Check1_CheckInst_2_n206 ), .A2(
        \Check1_CheckInst_2_n205 ), .ZN(\Check1_CheckInst_2_n207 ) );
  XNOR2_X1 \Check1_CheckInst_2_U213  ( .A(Red_Feedback3[38]), .B(
        Red_SignaltoCheck[230]), .ZN(\Check1_CheckInst_2_n205 ) );
  XNOR2_X1 \Check1_CheckInst_2_U212  ( .A(Red_Feedback3[46]), .B(
        Red_SignaltoCheck[238]), .ZN(\Check1_CheckInst_2_n206 ) );
  NAND2_X1 \Check1_CheckInst_2_U211  ( .A1(\Check1_CheckInst_2_n204 ), .A2(
        \Check1_CheckInst_2_n203 ), .ZN(\Check1_CheckInst_2_n208 ) );
  XNOR2_X1 \Check1_CheckInst_2_U210  ( .A(Red_Feedback3[30]), .B(
        Red_SignaltoCheck[222]), .ZN(\Check1_CheckInst_2_n203 ) );
  XNOR2_X1 \Check1_CheckInst_2_U209  ( .A(Red_Feedback3[42]), .B(
        Red_SignaltoCheck[234]), .ZN(\Check1_CheckInst_2_n204 ) );
  NOR2_X1 \Check1_CheckInst_2_U208  ( .A1(\Check1_CheckInst_2_n202 ), .A2(
        \Check1_CheckInst_2_n201 ), .ZN(\Check1_CheckInst_2_n210 ) );
  XOR2_X1 \Check1_CheckInst_2_U207  ( .A(Red_StateRegOutput3[14]), .B(
        Red_SignaltoCheck[270]), .Z(\Check1_CheckInst_2_n201 ) );
  XOR2_X1 \Check1_CheckInst_2_U206  ( .A(Red_Feedback3[34]), .B(
        Red_SignaltoCheck[226]), .Z(\Check1_CheckInst_2_n202 ) );
  NAND2_X1 \Check1_CheckInst_2_U205  ( .A1(\Check1_CheckInst_2_n200 ), .A2(
        \Check1_CheckInst_2_n199 ), .ZN(\Check1_CheckInst_2_n212 ) );
  XNOR2_X1 \Check1_CheckInst_2_U204  ( .A(Red_StateRegOutput3[10]), .B(
        Red_SignaltoCheck[266]), .ZN(\Check1_CheckInst_2_n199 ) );
  XNOR2_X1 \Check1_CheckInst_2_U203  ( .A(Red_StateRegOutput3[18]), .B(
        Red_SignaltoCheck[274]), .ZN(\Check1_CheckInst_2_n200 ) );
  NOR2_X1 \Check1_CheckInst_2_U202  ( .A1(\Check1_CheckInst_2_n198 ), .A2(
        \Check1_CheckInst_2_n197 ), .ZN(\Check1_CheckInst_2_n214 ) );
  NAND2_X1 \Check1_CheckInst_2_U201  ( .A1(\Check1_CheckInst_2_n196 ), .A2(
        \Check1_CheckInst_2_n195 ), .ZN(\Check1_CheckInst_2_n197 ) );
  NOR2_X1 \Check1_CheckInst_2_U200  ( .A1(\Check1_CheckInst_2_n194 ), .A2(
        \Check1_CheckInst_2_n193 ), .ZN(\Check1_CheckInst_2_n195 ) );
  NAND2_X1 \Check1_CheckInst_2_U199  ( .A1(\Check1_CheckInst_2_n192 ), .A2(
        \Check1_CheckInst_2_n191 ), .ZN(\Check1_CheckInst_2_n193 ) );
  XNOR2_X1 \Check1_CheckInst_2_U198  ( .A(Red_StateRegOutput3[6]), .B(
        Red_SignaltoCheck[262]), .ZN(\Check1_CheckInst_2_n191 ) );
  XNOR2_X1 \Check1_CheckInst_2_U197  ( .A(Red_StateRegOutput3[2]), .B(
        Red_SignaltoCheck[258]), .ZN(\Check1_CheckInst_2_n192 ) );
  NAND2_X1 \Check1_CheckInst_2_U196  ( .A1(\Check1_CheckInst_2_n190 ), .A2(
        \Check1_CheckInst_2_n189 ), .ZN(\Check1_CheckInst_2_n194 ) );
  XNOR2_X1 \Check1_CheckInst_2_U195  ( .A(Red_Feedback3[62]), .B(
        Red_SignaltoCheck[254]), .ZN(\Check1_CheckInst_2_n189 ) );
  XNOR2_X1 \Check1_CheckInst_2_U194  ( .A(Red_Feedback3[58]), .B(
        Red_SignaltoCheck[250]), .ZN(\Check1_CheckInst_2_n190 ) );
  NOR2_X1 \Check1_CheckInst_2_U193  ( .A1(\Check1_CheckInst_2_n188 ), .A2(
        \Check1_CheckInst_2_n187 ), .ZN(\Check1_CheckInst_2_n196 ) );
  XOR2_X1 \Check1_CheckInst_2_U192  ( .A(Red_StateRegOutput[30]), .B(
        Red_SignaltoCheck[414]), .Z(\Check1_CheckInst_2_n187 ) );
  XOR2_X1 \Check1_CheckInst_2_U191  ( .A(Red_StateRegOutput[26]), .B(
        Red_SignaltoCheck[410]), .Z(\Check1_CheckInst_2_n188 ) );
  NAND2_X1 \Check1_CheckInst_2_U190  ( .A1(\Check1_CheckInst_2_n186 ), .A2(
        \Check1_CheckInst_2_n185 ), .ZN(\Check1_CheckInst_2_n198 ) );
  XNOR2_X1 \Check1_CheckInst_2_U189  ( .A(Red_StateRegOutput[14]), .B(
        Red_SignaltoCheck[398]), .ZN(\Check1_CheckInst_2_n185 ) );
  XNOR2_X1 \Check1_CheckInst_2_U188  ( .A(Red_StateRegOutput[22]), .B(
        Red_SignaltoCheck[406]), .ZN(\Check1_CheckInst_2_n186 ) );
  NAND2_X1 \Check1_CheckInst_2_U187  ( .A1(\Check1_CheckInst_2_n184 ), .A2(
        \Check1_CheckInst_2_n183 ), .ZN(\Check1_CheckInst_2_n216 ) );
  NOR2_X1 \Check1_CheckInst_2_U186  ( .A1(\Check1_CheckInst_2_n182 ), .A2(
        \Check1_CheckInst_2_n181 ), .ZN(\Check1_CheckInst_2_n183 ) );
  NAND2_X1 \Check1_CheckInst_2_U185  ( .A1(\Check1_CheckInst_2_n180 ), .A2(
        \Check1_CheckInst_2_n179 ), .ZN(\Check1_CheckInst_2_n181 ) );
  NOR2_X1 \Check1_CheckInst_2_U184  ( .A1(\Check1_CheckInst_2_n178 ), .A2(
        \Check1_CheckInst_2_n177 ), .ZN(\Check1_CheckInst_2_n179 ) );
  XOR2_X1 \Check1_CheckInst_2_U183  ( .A(Red_StateRegOutput[6]), .B(
        Red_SignaltoCheck[390]), .Z(\Check1_CheckInst_2_n177 ) );
  XOR2_X1 \Check1_CheckInst_2_U182  ( .A(Red_StateRegOutput[18]), .B(
        Red_SignaltoCheck[402]), .Z(\Check1_CheckInst_2_n178 ) );
  NOR2_X1 \Check1_CheckInst_2_U181  ( .A1(\Check1_CheckInst_2_n176 ), .A2(
        \Check1_CheckInst_2_n175 ), .ZN(\Check1_CheckInst_2_n180 ) );
  XOR2_X1 \Check1_CheckInst_2_U180  ( .A(Red_StateRegOutput[54]), .B(
        Red_SignaltoCheck[438]), .Z(\Check1_CheckInst_2_n175 ) );
  XOR2_X1 \Check1_CheckInst_2_U179  ( .A(Red_StateRegOutput[10]), .B(
        Red_SignaltoCheck[394]), .Z(\Check1_CheckInst_2_n176 ) );
  NAND2_X1 \Check1_CheckInst_2_U178  ( .A1(\Check1_CheckInst_2_n174 ), .A2(
        \Check1_CheckInst_2_n173 ), .ZN(\Check1_CheckInst_2_n182 ) );
  XNOR2_X1 \Check1_CheckInst_2_U177  ( .A(Red_StateRegOutput[50]), .B(
        Red_SignaltoCheck[434]), .ZN(\Check1_CheckInst_2_n173 ) );
  XNOR2_X1 \Check1_CheckInst_2_U176  ( .A(Red_StateRegOutput[58]), .B(
        Red_SignaltoCheck[442]), .ZN(\Check1_CheckInst_2_n174 ) );
  NOR2_X1 \Check1_CheckInst_2_U175  ( .A1(\Check1_CheckInst_2_n172 ), .A2(
        \Check1_CheckInst_2_n171 ), .ZN(\Check1_CheckInst_2_n184 ) );
  XOR2_X1 \Check1_CheckInst_2_U174  ( .A(Red_StateRegOutput[46]), .B(
        Red_SignaltoCheck[430]), .Z(\Check1_CheckInst_2_n171 ) );
  XOR2_X1 \Check1_CheckInst_2_U173  ( .A(Red_StateRegOutput[42]), .B(
        Red_SignaltoCheck[426]), .Z(\Check1_CheckInst_2_n172 ) );
  NOR2_X1 \Check1_CheckInst_2_U172  ( .A1(\Check1_CheckInst_2_n170 ), .A2(
        \Check1_CheckInst_2_n169 ), .ZN(\Check1_CheckInst_2_n218 ) );
  NAND2_X1 \Check1_CheckInst_2_U171  ( .A1(\Check1_CheckInst_2_n168 ), .A2(
        \Check1_CheckInst_2_n167 ), .ZN(\Check1_CheckInst_2_n169 ) );
  NOR2_X1 \Check1_CheckInst_2_U170  ( .A1(\Check1_CheckInst_2_n166 ), .A2(
        \Check1_CheckInst_2_n165 ), .ZN(\Check1_CheckInst_2_n167 ) );
  NAND2_X1 \Check1_CheckInst_2_U169  ( .A1(\Check1_CheckInst_2_n164 ), .A2(
        \Check1_CheckInst_2_n163 ), .ZN(\Check1_CheckInst_2_n165 ) );
  XNOR2_X1 \Check1_CheckInst_2_U168  ( .A(Red_StateRegOutput[38]), .B(
        Red_SignaltoCheck[422]), .ZN(\Check1_CheckInst_2_n163 ) );
  XNOR2_X1 \Check1_CheckInst_2_U167  ( .A(Red_StateRegOutput[34]), .B(
        Red_SignaltoCheck[418]), .ZN(\Check1_CheckInst_2_n164 ) );
  NAND2_X1 \Check1_CheckInst_2_U166  ( .A1(\Check1_CheckInst_2_n162 ), .A2(
        \Check1_CheckInst_2_n161 ), .ZN(\Check1_CheckInst_2_n166 ) );
  XNOR2_X1 \Check1_CheckInst_2_U165  ( .A(Red_StateRegOutput2[38]), .B(
        Red_SignaltoCheck[358]), .ZN(\Check1_CheckInst_2_n161 ) );
  XNOR2_X1 \Check1_CheckInst_2_U164  ( .A(Red_StateRegOutput2[34]), .B(
        Red_SignaltoCheck[354]), .ZN(\Check1_CheckInst_2_n162 ) );
  NOR2_X1 \Check1_CheckInst_2_U163  ( .A1(\Check1_CheckInst_2_n160 ), .A2(
        \Check1_CheckInst_2_n159 ), .ZN(\Check1_CheckInst_2_n168 ) );
  XOR2_X1 \Check1_CheckInst_2_U162  ( .A(Red_StateRegOutput2[22]), .B(
        Red_SignaltoCheck[342]), .Z(\Check1_CheckInst_2_n159 ) );
  XOR2_X1 \Check1_CheckInst_2_U161  ( .A(Red_StateRegOutput2[30]), .B(
        Red_SignaltoCheck[350]), .Z(\Check1_CheckInst_2_n160 ) );
  NAND2_X1 \Check1_CheckInst_2_U160  ( .A1(\Check1_CheckInst_2_n158 ), .A2(
        \Check1_CheckInst_2_n157 ), .ZN(\Check1_CheckInst_2_n170 ) );
  XNOR2_X1 \Check1_CheckInst_2_U159  ( .A(Red_StateRegOutput2[14]), .B(
        Red_SignaltoCheck[334]), .ZN(\Check1_CheckInst_2_n157 ) );
  XNOR2_X1 \Check1_CheckInst_2_U158  ( .A(Red_StateRegOutput2[26]), .B(
        Red_SignaltoCheck[346]), .ZN(\Check1_CheckInst_2_n158 ) );
  NAND2_X1 \Check1_CheckInst_2_U157  ( .A1(\Check1_CheckInst_2_n156 ), .A2(
        \Check1_CheckInst_2_n155 ), .ZN(\Check1_CheckInst_2_n220 ) );
  NOR2_X1 \Check1_CheckInst_2_U156  ( .A1(\Check1_CheckInst_2_n154 ), .A2(
        \Check1_CheckInst_2_n153 ), .ZN(\Check1_CheckInst_2_n155 ) );
  NAND2_X1 \Check1_CheckInst_2_U155  ( .A1(\Check1_CheckInst_2_n152 ), .A2(
        \Check1_CheckInst_2_n151 ), .ZN(\Check1_CheckInst_2_n153 ) );
  NOR2_X1 \Check1_CheckInst_2_U154  ( .A1(\Check1_CheckInst_2_n150 ), .A2(
        \Check1_CheckInst_2_n149 ), .ZN(\Check1_CheckInst_2_n151 ) );
  NAND2_X1 \Check1_CheckInst_2_U153  ( .A1(\Check1_CheckInst_2_n148 ), .A2(
        \Check1_CheckInst_2_n147 ), .ZN(\Check1_CheckInst_2_n149 ) );
  NOR2_X1 \Check1_CheckInst_2_U152  ( .A1(\Check1_CheckInst_2_n146 ), .A2(
        \Check1_CheckInst_2_n145 ), .ZN(\Check1_CheckInst_2_n147 ) );
  NAND2_X1 \Check1_CheckInst_2_U151  ( .A1(\Check1_CheckInst_2_n144 ), .A2(
        \Check1_CheckInst_2_n143 ), .ZN(\Check1_CheckInst_2_n145 ) );
  XNOR2_X1 \Check1_CheckInst_2_U150  ( .A(Red_StateRegOutput2[62]), .B(
        Red_SignaltoCheck[382]), .ZN(\Check1_CheckInst_2_n143 ) );
  XNOR2_X1 \Check1_CheckInst_2_U149  ( .A(Red_StateRegOutput2[18]), .B(
        Red_SignaltoCheck[338]), .ZN(\Check1_CheckInst_2_n144 ) );
  NAND2_X1 \Check1_CheckInst_2_U148  ( .A1(\Check1_CheckInst_2_n142 ), .A2(
        \Check1_CheckInst_2_n141 ), .ZN(\Check1_CheckInst_2_n146 ) );
  XNOR2_X1 \Check1_CheckInst_2_U147  ( .A(Red_StateRegOutput2[58]), .B(
        Red_SignaltoCheck[378]), .ZN(\Check1_CheckInst_2_n141 ) );
  XNOR2_X1 \Check1_CheckInst_2_U146  ( .A(Red_StateRegOutput[2]), .B(
        Red_SignaltoCheck[386]), .ZN(\Check1_CheckInst_2_n142 ) );
  NOR2_X1 \Check1_CheckInst_2_U145  ( .A1(\Check1_CheckInst_2_n140 ), .A2(
        \Check1_CheckInst_2_n139 ), .ZN(\Check1_CheckInst_2_n148 ) );
  XOR2_X1 \Check1_CheckInst_2_U144  ( .A(Red_StateRegOutput2[54]), .B(
        Red_SignaltoCheck[374]), .Z(\Check1_CheckInst_2_n139 ) );
  XOR2_X1 \Check1_CheckInst_2_U143  ( .A(Red_StateRegOutput2[50]), .B(
        Red_SignaltoCheck[370]), .Z(\Check1_CheckInst_2_n140 ) );
  NAND2_X1 \Check1_CheckInst_2_U142  ( .A1(\Check1_CheckInst_2_n138 ), .A2(
        \Check1_CheckInst_2_n137 ), .ZN(\Check1_CheckInst_2_n150 ) );
  XNOR2_X1 \Check1_CheckInst_2_U141  ( .A(Red_StateRegOutput2[46]), .B(
        Red_SignaltoCheck[366]), .ZN(\Check1_CheckInst_2_n137 ) );
  XNOR2_X1 \Check1_CheckInst_2_U140  ( .A(Red_StateRegOutput2[42]), .B(
        Red_SignaltoCheck[362]), .ZN(\Check1_CheckInst_2_n138 ) );
  NOR2_X1 \Check1_CheckInst_2_U139  ( .A1(\Check1_CheckInst_2_n136 ), .A2(
        \Check1_CheckInst_2_n135 ), .ZN(\Check1_CheckInst_2_n152 ) );
  NAND2_X1 \Check1_CheckInst_2_U138  ( .A1(\Check1_CheckInst_2_n134 ), .A2(
        \Check1_CheckInst_2_n133 ), .ZN(\Check1_CheckInst_2_n135 ) );
  NOR2_X1 \Check1_CheckInst_2_U137  ( .A1(\Check1_CheckInst_2_n132 ), .A2(
        \Check1_CheckInst_2_n131 ), .ZN(\Check1_CheckInst_2_n133 ) );
  NAND2_X1 \Check1_CheckInst_2_U136  ( .A1(\Check1_CheckInst_2_n130 ), .A2(
        \Check1_CheckInst_2_n129 ), .ZN(\Check1_CheckInst_2_n131 ) );
  XNOR2_X1 \Check1_CheckInst_2_U135  ( .A(Red_AddRoundKeyOutput2[14]), .B(
        Red_SignaltoCheck[78]), .ZN(\Check1_CheckInst_2_n129 ) );
  XNOR2_X1 \Check1_CheckInst_2_U134  ( .A(Red_AddRoundKeyOutput2[10]), .B(
        Red_SignaltoCheck[74]), .ZN(\Check1_CheckInst_2_n130 ) );
  NAND2_X1 \Check1_CheckInst_2_U133  ( .A1(\Check1_CheckInst_2_n128 ), .A2(
        \Check1_CheckInst_2_n127 ), .ZN(\Check1_CheckInst_2_n132 ) );
  XNOR2_X1 \Check1_CheckInst_2_U132  ( .A(Red_AddRoundKeyOutput3[62]), .B(
        Red_SignaltoCheck[62]), .ZN(\Check1_CheckInst_2_n127 ) );
  XNOR2_X1 \Check1_CheckInst_2_U131  ( .A(Red_AddRoundKeyOutput2[6]), .B(
        Red_SignaltoCheck[70]), .ZN(\Check1_CheckInst_2_n128 ) );
  NOR2_X1 \Check1_CheckInst_2_U130  ( .A1(\Check1_CheckInst_2_n126 ), .A2(
        \Check1_CheckInst_2_n125 ), .ZN(\Check1_CheckInst_2_n134 ) );
  XOR2_X1 \Check1_CheckInst_2_U129  ( .A(Red_AddRoundKeyOutput3[54]), .B(
        Red_SignaltoCheck[54]), .Z(\Check1_CheckInst_2_n125 ) );
  XOR2_X1 \Check1_CheckInst_2_U128  ( .A(Red_AddRoundKeyOutput2[2]), .B(
        Red_SignaltoCheck[66]), .Z(\Check1_CheckInst_2_n126 ) );
  NAND2_X1 \Check1_CheckInst_2_U127  ( .A1(\Check1_CheckInst_2_n124 ), .A2(
        \Check1_CheckInst_2_n123 ), .ZN(\Check1_CheckInst_2_n136 ) );
  XNOR2_X1 \Check1_CheckInst_2_U126  ( .A(Red_AddRoundKeyOutput2[38]), .B(
        Red_SignaltoCheck[102]), .ZN(\Check1_CheckInst_2_n123 ) );
  XNOR2_X1 \Check1_CheckInst_2_U125  ( .A(Red_AddRoundKeyOutput3[58]), .B(
        Red_SignaltoCheck[58]), .ZN(\Check1_CheckInst_2_n124 ) );
  NAND2_X1 \Check1_CheckInst_2_U124  ( .A1(\Check1_CheckInst_2_n122 ), .A2(
        \Check1_CheckInst_2_n121 ), .ZN(\Check1_CheckInst_2_n154 ) );
  NOR2_X1 \Check1_CheckInst_2_U123  ( .A1(\Check1_CheckInst_2_n120 ), .A2(
        \Check1_CheckInst_2_n119 ), .ZN(\Check1_CheckInst_2_n121 ) );
  NAND2_X1 \Check1_CheckInst_2_U122  ( .A1(\Check1_CheckInst_2_n118 ), .A2(
        \Check1_CheckInst_2_n117 ), .ZN(\Check1_CheckInst_2_n119 ) );
  NOR2_X1 \Check1_CheckInst_2_U121  ( .A1(\Check1_CheckInst_2_n116 ), .A2(
        \Check1_CheckInst_2_n115 ), .ZN(\Check1_CheckInst_2_n117 ) );
  XOR2_X1 \Check1_CheckInst_2_U120  ( .A(Red_AddRoundKeyOutput2[34]), .B(
        Red_SignaltoCheck[98]), .Z(\Check1_CheckInst_2_n115 ) );
  XOR2_X1 \Check1_CheckInst_2_U119  ( .A(Red_AddRoundKeyOutput2[42]), .B(
        Red_SignaltoCheck[106]), .Z(\Check1_CheckInst_2_n116 ) );
  NOR2_X1 \Check1_CheckInst_2_U118  ( .A1(\Check1_CheckInst_2_n114 ), .A2(
        \Check1_CheckInst_2_n113 ), .ZN(\Check1_CheckInst_2_n118 ) );
  XOR2_X1 \Check1_CheckInst_2_U117  ( .A(Red_AddRoundKeyOutput2[30]), .B(
        Red_SignaltoCheck[94]), .Z(\Check1_CheckInst_2_n113 ) );
  XOR2_X1 \Check1_CheckInst_2_U116  ( .A(Red_AddRoundKeyOutput2[26]), .B(
        Red_SignaltoCheck[90]), .Z(\Check1_CheckInst_2_n114 ) );
  NAND2_X1 \Check1_CheckInst_2_U115  ( .A1(\Check1_CheckInst_2_n112 ), .A2(
        \Check1_CheckInst_2_n111 ), .ZN(\Check1_CheckInst_2_n120 ) );
  XNOR2_X1 \Check1_CheckInst_2_U114  ( .A(Red_AddRoundKeyOutput2[22]), .B(
        Red_SignaltoCheck[86]), .ZN(\Check1_CheckInst_2_n111 ) );
  XNOR2_X1 \Check1_CheckInst_2_U113  ( .A(Red_AddRoundKeyOutput2[18]), .B(
        Red_SignaltoCheck[82]), .ZN(\Check1_CheckInst_2_n112 ) );
  NOR2_X1 \Check1_CheckInst_2_U112  ( .A1(\Check1_CheckInst_2_n110 ), .A2(
        \Check1_CheckInst_2_n109 ), .ZN(\Check1_CheckInst_2_n122 ) );
  XOR2_X1 \Check1_CheckInst_2_U111  ( .A(Red_AddRoundKeyOutput3[26]), .B(
        Red_SignaltoCheck[26]), .Z(\Check1_CheckInst_2_n109 ) );
  XOR2_X1 \Check1_CheckInst_2_U110  ( .A(Red_AddRoundKeyOutput3[38]), .B(
        Red_SignaltoCheck[38]), .Z(\Check1_CheckInst_2_n110 ) );
  NOR2_X1 \Check1_CheckInst_2_U109  ( .A1(\Check1_CheckInst_2_n108 ), .A2(
        \Check1_CheckInst_2_n107 ), .ZN(\Check1_CheckInst_2_n156 ) );
  NAND2_X1 \Check1_CheckInst_2_U108  ( .A1(\Check1_CheckInst_2_n106 ), .A2(
        \Check1_CheckInst_2_n105 ), .ZN(\Check1_CheckInst_2_n107 ) );
  NOR2_X1 \Check1_CheckInst_2_U107  ( .A1(\Check1_CheckInst_2_n104 ), .A2(
        \Check1_CheckInst_2_n103 ), .ZN(\Check1_CheckInst_2_n105 ) );
  NAND2_X1 \Check1_CheckInst_2_U106  ( .A1(\Check1_CheckInst_2_n102 ), .A2(
        \Check1_CheckInst_2_n101 ), .ZN(\Check1_CheckInst_2_n103 ) );
  XNOR2_X1 \Check1_CheckInst_2_U105  ( .A(Red_AddRoundKeyOutput3[30]), .B(
        Red_SignaltoCheck[30]), .ZN(\Check1_CheckInst_2_n101 ) );
  XNOR2_X1 \Check1_CheckInst_2_U104  ( .A(Red_AddRoundKeyOutput3[34]), .B(
        Red_SignaltoCheck[34]), .ZN(\Check1_CheckInst_2_n102 ) );
  NAND2_X1 \Check1_CheckInst_2_U103  ( .A1(\Check1_CheckInst_2_n100 ), .A2(
        \Check1_CheckInst_2_n99 ), .ZN(\Check1_CheckInst_2_n104 ) );
  XNOR2_X1 \Check1_CheckInst_2_U102  ( .A(Red_AddRoundKeyOutput3[46]), .B(
        Red_SignaltoCheck[46]), .ZN(\Check1_CheckInst_2_n99 ) );
  XNOR2_X1 \Check1_CheckInst_2_U101  ( .A(Red_AddRoundKeyOutput3[42]), .B(
        Red_SignaltoCheck[42]), .ZN(\Check1_CheckInst_2_n100 ) );
  NOR2_X1 \Check1_CheckInst_2_U100  ( .A1(\Check1_CheckInst_2_n98 ), .A2(
        \Check1_CheckInst_2_n97 ), .ZN(\Check1_CheckInst_2_n106 ) );
  XOR2_X1 \Check1_CheckInst_2_U99  ( .A(Red_AddRoundKeyOutput3[10]), .B(
        Red_SignaltoCheck[10]), .Z(\Check1_CheckInst_2_n97 ) );
  XOR2_X1 \Check1_CheckInst_2_U98  ( .A(Red_AddRoundKeyOutput3[50]), .B(
        Red_SignaltoCheck[50]), .Z(\Check1_CheckInst_2_n98 ) );
  NAND2_X1 \Check1_CheckInst_2_U97  ( .A1(\Check1_CheckInst_2_n96 ), .A2(
        \Check1_CheckInst_2_n95 ), .ZN(\Check1_CheckInst_2_n108 ) );
  XNOR2_X1 \Check1_CheckInst_2_U96  ( .A(Red_StateRegOutput[62]), .B(
        Red_SignaltoCheck[446]), .ZN(\Check1_CheckInst_2_n95 ) );
  XNOR2_X1 \Check1_CheckInst_2_U95  ( .A(Red_SignaltoCheck[2]), .B(
        Red_AddRoundKeyOutput3[2]), .ZN(\Check1_CheckInst_2_n96 ) );
  NOR2_X1 \Check1_CheckInst_2_U94  ( .A1(\Check1_CheckInst_2_n94 ), .A2(
        \Check1_CheckInst_2_n93 ), .ZN(\Check1_CheckInst_2_n222 ) );
  NAND2_X1 \Check1_CheckInst_2_U93  ( .A1(\Check1_CheckInst_2_n92 ), .A2(
        \Check1_CheckInst_2_n91 ), .ZN(\Check1_CheckInst_2_n93 ) );
  NOR2_X1 \Check1_CheckInst_2_U92  ( .A1(\Check1_CheckInst_2_n90 ), .A2(
        \Check1_CheckInst_2_n89 ), .ZN(\Check1_CheckInst_2_n91 ) );
  NAND2_X1 \Check1_CheckInst_2_U91  ( .A1(\Check1_CheckInst_2_n88 ), .A2(
        \Check1_CheckInst_2_n87 ), .ZN(\Check1_CheckInst_2_n89 ) );
  NOR2_X1 \Check1_CheckInst_2_U90  ( .A1(\Check1_CheckInst_2_n86 ), .A2(
        \Check1_CheckInst_2_n85 ), .ZN(\Check1_CheckInst_2_n87 ) );
  NAND2_X1 \Check1_CheckInst_2_U89  ( .A1(\Check1_CheckInst_2_n84 ), .A2(
        \Check1_CheckInst_2_n83 ), .ZN(\Check1_CheckInst_2_n85 ) );
  NOR2_X1 \Check1_CheckInst_2_U88  ( .A1(\Check1_CheckInst_2_n82 ), .A2(
        \Check1_CheckInst_2_n81 ), .ZN(\Check1_CheckInst_2_n83 ) );
  XOR2_X1 \Check1_CheckInst_2_U87  ( .A(Red_AddRoundKeyOutput3[14]), .B(
        Red_SignaltoCheck[14]), .Z(\Check1_CheckInst_2_n81 ) );
  XOR2_X1 \Check1_CheckInst_2_U86  ( .A(Red_SignaltoCheck[6]), .B(
        Red_AddRoundKeyOutput3[6]), .Z(\Check1_CheckInst_2_n82 ) );
  NOR2_X1 \Check1_CheckInst_2_U85  ( .A1(\Check1_CheckInst_2_n80 ), .A2(
        \Check1_CheckInst_2_n79 ), .ZN(\Check1_CheckInst_2_n84 ) );
  XOR2_X1 \Check1_CheckInst_2_U84  ( .A(Red_AddRoundKeyOutput3[22]), .B(
        Red_SignaltoCheck[22]), .Z(\Check1_CheckInst_2_n79 ) );
  XOR2_X1 \Check1_CheckInst_2_U83  ( .A(Red_AddRoundKeyOutput3[18]), .B(
        Red_SignaltoCheck[18]), .Z(\Check1_CheckInst_2_n80 ) );
  NAND2_X1 \Check1_CheckInst_2_U82  ( .A1(\Check1_CheckInst_2_n78 ), .A2(
        \Check1_CheckInst_2_n77 ), .ZN(\Check1_CheckInst_2_n86 ) );
  XNOR2_X1 \Check1_CheckInst_2_U81  ( .A(Red_AddRoundKeyOutput[62]), .B(
        Red_SignaltoCheck[190]), .ZN(\Check1_CheckInst_2_n77 ) );
  XNOR2_X1 \Check1_CheckInst_2_U80  ( .A(Red_AddRoundKeyOutput[58]), .B(
        Red_SignaltoCheck[186]), .ZN(\Check1_CheckInst_2_n78 ) );
  NOR2_X1 \Check1_CheckInst_2_U79  ( .A1(\Check1_CheckInst_2_n76 ), .A2(
        \Check1_CheckInst_2_n75 ), .ZN(\Check1_CheckInst_2_n88 ) );
  XOR2_X1 \Check1_CheckInst_2_U78  ( .A(Red_AddRoundKeyOutput[46]), .B(
        Red_SignaltoCheck[174]), .Z(\Check1_CheckInst_2_n75 ) );
  XOR2_X1 \Check1_CheckInst_2_U77  ( .A(Red_AddRoundKeyOutput[54]), .B(
        Red_SignaltoCheck[182]), .Z(\Check1_CheckInst_2_n76 ) );
  NAND2_X1 \Check1_CheckInst_2_U76  ( .A1(\Check1_CheckInst_2_n74 ), .A2(
        \Check1_CheckInst_2_n73 ), .ZN(\Check1_CheckInst_2_n90 ) );
  NOR2_X1 \Check1_CheckInst_2_U75  ( .A1(\Check1_CheckInst_2_n72 ), .A2(
        \Check1_CheckInst_2_n71 ), .ZN(\Check1_CheckInst_2_n73 ) );
  NAND2_X1 \Check1_CheckInst_2_U74  ( .A1(\Check1_CheckInst_2_n70 ), .A2(
        \Check1_CheckInst_2_n69 ), .ZN(\Check1_CheckInst_2_n71 ) );
  NOR2_X1 \Check1_CheckInst_2_U73  ( .A1(\Check1_CheckInst_2_n68 ), .A2(
        \Check1_CheckInst_2_n67 ), .ZN(\Check1_CheckInst_2_n69 ) );
  XOR2_X1 \Check1_CheckInst_2_U72  ( .A(Red_AddRoundKeyOutput[38]), .B(
        Red_SignaltoCheck[166]), .Z(\Check1_CheckInst_2_n67 ) );
  XOR2_X1 \Check1_CheckInst_2_U71  ( .A(Red_AddRoundKeyOutput[50]), .B(
        Red_SignaltoCheck[178]), .Z(\Check1_CheckInst_2_n68 ) );
  NOR2_X1 \Check1_CheckInst_2_U70  ( .A1(\Check1_CheckInst_2_n66 ), .A2(
        \Check1_CheckInst_2_n65 ), .ZN(\Check1_CheckInst_2_n70 ) );
  XOR2_X1 \Check1_CheckInst_2_U69  ( .A(Red_Feedback3[22]), .B(
        Red_SignaltoCheck[214]), .Z(\Check1_CheckInst_2_n65 ) );
  XOR2_X1 \Check1_CheckInst_2_U68  ( .A(Red_AddRoundKeyOutput[42]), .B(
        Red_SignaltoCheck[170]), .Z(\Check1_CheckInst_2_n66 ) );
  NAND2_X1 \Check1_CheckInst_2_U67  ( .A1(\Check1_CheckInst_2_n64 ), .A2(
        \Check1_CheckInst_2_n63 ), .ZN(\Check1_CheckInst_2_n72 ) );
  XNOR2_X1 \Check1_CheckInst_2_U66  ( .A(Red_Feedback3[18]), .B(
        Red_SignaltoCheck[210]), .ZN(\Check1_CheckInst_2_n63 ) );
  XNOR2_X1 \Check1_CheckInst_2_U65  ( .A(Red_Feedback3[26]), .B(
        Red_SignaltoCheck[218]), .ZN(\Check1_CheckInst_2_n64 ) );
  NOR2_X1 \Check1_CheckInst_2_U64  ( .A1(\Check1_CheckInst_2_n62 ), .A2(
        \Check1_CheckInst_2_n61 ), .ZN(\Check1_CheckInst_2_n74 ) );
  XOR2_X1 \Check1_CheckInst_2_U63  ( .A(Red_Feedback3[14]), .B(
        Red_SignaltoCheck[206]), .Z(\Check1_CheckInst_2_n61 ) );
  XOR2_X1 \Check1_CheckInst_2_U62  ( .A(Red_Feedback3[10]), .B(
        Red_SignaltoCheck[202]), .Z(\Check1_CheckInst_2_n62 ) );
  NOR2_X1 \Check1_CheckInst_2_U61  ( .A1(\Check1_CheckInst_2_n60 ), .A2(
        \Check1_CheckInst_2_n59 ), .ZN(\Check1_CheckInst_2_n92 ) );
  NAND2_X1 \Check1_CheckInst_2_U60  ( .A1(\Check1_CheckInst_2_n58 ), .A2(
        \Check1_CheckInst_2_n57 ), .ZN(\Check1_CheckInst_2_n59 ) );
  NOR2_X1 \Check1_CheckInst_2_U59  ( .A1(\Check1_CheckInst_2_n56 ), .A2(
        \Check1_CheckInst_2_n55 ), .ZN(\Check1_CheckInst_2_n57 ) );
  NAND2_X1 \Check1_CheckInst_2_U58  ( .A1(\Check1_CheckInst_2_n54 ), .A2(
        \Check1_CheckInst_2_n53 ), .ZN(\Check1_CheckInst_2_n55 ) );
  XNOR2_X1 \Check1_CheckInst_2_U57  ( .A(Red_Feedback3[6]), .B(
        Red_SignaltoCheck[198]), .ZN(\Check1_CheckInst_2_n53 ) );
  XNOR2_X1 \Check1_CheckInst_2_U56  ( .A(Red_Feedback3[2]), .B(
        Red_SignaltoCheck[194]), .ZN(\Check1_CheckInst_2_n54 ) );
  NAND2_X1 \Check1_CheckInst_2_U55  ( .A1(\Check1_CheckInst_2_n52 ), .A2(
        \Check1_CheckInst_2_n51 ), .ZN(\Check1_CheckInst_2_n56 ) );
  XNOR2_X1 \Check1_CheckInst_2_U54  ( .A(Red_AddRoundKeyOutput[6]), .B(
        Red_SignaltoCheck[134]), .ZN(\Check1_CheckInst_2_n51 ) );
  XNOR2_X1 \Check1_CheckInst_2_U53  ( .A(Red_AddRoundKeyOutput[2]), .B(
        Red_SignaltoCheck[130]), .ZN(\Check1_CheckInst_2_n52 ) );
  NOR2_X1 \Check1_CheckInst_2_U52  ( .A1(\Check1_CheckInst_2_n50 ), .A2(
        \Check1_CheckInst_2_n49 ), .ZN(\Check1_CheckInst_2_n58 ) );
  XOR2_X1 \Check1_CheckInst_2_U51  ( .A(Red_AddRoundKeyOutput2[54]), .B(
        Red_SignaltoCheck[118]), .Z(\Check1_CheckInst_2_n49 ) );
  XOR2_X1 \Check1_CheckInst_2_U50  ( .A(Red_AddRoundKeyOutput2[62]), .B(
        Red_SignaltoCheck[126]), .Z(\Check1_CheckInst_2_n50 ) );
  NAND2_X1 \Check1_CheckInst_2_U49  ( .A1(\Check1_CheckInst_2_n48 ), .A2(
        \Check1_CheckInst_2_n47 ), .ZN(\Check1_CheckInst_2_n60 ) );
  XNOR2_X1 \Check1_CheckInst_2_U48  ( .A(Red_AddRoundKeyOutput2[46]), .B(
        Red_SignaltoCheck[110]), .ZN(\Check1_CheckInst_2_n47 ) );
  XNOR2_X1 \Check1_CheckInst_2_U47  ( .A(Red_AddRoundKeyOutput2[58]), .B(
        Red_SignaltoCheck[122]), .ZN(\Check1_CheckInst_2_n48 ) );
  NAND2_X1 \Check1_CheckInst_2_U46  ( .A1(\Check1_CheckInst_2_n46 ), .A2(
        \Check1_CheckInst_2_n45 ), .ZN(\Check1_CheckInst_2_n94 ) );
  NOR2_X1 \Check1_CheckInst_2_U45  ( .A1(\Check1_CheckInst_2_n44 ), .A2(
        \Check1_CheckInst_2_n43 ), .ZN(\Check1_CheckInst_2_n45 ) );
  NAND2_X1 \Check1_CheckInst_2_U44  ( .A1(\Check1_CheckInst_2_n42 ), .A2(
        \Check1_CheckInst_2_n41 ), .ZN(\Check1_CheckInst_2_n43 ) );
  NOR2_X1 \Check1_CheckInst_2_U43  ( .A1(\Check1_CheckInst_2_n40 ), .A2(
        \Check1_CheckInst_2_n39 ), .ZN(\Check1_CheckInst_2_n41 ) );
  XOR2_X1 \Check1_CheckInst_2_U42  ( .A(Red_AddRoundKeyOutput[30]), .B(
        Red_SignaltoCheck[158]), .Z(\Check1_CheckInst_2_n39 ) );
  XOR2_X1 \Check1_CheckInst_2_U41  ( .A(Red_AddRoundKeyOutput2[50]), .B(
        Red_SignaltoCheck[114]), .Z(\Check1_CheckInst_2_n40 ) );
  NOR2_X1 \Check1_CheckInst_2_U40  ( .A1(\Check1_CheckInst_2_n38 ), .A2(
        \Check1_CheckInst_2_n37 ), .ZN(\Check1_CheckInst_2_n42 ) );
  XOR2_X1 \Check1_CheckInst_2_U39  ( .A(Red_AddRoundKeyOutput[26]), .B(
        Red_SignaltoCheck[154]), .Z(\Check1_CheckInst_2_n37 ) );
  XOR2_X1 \Check1_CheckInst_2_U38  ( .A(Red_AddRoundKeyOutput[34]), .B(
        Red_SignaltoCheck[162]), .Z(\Check1_CheckInst_2_n38 ) );
  NAND2_X1 \Check1_CheckInst_2_U37  ( .A1(\Check1_CheckInst_2_n36 ), .A2(
        \Check1_CheckInst_2_n35 ), .ZN(\Check1_CheckInst_2_n44 ) );
  XNOR2_X1 \Check1_CheckInst_2_U36  ( .A(Red_AddRoundKeyOutput[22]), .B(
        Red_SignaltoCheck[150]), .ZN(\Check1_CheckInst_2_n35 ) );
  XNOR2_X1 \Check1_CheckInst_2_U35  ( .A(Red_AddRoundKeyOutput[18]), .B(
        Red_SignaltoCheck[146]), .ZN(\Check1_CheckInst_2_n36 ) );
  NOR2_X1 \Check1_CheckInst_2_U34  ( .A1(\Check1_CheckInst_2_n34 ), .A2(
        \Check1_CheckInst_2_n33 ), .ZN(\Check1_CheckInst_2_n46 ) );
  XOR2_X1 \Check1_CheckInst_2_U33  ( .A(Red_AddRoundKeyOutput[14]), .B(
        Red_SignaltoCheck[142]), .Z(\Check1_CheckInst_2_n33 ) );
  XOR2_X1 \Check1_CheckInst_2_U32  ( .A(Red_AddRoundKeyOutput[10]), .B(
        Red_SignaltoCheck[138]), .Z(\Check1_CheckInst_2_n34 ) );
  NAND2_X1 \Check1_CheckInst_2_U31  ( .A1(\Check1_CheckInst_2_n32 ), .A2(
        \Check1_CheckInst_2_n31 ), .ZN(\Check1_CheckInst_2_n224 ) );
  NOR2_X1 \Check1_CheckInst_2_U30  ( .A1(\Check1_CheckInst_2_n30 ), .A2(
        \Check1_CheckInst_2_n29 ), .ZN(\Check1_CheckInst_2_n31 ) );
  NAND2_X1 \Check1_CheckInst_2_U29  ( .A1(\Check1_CheckInst_2_n28 ), .A2(
        \Check1_CheckInst_2_n27 ), .ZN(\Check1_CheckInst_2_n29 ) );
  NOR2_X1 \Check1_CheckInst_2_U28  ( .A1(\Check1_CheckInst_2_n26 ), .A2(
        \Check1_CheckInst_2_n25 ), .ZN(\Check1_CheckInst_2_n27 ) );
  NAND2_X1 \Check1_CheckInst_2_U27  ( .A1(\Check1_CheckInst_2_n24 ), .A2(
        \Check1_CheckInst_2_n23 ), .ZN(\Check1_CheckInst_2_n25 ) );
  XNOR2_X1 \Check1_CheckInst_2_U26  ( .A(Red_StateRegOutput3[30]), .B(
        Red_SignaltoCheck[286]), .ZN(\Check1_CheckInst_2_n23 ) );
  XNOR2_X1 \Check1_CheckInst_2_U25  ( .A(Red_StateRegOutput3[38]), .B(
        Red_SignaltoCheck[294]), .ZN(\Check1_CheckInst_2_n24 ) );
  NAND2_X1 \Check1_CheckInst_2_U24  ( .A1(\Check1_CheckInst_2_n22 ), .A2(
        \Check1_CheckInst_2_n21 ), .ZN(\Check1_CheckInst_2_n26 ) );
  XNOR2_X1 \Check1_CheckInst_2_U23  ( .A(Red_StateRegOutput3[46]), .B(
        Red_SignaltoCheck[302]), .ZN(\Check1_CheckInst_2_n21 ) );
  XNOR2_X1 \Check1_CheckInst_2_U22  ( .A(Red_StateRegOutput3[42]), .B(
        Red_SignaltoCheck[298]), .ZN(\Check1_CheckInst_2_n22 ) );
  NOR2_X1 \Check1_CheckInst_2_U21  ( .A1(\Check1_CheckInst_2_n20 ), .A2(
        \Check1_CheckInst_2_n19 ), .ZN(\Check1_CheckInst_2_n28 ) );
  NAND2_X1 \Check1_CheckInst_2_U20  ( .A1(\Check1_CheckInst_2_n18 ), .A2(
        \Check1_CheckInst_2_n17 ), .ZN(\Check1_CheckInst_2_n19 ) );
  XNOR2_X1 \Check1_CheckInst_2_U19  ( .A(Red_StateRegOutput2[6]), .B(
        Red_SignaltoCheck[326]), .ZN(\Check1_CheckInst_2_n17 ) );
  XNOR2_X1 \Check1_CheckInst_2_U18  ( .A(Red_StateRegOutput3[26]), .B(
        Red_SignaltoCheck[282]), .ZN(\Check1_CheckInst_2_n18 ) );
  NAND2_X1 \Check1_CheckInst_2_U17  ( .A1(\Check1_CheckInst_2_n16 ), .A2(
        \Check1_CheckInst_2_n15 ), .ZN(\Check1_CheckInst_2_n20 ) );
  XNOR2_X1 \Check1_CheckInst_2_U16  ( .A(Red_StateRegOutput3[22]), .B(
        Red_SignaltoCheck[278]), .ZN(\Check1_CheckInst_2_n15 ) );
  XNOR2_X1 \Check1_CheckInst_2_U15  ( .A(Red_StateRegOutput3[34]), .B(
        Red_SignaltoCheck[290]), .ZN(\Check1_CheckInst_2_n16 ) );
  NAND2_X1 \Check1_CheckInst_2_U14  ( .A1(\Check1_CheckInst_2_n14 ), .A2(
        \Check1_CheckInst_2_n13 ), .ZN(\Check1_CheckInst_2_n30 ) );
  NOR2_X1 \Check1_CheckInst_2_U13  ( .A1(\Check1_CheckInst_2_n12 ), .A2(
        \Check1_CheckInst_2_n11 ), .ZN(\Check1_CheckInst_2_n13 ) );
  XOR2_X1 \Check1_CheckInst_2_U12  ( .A(Red_StateRegOutput3[62]), .B(
        Red_SignaltoCheck[318]), .Z(\Check1_CheckInst_2_n11 ) );
  XOR2_X1 \Check1_CheckInst_2_U11  ( .A(Red_StateRegOutput3[58]), .B(
        Red_SignaltoCheck[314]), .Z(\Check1_CheckInst_2_n12 ) );
  NOR2_X1 \Check1_CheckInst_2_U10  ( .A1(\Check1_CheckInst_2_n10 ), .A2(
        \Check1_CheckInst_2_n9 ), .ZN(\Check1_CheckInst_2_n14 ) );
  XOR2_X1 \Check1_CheckInst_2_U9  ( .A(Red_StateRegOutput2[2]), .B(
        Red_SignaltoCheck[322]), .Z(\Check1_CheckInst_2_n9 ) );
  XOR2_X1 \Check1_CheckInst_2_U8  ( .A(Red_StateRegOutput2[10]), .B(
        Red_SignaltoCheck[330]), .Z(\Check1_CheckInst_2_n10 ) );
  NOR2_X1 \Check1_CheckInst_2_U7  ( .A1(\Check1_CheckInst_2_n8 ), .A2(
        \Check1_CheckInst_2_n7 ), .ZN(\Check1_CheckInst_2_n32 ) );
  NAND2_X1 \Check1_CheckInst_2_U6  ( .A1(\Check1_CheckInst_2_n6 ), .A2(
        \Check1_CheckInst_2_n5 ), .ZN(\Check1_CheckInst_2_n7 ) );
  XNOR2_X1 \Check1_CheckInst_2_U5  ( .A(Red_Feedback3[54]), .B(
        Red_SignaltoCheck[246]), .ZN(\Check1_CheckInst_2_n5 ) );
  XNOR2_X1 \Check1_CheckInst_2_U4  ( .A(Red_Feedback3[50]), .B(
        Red_SignaltoCheck[242]), .ZN(\Check1_CheckInst_2_n6 ) );
  NAND2_X1 \Check1_CheckInst_2_U3  ( .A1(\Check1_CheckInst_2_n4 ), .A2(
        \Check1_CheckInst_2_n3 ), .ZN(\Check1_CheckInst_2_n8 ) );
  XNOR2_X1 \Check1_CheckInst_2_U2  ( .A(Red_StateRegOutput3[54]), .B(
        Red_SignaltoCheck[310]), .ZN(\Check1_CheckInst_2_n3 ) );
  XNOR2_X1 \Check1_CheckInst_2_U1  ( .A(Red_StateRegOutput3[50]), .B(
        Red_SignaltoCheck[306]), .ZN(\Check1_CheckInst_2_n4 ) );
  NOR2_X1 \Check1_CheckInst_3_U223  ( .A1(\Check1_CheckInst_3_n224 ), .A2(
        \Check1_CheckInst_3_n223 ), .ZN(Error[3]) );
  NAND2_X1 \Check1_CheckInst_3_U222  ( .A1(\Check1_CheckInst_3_n222 ), .A2(
        \Check1_CheckInst_3_n221 ), .ZN(\Check1_CheckInst_3_n223 ) );
  NOR2_X1 \Check1_CheckInst_3_U221  ( .A1(\Check1_CheckInst_3_n220 ), .A2(
        \Check1_CheckInst_3_n219 ), .ZN(\Check1_CheckInst_3_n221 ) );
  NAND2_X1 \Check1_CheckInst_3_U220  ( .A1(\Check1_CheckInst_3_n218 ), .A2(
        \Check1_CheckInst_3_n217 ), .ZN(\Check1_CheckInst_3_n219 ) );
  NOR2_X1 \Check1_CheckInst_3_U219  ( .A1(\Check1_CheckInst_3_n216 ), .A2(
        \Check1_CheckInst_3_n215 ), .ZN(\Check1_CheckInst_3_n217 ) );
  NAND2_X1 \Check1_CheckInst_3_U218  ( .A1(\Check1_CheckInst_3_n214 ), .A2(
        \Check1_CheckInst_3_n213 ), .ZN(\Check1_CheckInst_3_n215 ) );
  NOR2_X1 \Check1_CheckInst_3_U217  ( .A1(\Check1_CheckInst_3_n212 ), .A2(
        \Check1_CheckInst_3_n211 ), .ZN(\Check1_CheckInst_3_n213 ) );
  NAND2_X1 \Check1_CheckInst_3_U216  ( .A1(\Check1_CheckInst_3_n210 ), .A2(
        \Check1_CheckInst_3_n209 ), .ZN(\Check1_CheckInst_3_n211 ) );
  NOR2_X1 \Check1_CheckInst_3_U215  ( .A1(\Check1_CheckInst_3_n208 ), .A2(
        \Check1_CheckInst_3_n207 ), .ZN(\Check1_CheckInst_3_n209 ) );
  NAND2_X1 \Check1_CheckInst_3_U214  ( .A1(\Check1_CheckInst_3_n206 ), .A2(
        \Check1_CheckInst_3_n205 ), .ZN(\Check1_CheckInst_3_n207 ) );
  XNOR2_X1 \Check1_CheckInst_3_U213  ( .A(Red_Feedback3[39]), .B(
        Red_SignaltoCheck[231]), .ZN(\Check1_CheckInst_3_n205 ) );
  XNOR2_X1 \Check1_CheckInst_3_U212  ( .A(Red_Feedback3[47]), .B(
        Red_SignaltoCheck[239]), .ZN(\Check1_CheckInst_3_n206 ) );
  NAND2_X1 \Check1_CheckInst_3_U211  ( .A1(\Check1_CheckInst_3_n204 ), .A2(
        \Check1_CheckInst_3_n203 ), .ZN(\Check1_CheckInst_3_n208 ) );
  XNOR2_X1 \Check1_CheckInst_3_U210  ( .A(Red_Feedback3[31]), .B(
        Red_SignaltoCheck[223]), .ZN(\Check1_CheckInst_3_n203 ) );
  XNOR2_X1 \Check1_CheckInst_3_U209  ( .A(Red_Feedback3[43]), .B(
        Red_SignaltoCheck[235]), .ZN(\Check1_CheckInst_3_n204 ) );
  NOR2_X1 \Check1_CheckInst_3_U208  ( .A1(\Check1_CheckInst_3_n202 ), .A2(
        \Check1_CheckInst_3_n201 ), .ZN(\Check1_CheckInst_3_n210 ) );
  XOR2_X1 \Check1_CheckInst_3_U207  ( .A(Red_StateRegOutput3[15]), .B(
        Red_SignaltoCheck[271]), .Z(\Check1_CheckInst_3_n201 ) );
  XOR2_X1 \Check1_CheckInst_3_U206  ( .A(Red_Feedback3[35]), .B(
        Red_SignaltoCheck[227]), .Z(\Check1_CheckInst_3_n202 ) );
  NAND2_X1 \Check1_CheckInst_3_U205  ( .A1(\Check1_CheckInst_3_n200 ), .A2(
        \Check1_CheckInst_3_n199 ), .ZN(\Check1_CheckInst_3_n212 ) );
  XNOR2_X1 \Check1_CheckInst_3_U204  ( .A(Red_StateRegOutput3[11]), .B(
        Red_SignaltoCheck[267]), .ZN(\Check1_CheckInst_3_n199 ) );
  XNOR2_X1 \Check1_CheckInst_3_U203  ( .A(Red_StateRegOutput3[19]), .B(
        Red_SignaltoCheck[275]), .ZN(\Check1_CheckInst_3_n200 ) );
  NOR2_X1 \Check1_CheckInst_3_U202  ( .A1(\Check1_CheckInst_3_n198 ), .A2(
        \Check1_CheckInst_3_n197 ), .ZN(\Check1_CheckInst_3_n214 ) );
  NAND2_X1 \Check1_CheckInst_3_U201  ( .A1(\Check1_CheckInst_3_n196 ), .A2(
        \Check1_CheckInst_3_n195 ), .ZN(\Check1_CheckInst_3_n197 ) );
  NOR2_X1 \Check1_CheckInst_3_U200  ( .A1(\Check1_CheckInst_3_n194 ), .A2(
        \Check1_CheckInst_3_n193 ), .ZN(\Check1_CheckInst_3_n195 ) );
  NAND2_X1 \Check1_CheckInst_3_U199  ( .A1(\Check1_CheckInst_3_n192 ), .A2(
        \Check1_CheckInst_3_n191 ), .ZN(\Check1_CheckInst_3_n193 ) );
  XNOR2_X1 \Check1_CheckInst_3_U198  ( .A(Red_StateRegOutput3[7]), .B(
        Red_SignaltoCheck[263]), .ZN(\Check1_CheckInst_3_n191 ) );
  XNOR2_X1 \Check1_CheckInst_3_U197  ( .A(Red_StateRegOutput3[3]), .B(
        Red_SignaltoCheck[259]), .ZN(\Check1_CheckInst_3_n192 ) );
  NAND2_X1 \Check1_CheckInst_3_U196  ( .A1(\Check1_CheckInst_3_n190 ), .A2(
        \Check1_CheckInst_3_n189 ), .ZN(\Check1_CheckInst_3_n194 ) );
  XNOR2_X1 \Check1_CheckInst_3_U195  ( .A(Red_Feedback3[63]), .B(
        Red_SignaltoCheck[255]), .ZN(\Check1_CheckInst_3_n189 ) );
  XNOR2_X1 \Check1_CheckInst_3_U194  ( .A(Red_Feedback3[59]), .B(
        Red_SignaltoCheck[251]), .ZN(\Check1_CheckInst_3_n190 ) );
  NOR2_X1 \Check1_CheckInst_3_U193  ( .A1(\Check1_CheckInst_3_n188 ), .A2(
        \Check1_CheckInst_3_n187 ), .ZN(\Check1_CheckInst_3_n196 ) );
  XOR2_X1 \Check1_CheckInst_3_U192  ( .A(Red_StateRegOutput[31]), .B(
        Red_SignaltoCheck[415]), .Z(\Check1_CheckInst_3_n187 ) );
  XOR2_X1 \Check1_CheckInst_3_U191  ( .A(Red_StateRegOutput[27]), .B(
        Red_SignaltoCheck[411]), .Z(\Check1_CheckInst_3_n188 ) );
  NAND2_X1 \Check1_CheckInst_3_U190  ( .A1(\Check1_CheckInst_3_n186 ), .A2(
        \Check1_CheckInst_3_n185 ), .ZN(\Check1_CheckInst_3_n198 ) );
  XNOR2_X1 \Check1_CheckInst_3_U189  ( .A(Red_StateRegOutput[15]), .B(
        Red_SignaltoCheck[399]), .ZN(\Check1_CheckInst_3_n185 ) );
  XNOR2_X1 \Check1_CheckInst_3_U188  ( .A(Red_StateRegOutput[23]), .B(
        Red_SignaltoCheck[407]), .ZN(\Check1_CheckInst_3_n186 ) );
  NAND2_X1 \Check1_CheckInst_3_U187  ( .A1(\Check1_CheckInst_3_n184 ), .A2(
        \Check1_CheckInst_3_n183 ), .ZN(\Check1_CheckInst_3_n216 ) );
  NOR2_X1 \Check1_CheckInst_3_U186  ( .A1(\Check1_CheckInst_3_n182 ), .A2(
        \Check1_CheckInst_3_n181 ), .ZN(\Check1_CheckInst_3_n183 ) );
  NAND2_X1 \Check1_CheckInst_3_U185  ( .A1(\Check1_CheckInst_3_n180 ), .A2(
        \Check1_CheckInst_3_n179 ), .ZN(\Check1_CheckInst_3_n181 ) );
  NOR2_X1 \Check1_CheckInst_3_U184  ( .A1(\Check1_CheckInst_3_n178 ), .A2(
        \Check1_CheckInst_3_n177 ), .ZN(\Check1_CheckInst_3_n179 ) );
  XOR2_X1 \Check1_CheckInst_3_U183  ( .A(Red_StateRegOutput[7]), .B(
        Red_SignaltoCheck[391]), .Z(\Check1_CheckInst_3_n177 ) );
  XOR2_X1 \Check1_CheckInst_3_U182  ( .A(Red_StateRegOutput[19]), .B(
        Red_SignaltoCheck[403]), .Z(\Check1_CheckInst_3_n178 ) );
  NOR2_X1 \Check1_CheckInst_3_U181  ( .A1(\Check1_CheckInst_3_n176 ), .A2(
        \Check1_CheckInst_3_n175 ), .ZN(\Check1_CheckInst_3_n180 ) );
  XOR2_X1 \Check1_CheckInst_3_U180  ( .A(Red_StateRegOutput[55]), .B(
        Red_SignaltoCheck[439]), .Z(\Check1_CheckInst_3_n175 ) );
  XOR2_X1 \Check1_CheckInst_3_U179  ( .A(Red_StateRegOutput[11]), .B(
        Red_SignaltoCheck[395]), .Z(\Check1_CheckInst_3_n176 ) );
  NAND2_X1 \Check1_CheckInst_3_U178  ( .A1(\Check1_CheckInst_3_n174 ), .A2(
        \Check1_CheckInst_3_n173 ), .ZN(\Check1_CheckInst_3_n182 ) );
  XNOR2_X1 \Check1_CheckInst_3_U177  ( .A(Red_StateRegOutput[51]), .B(
        Red_SignaltoCheck[435]), .ZN(\Check1_CheckInst_3_n173 ) );
  XNOR2_X1 \Check1_CheckInst_3_U176  ( .A(Red_StateRegOutput[59]), .B(
        Red_SignaltoCheck[443]), .ZN(\Check1_CheckInst_3_n174 ) );
  NOR2_X1 \Check1_CheckInst_3_U175  ( .A1(\Check1_CheckInst_3_n172 ), .A2(
        \Check1_CheckInst_3_n171 ), .ZN(\Check1_CheckInst_3_n184 ) );
  XOR2_X1 \Check1_CheckInst_3_U174  ( .A(Red_StateRegOutput[47]), .B(
        Red_SignaltoCheck[431]), .Z(\Check1_CheckInst_3_n171 ) );
  XOR2_X1 \Check1_CheckInst_3_U173  ( .A(Red_StateRegOutput[43]), .B(
        Red_SignaltoCheck[427]), .Z(\Check1_CheckInst_3_n172 ) );
  NOR2_X1 \Check1_CheckInst_3_U172  ( .A1(\Check1_CheckInst_3_n170 ), .A2(
        \Check1_CheckInst_3_n169 ), .ZN(\Check1_CheckInst_3_n218 ) );
  NAND2_X1 \Check1_CheckInst_3_U171  ( .A1(\Check1_CheckInst_3_n168 ), .A2(
        \Check1_CheckInst_3_n167 ), .ZN(\Check1_CheckInst_3_n169 ) );
  NOR2_X1 \Check1_CheckInst_3_U170  ( .A1(\Check1_CheckInst_3_n166 ), .A2(
        \Check1_CheckInst_3_n165 ), .ZN(\Check1_CheckInst_3_n167 ) );
  NAND2_X1 \Check1_CheckInst_3_U169  ( .A1(\Check1_CheckInst_3_n164 ), .A2(
        \Check1_CheckInst_3_n163 ), .ZN(\Check1_CheckInst_3_n165 ) );
  XNOR2_X1 \Check1_CheckInst_3_U168  ( .A(Red_StateRegOutput[39]), .B(
        Red_SignaltoCheck[423]), .ZN(\Check1_CheckInst_3_n163 ) );
  XNOR2_X1 \Check1_CheckInst_3_U167  ( .A(Red_StateRegOutput[35]), .B(
        Red_SignaltoCheck[419]), .ZN(\Check1_CheckInst_3_n164 ) );
  NAND2_X1 \Check1_CheckInst_3_U166  ( .A1(\Check1_CheckInst_3_n162 ), .A2(
        \Check1_CheckInst_3_n161 ), .ZN(\Check1_CheckInst_3_n166 ) );
  XNOR2_X1 \Check1_CheckInst_3_U165  ( .A(Red_StateRegOutput2[39]), .B(
        Red_SignaltoCheck[359]), .ZN(\Check1_CheckInst_3_n161 ) );
  XNOR2_X1 \Check1_CheckInst_3_U164  ( .A(Red_StateRegOutput2[35]), .B(
        Red_SignaltoCheck[355]), .ZN(\Check1_CheckInst_3_n162 ) );
  NOR2_X1 \Check1_CheckInst_3_U163  ( .A1(\Check1_CheckInst_3_n160 ), .A2(
        \Check1_CheckInst_3_n159 ), .ZN(\Check1_CheckInst_3_n168 ) );
  XOR2_X1 \Check1_CheckInst_3_U162  ( .A(Red_StateRegOutput2[23]), .B(
        Red_SignaltoCheck[343]), .Z(\Check1_CheckInst_3_n159 ) );
  XOR2_X1 \Check1_CheckInst_3_U161  ( .A(Red_StateRegOutput2[31]), .B(
        Red_SignaltoCheck[351]), .Z(\Check1_CheckInst_3_n160 ) );
  NAND2_X1 \Check1_CheckInst_3_U160  ( .A1(\Check1_CheckInst_3_n158 ), .A2(
        \Check1_CheckInst_3_n157 ), .ZN(\Check1_CheckInst_3_n170 ) );
  XNOR2_X1 \Check1_CheckInst_3_U159  ( .A(Red_StateRegOutput2[15]), .B(
        Red_SignaltoCheck[335]), .ZN(\Check1_CheckInst_3_n157 ) );
  XNOR2_X1 \Check1_CheckInst_3_U158  ( .A(Red_StateRegOutput2[27]), .B(
        Red_SignaltoCheck[347]), .ZN(\Check1_CheckInst_3_n158 ) );
  NAND2_X1 \Check1_CheckInst_3_U157  ( .A1(\Check1_CheckInst_3_n156 ), .A2(
        \Check1_CheckInst_3_n155 ), .ZN(\Check1_CheckInst_3_n220 ) );
  NOR2_X1 \Check1_CheckInst_3_U156  ( .A1(\Check1_CheckInst_3_n154 ), .A2(
        \Check1_CheckInst_3_n153 ), .ZN(\Check1_CheckInst_3_n155 ) );
  NAND2_X1 \Check1_CheckInst_3_U155  ( .A1(\Check1_CheckInst_3_n152 ), .A2(
        \Check1_CheckInst_3_n151 ), .ZN(\Check1_CheckInst_3_n153 ) );
  NOR2_X1 \Check1_CheckInst_3_U154  ( .A1(\Check1_CheckInst_3_n150 ), .A2(
        \Check1_CheckInst_3_n149 ), .ZN(\Check1_CheckInst_3_n151 ) );
  NAND2_X1 \Check1_CheckInst_3_U153  ( .A1(\Check1_CheckInst_3_n148 ), .A2(
        \Check1_CheckInst_3_n147 ), .ZN(\Check1_CheckInst_3_n149 ) );
  NOR2_X1 \Check1_CheckInst_3_U152  ( .A1(\Check1_CheckInst_3_n146 ), .A2(
        \Check1_CheckInst_3_n145 ), .ZN(\Check1_CheckInst_3_n147 ) );
  NAND2_X1 \Check1_CheckInst_3_U151  ( .A1(\Check1_CheckInst_3_n144 ), .A2(
        \Check1_CheckInst_3_n143 ), .ZN(\Check1_CheckInst_3_n145 ) );
  XNOR2_X1 \Check1_CheckInst_3_U150  ( .A(Red_StateRegOutput2[63]), .B(
        Red_SignaltoCheck[383]), .ZN(\Check1_CheckInst_3_n143 ) );
  XNOR2_X1 \Check1_CheckInst_3_U149  ( .A(Red_StateRegOutput2[19]), .B(
        Red_SignaltoCheck[339]), .ZN(\Check1_CheckInst_3_n144 ) );
  NAND2_X1 \Check1_CheckInst_3_U148  ( .A1(\Check1_CheckInst_3_n142 ), .A2(
        \Check1_CheckInst_3_n141 ), .ZN(\Check1_CheckInst_3_n146 ) );
  XNOR2_X1 \Check1_CheckInst_3_U147  ( .A(Red_StateRegOutput2[59]), .B(
        Red_SignaltoCheck[379]), .ZN(\Check1_CheckInst_3_n141 ) );
  XNOR2_X1 \Check1_CheckInst_3_U146  ( .A(Red_StateRegOutput[3]), .B(
        Red_SignaltoCheck[387]), .ZN(\Check1_CheckInst_3_n142 ) );
  NOR2_X1 \Check1_CheckInst_3_U145  ( .A1(\Check1_CheckInst_3_n140 ), .A2(
        \Check1_CheckInst_3_n139 ), .ZN(\Check1_CheckInst_3_n148 ) );
  XOR2_X1 \Check1_CheckInst_3_U144  ( .A(Red_StateRegOutput2[55]), .B(
        Red_SignaltoCheck[375]), .Z(\Check1_CheckInst_3_n139 ) );
  XOR2_X1 \Check1_CheckInst_3_U143  ( .A(Red_StateRegOutput2[51]), .B(
        Red_SignaltoCheck[371]), .Z(\Check1_CheckInst_3_n140 ) );
  NAND2_X1 \Check1_CheckInst_3_U142  ( .A1(\Check1_CheckInst_3_n138 ), .A2(
        \Check1_CheckInst_3_n137 ), .ZN(\Check1_CheckInst_3_n150 ) );
  XNOR2_X1 \Check1_CheckInst_3_U141  ( .A(Red_StateRegOutput2[47]), .B(
        Red_SignaltoCheck[367]), .ZN(\Check1_CheckInst_3_n137 ) );
  XNOR2_X1 \Check1_CheckInst_3_U140  ( .A(Red_StateRegOutput2[43]), .B(
        Red_SignaltoCheck[363]), .ZN(\Check1_CheckInst_3_n138 ) );
  NOR2_X1 \Check1_CheckInst_3_U139  ( .A1(\Check1_CheckInst_3_n136 ), .A2(
        \Check1_CheckInst_3_n135 ), .ZN(\Check1_CheckInst_3_n152 ) );
  NAND2_X1 \Check1_CheckInst_3_U138  ( .A1(\Check1_CheckInst_3_n134 ), .A2(
        \Check1_CheckInst_3_n133 ), .ZN(\Check1_CheckInst_3_n135 ) );
  NOR2_X1 \Check1_CheckInst_3_U137  ( .A1(\Check1_CheckInst_3_n132 ), .A2(
        \Check1_CheckInst_3_n131 ), .ZN(\Check1_CheckInst_3_n133 ) );
  NAND2_X1 \Check1_CheckInst_3_U136  ( .A1(\Check1_CheckInst_3_n130 ), .A2(
        \Check1_CheckInst_3_n129 ), .ZN(\Check1_CheckInst_3_n131 ) );
  XNOR2_X1 \Check1_CheckInst_3_U135  ( .A(Red_AddRoundKeyOutput2[15]), .B(
        Red_SignaltoCheck[79]), .ZN(\Check1_CheckInst_3_n129 ) );
  XNOR2_X1 \Check1_CheckInst_3_U134  ( .A(Red_AddRoundKeyOutput2[11]), .B(
        Red_SignaltoCheck[75]), .ZN(\Check1_CheckInst_3_n130 ) );
  NAND2_X1 \Check1_CheckInst_3_U133  ( .A1(\Check1_CheckInst_3_n128 ), .A2(
        \Check1_CheckInst_3_n127 ), .ZN(\Check1_CheckInst_3_n132 ) );
  XNOR2_X1 \Check1_CheckInst_3_U132  ( .A(Red_AddRoundKeyOutput3[63]), .B(
        Red_SignaltoCheck[63]), .ZN(\Check1_CheckInst_3_n127 ) );
  XNOR2_X1 \Check1_CheckInst_3_U131  ( .A(Red_AddRoundKeyOutput2[7]), .B(
        Red_SignaltoCheck[71]), .ZN(\Check1_CheckInst_3_n128 ) );
  NOR2_X1 \Check1_CheckInst_3_U130  ( .A1(\Check1_CheckInst_3_n126 ), .A2(
        \Check1_CheckInst_3_n125 ), .ZN(\Check1_CheckInst_3_n134 ) );
  XOR2_X1 \Check1_CheckInst_3_U129  ( .A(Red_AddRoundKeyOutput3[55]), .B(
        Red_SignaltoCheck[55]), .Z(\Check1_CheckInst_3_n125 ) );
  XOR2_X1 \Check1_CheckInst_3_U128  ( .A(Red_AddRoundKeyOutput2[3]), .B(
        Red_SignaltoCheck[67]), .Z(\Check1_CheckInst_3_n126 ) );
  NAND2_X1 \Check1_CheckInst_3_U127  ( .A1(\Check1_CheckInst_3_n124 ), .A2(
        \Check1_CheckInst_3_n123 ), .ZN(\Check1_CheckInst_3_n136 ) );
  XNOR2_X1 \Check1_CheckInst_3_U126  ( .A(Red_AddRoundKeyOutput2[39]), .B(
        Red_SignaltoCheck[103]), .ZN(\Check1_CheckInst_3_n123 ) );
  XNOR2_X1 \Check1_CheckInst_3_U125  ( .A(Red_AddRoundKeyOutput3[59]), .B(
        Red_SignaltoCheck[59]), .ZN(\Check1_CheckInst_3_n124 ) );
  NAND2_X1 \Check1_CheckInst_3_U124  ( .A1(\Check1_CheckInst_3_n122 ), .A2(
        \Check1_CheckInst_3_n121 ), .ZN(\Check1_CheckInst_3_n154 ) );
  NOR2_X1 \Check1_CheckInst_3_U123  ( .A1(\Check1_CheckInst_3_n120 ), .A2(
        \Check1_CheckInst_3_n119 ), .ZN(\Check1_CheckInst_3_n121 ) );
  NAND2_X1 \Check1_CheckInst_3_U122  ( .A1(\Check1_CheckInst_3_n118 ), .A2(
        \Check1_CheckInst_3_n117 ), .ZN(\Check1_CheckInst_3_n119 ) );
  NOR2_X1 \Check1_CheckInst_3_U121  ( .A1(\Check1_CheckInst_3_n116 ), .A2(
        \Check1_CheckInst_3_n115 ), .ZN(\Check1_CheckInst_3_n117 ) );
  XOR2_X1 \Check1_CheckInst_3_U120  ( .A(Red_AddRoundKeyOutput2[35]), .B(
        Red_SignaltoCheck[99]), .Z(\Check1_CheckInst_3_n115 ) );
  XOR2_X1 \Check1_CheckInst_3_U119  ( .A(Red_AddRoundKeyOutput2[43]), .B(
        Red_SignaltoCheck[107]), .Z(\Check1_CheckInst_3_n116 ) );
  NOR2_X1 \Check1_CheckInst_3_U118  ( .A1(\Check1_CheckInst_3_n114 ), .A2(
        \Check1_CheckInst_3_n113 ), .ZN(\Check1_CheckInst_3_n118 ) );
  XOR2_X1 \Check1_CheckInst_3_U117  ( .A(Red_AddRoundKeyOutput2[31]), .B(
        Red_SignaltoCheck[95]), .Z(\Check1_CheckInst_3_n113 ) );
  XOR2_X1 \Check1_CheckInst_3_U116  ( .A(Red_AddRoundKeyOutput2[27]), .B(
        Red_SignaltoCheck[91]), .Z(\Check1_CheckInst_3_n114 ) );
  NAND2_X1 \Check1_CheckInst_3_U115  ( .A1(\Check1_CheckInst_3_n112 ), .A2(
        \Check1_CheckInst_3_n111 ), .ZN(\Check1_CheckInst_3_n120 ) );
  XNOR2_X1 \Check1_CheckInst_3_U114  ( .A(Red_AddRoundKeyOutput2[23]), .B(
        Red_SignaltoCheck[87]), .ZN(\Check1_CheckInst_3_n111 ) );
  XNOR2_X1 \Check1_CheckInst_3_U113  ( .A(Red_AddRoundKeyOutput2[19]), .B(
        Red_SignaltoCheck[83]), .ZN(\Check1_CheckInst_3_n112 ) );
  NOR2_X1 \Check1_CheckInst_3_U112  ( .A1(\Check1_CheckInst_3_n110 ), .A2(
        \Check1_CheckInst_3_n109 ), .ZN(\Check1_CheckInst_3_n122 ) );
  XOR2_X1 \Check1_CheckInst_3_U111  ( .A(Red_AddRoundKeyOutput3[27]), .B(
        Red_SignaltoCheck[27]), .Z(\Check1_CheckInst_3_n109 ) );
  XOR2_X1 \Check1_CheckInst_3_U110  ( .A(Red_AddRoundKeyOutput3[39]), .B(
        Red_SignaltoCheck[39]), .Z(\Check1_CheckInst_3_n110 ) );
  NOR2_X1 \Check1_CheckInst_3_U109  ( .A1(\Check1_CheckInst_3_n108 ), .A2(
        \Check1_CheckInst_3_n107 ), .ZN(\Check1_CheckInst_3_n156 ) );
  NAND2_X1 \Check1_CheckInst_3_U108  ( .A1(\Check1_CheckInst_3_n106 ), .A2(
        \Check1_CheckInst_3_n105 ), .ZN(\Check1_CheckInst_3_n107 ) );
  NOR2_X1 \Check1_CheckInst_3_U107  ( .A1(\Check1_CheckInst_3_n104 ), .A2(
        \Check1_CheckInst_3_n103 ), .ZN(\Check1_CheckInst_3_n105 ) );
  NAND2_X1 \Check1_CheckInst_3_U106  ( .A1(\Check1_CheckInst_3_n102 ), .A2(
        \Check1_CheckInst_3_n101 ), .ZN(\Check1_CheckInst_3_n103 ) );
  XNOR2_X1 \Check1_CheckInst_3_U105  ( .A(Red_AddRoundKeyOutput3[31]), .B(
        Red_SignaltoCheck[31]), .ZN(\Check1_CheckInst_3_n101 ) );
  XNOR2_X1 \Check1_CheckInst_3_U104  ( .A(Red_AddRoundKeyOutput3[35]), .B(
        Red_SignaltoCheck[35]), .ZN(\Check1_CheckInst_3_n102 ) );
  NAND2_X1 \Check1_CheckInst_3_U103  ( .A1(\Check1_CheckInst_3_n100 ), .A2(
        \Check1_CheckInst_3_n99 ), .ZN(\Check1_CheckInst_3_n104 ) );
  XNOR2_X1 \Check1_CheckInst_3_U102  ( .A(Red_AddRoundKeyOutput3[47]), .B(
        Red_SignaltoCheck[47]), .ZN(\Check1_CheckInst_3_n99 ) );
  XNOR2_X1 \Check1_CheckInst_3_U101  ( .A(Red_AddRoundKeyOutput3[43]), .B(
        Red_SignaltoCheck[43]), .ZN(\Check1_CheckInst_3_n100 ) );
  NOR2_X1 \Check1_CheckInst_3_U100  ( .A1(\Check1_CheckInst_3_n98 ), .A2(
        \Check1_CheckInst_3_n97 ), .ZN(\Check1_CheckInst_3_n106 ) );
  XOR2_X1 \Check1_CheckInst_3_U99  ( .A(Red_AddRoundKeyOutput3[11]), .B(
        Red_SignaltoCheck[11]), .Z(\Check1_CheckInst_3_n97 ) );
  XOR2_X1 \Check1_CheckInst_3_U98  ( .A(Red_AddRoundKeyOutput3[51]), .B(
        Red_SignaltoCheck[51]), .Z(\Check1_CheckInst_3_n98 ) );
  NAND2_X1 \Check1_CheckInst_3_U97  ( .A1(\Check1_CheckInst_3_n96 ), .A2(
        \Check1_CheckInst_3_n95 ), .ZN(\Check1_CheckInst_3_n108 ) );
  XNOR2_X1 \Check1_CheckInst_3_U96  ( .A(Red_StateRegOutput[63]), .B(
        Red_SignaltoCheck[447]), .ZN(\Check1_CheckInst_3_n95 ) );
  XNOR2_X1 \Check1_CheckInst_3_U95  ( .A(Red_SignaltoCheck[3]), .B(
        Red_AddRoundKeyOutput3[3]), .ZN(\Check1_CheckInst_3_n96 ) );
  NOR2_X1 \Check1_CheckInst_3_U94  ( .A1(\Check1_CheckInst_3_n94 ), .A2(
        \Check1_CheckInst_3_n93 ), .ZN(\Check1_CheckInst_3_n222 ) );
  NAND2_X1 \Check1_CheckInst_3_U93  ( .A1(\Check1_CheckInst_3_n92 ), .A2(
        \Check1_CheckInst_3_n91 ), .ZN(\Check1_CheckInst_3_n93 ) );
  NOR2_X1 \Check1_CheckInst_3_U92  ( .A1(\Check1_CheckInst_3_n90 ), .A2(
        \Check1_CheckInst_3_n89 ), .ZN(\Check1_CheckInst_3_n91 ) );
  NAND2_X1 \Check1_CheckInst_3_U91  ( .A1(\Check1_CheckInst_3_n88 ), .A2(
        \Check1_CheckInst_3_n87 ), .ZN(\Check1_CheckInst_3_n89 ) );
  NOR2_X1 \Check1_CheckInst_3_U90  ( .A1(\Check1_CheckInst_3_n86 ), .A2(
        \Check1_CheckInst_3_n85 ), .ZN(\Check1_CheckInst_3_n87 ) );
  NAND2_X1 \Check1_CheckInst_3_U89  ( .A1(\Check1_CheckInst_3_n84 ), .A2(
        \Check1_CheckInst_3_n83 ), .ZN(\Check1_CheckInst_3_n85 ) );
  NOR2_X1 \Check1_CheckInst_3_U88  ( .A1(\Check1_CheckInst_3_n82 ), .A2(
        \Check1_CheckInst_3_n81 ), .ZN(\Check1_CheckInst_3_n83 ) );
  XOR2_X1 \Check1_CheckInst_3_U87  ( .A(Red_AddRoundKeyOutput3[15]), .B(
        Red_SignaltoCheck[15]), .Z(\Check1_CheckInst_3_n81 ) );
  XOR2_X1 \Check1_CheckInst_3_U86  ( .A(Red_SignaltoCheck[7]), .B(
        Red_AddRoundKeyOutput3[7]), .Z(\Check1_CheckInst_3_n82 ) );
  NOR2_X1 \Check1_CheckInst_3_U85  ( .A1(\Check1_CheckInst_3_n80 ), .A2(
        \Check1_CheckInst_3_n79 ), .ZN(\Check1_CheckInst_3_n84 ) );
  XOR2_X1 \Check1_CheckInst_3_U84  ( .A(Red_AddRoundKeyOutput3[23]), .B(
        Red_SignaltoCheck[23]), .Z(\Check1_CheckInst_3_n79 ) );
  XOR2_X1 \Check1_CheckInst_3_U83  ( .A(Red_AddRoundKeyOutput3[19]), .B(
        Red_SignaltoCheck[19]), .Z(\Check1_CheckInst_3_n80 ) );
  NAND2_X1 \Check1_CheckInst_3_U82  ( .A1(\Check1_CheckInst_3_n78 ), .A2(
        \Check1_CheckInst_3_n77 ), .ZN(\Check1_CheckInst_3_n86 ) );
  XNOR2_X1 \Check1_CheckInst_3_U81  ( .A(Red_AddRoundKeyOutput[63]), .B(
        Red_SignaltoCheck[191]), .ZN(\Check1_CheckInst_3_n77 ) );
  XNOR2_X1 \Check1_CheckInst_3_U80  ( .A(Red_AddRoundKeyOutput[59]), .B(
        Red_SignaltoCheck[187]), .ZN(\Check1_CheckInst_3_n78 ) );
  NOR2_X1 \Check1_CheckInst_3_U79  ( .A1(\Check1_CheckInst_3_n76 ), .A2(
        \Check1_CheckInst_3_n75 ), .ZN(\Check1_CheckInst_3_n88 ) );
  XOR2_X1 \Check1_CheckInst_3_U78  ( .A(Red_AddRoundKeyOutput[47]), .B(
        Red_SignaltoCheck[175]), .Z(\Check1_CheckInst_3_n75 ) );
  XOR2_X1 \Check1_CheckInst_3_U77  ( .A(Red_AddRoundKeyOutput[55]), .B(
        Red_SignaltoCheck[183]), .Z(\Check1_CheckInst_3_n76 ) );
  NAND2_X1 \Check1_CheckInst_3_U76  ( .A1(\Check1_CheckInst_3_n74 ), .A2(
        \Check1_CheckInst_3_n73 ), .ZN(\Check1_CheckInst_3_n90 ) );
  NOR2_X1 \Check1_CheckInst_3_U75  ( .A1(\Check1_CheckInst_3_n72 ), .A2(
        \Check1_CheckInst_3_n71 ), .ZN(\Check1_CheckInst_3_n73 ) );
  NAND2_X1 \Check1_CheckInst_3_U74  ( .A1(\Check1_CheckInst_3_n70 ), .A2(
        \Check1_CheckInst_3_n69 ), .ZN(\Check1_CheckInst_3_n71 ) );
  NOR2_X1 \Check1_CheckInst_3_U73  ( .A1(\Check1_CheckInst_3_n68 ), .A2(
        \Check1_CheckInst_3_n67 ), .ZN(\Check1_CheckInst_3_n69 ) );
  XOR2_X1 \Check1_CheckInst_3_U72  ( .A(Red_AddRoundKeyOutput[39]), .B(
        Red_SignaltoCheck[167]), .Z(\Check1_CheckInst_3_n67 ) );
  XOR2_X1 \Check1_CheckInst_3_U71  ( .A(Red_AddRoundKeyOutput[51]), .B(
        Red_SignaltoCheck[179]), .Z(\Check1_CheckInst_3_n68 ) );
  NOR2_X1 \Check1_CheckInst_3_U70  ( .A1(\Check1_CheckInst_3_n66 ), .A2(
        \Check1_CheckInst_3_n65 ), .ZN(\Check1_CheckInst_3_n70 ) );
  XOR2_X1 \Check1_CheckInst_3_U69  ( .A(Red_Feedback3[23]), .B(
        Red_SignaltoCheck[215]), .Z(\Check1_CheckInst_3_n65 ) );
  XOR2_X1 \Check1_CheckInst_3_U68  ( .A(Red_AddRoundKeyOutput[43]), .B(
        Red_SignaltoCheck[171]), .Z(\Check1_CheckInst_3_n66 ) );
  NAND2_X1 \Check1_CheckInst_3_U67  ( .A1(\Check1_CheckInst_3_n64 ), .A2(
        \Check1_CheckInst_3_n63 ), .ZN(\Check1_CheckInst_3_n72 ) );
  XNOR2_X1 \Check1_CheckInst_3_U66  ( .A(Red_Feedback3[19]), .B(
        Red_SignaltoCheck[211]), .ZN(\Check1_CheckInst_3_n63 ) );
  XNOR2_X1 \Check1_CheckInst_3_U65  ( .A(Red_Feedback3[27]), .B(
        Red_SignaltoCheck[219]), .ZN(\Check1_CheckInst_3_n64 ) );
  NOR2_X1 \Check1_CheckInst_3_U64  ( .A1(\Check1_CheckInst_3_n62 ), .A2(
        \Check1_CheckInst_3_n61 ), .ZN(\Check1_CheckInst_3_n74 ) );
  XOR2_X1 \Check1_CheckInst_3_U63  ( .A(Red_Feedback3[15]), .B(
        Red_SignaltoCheck[207]), .Z(\Check1_CheckInst_3_n61 ) );
  XOR2_X1 \Check1_CheckInst_3_U62  ( .A(Red_Feedback3[11]), .B(
        Red_SignaltoCheck[203]), .Z(\Check1_CheckInst_3_n62 ) );
  NOR2_X1 \Check1_CheckInst_3_U61  ( .A1(\Check1_CheckInst_3_n60 ), .A2(
        \Check1_CheckInst_3_n59 ), .ZN(\Check1_CheckInst_3_n92 ) );
  NAND2_X1 \Check1_CheckInst_3_U60  ( .A1(\Check1_CheckInst_3_n58 ), .A2(
        \Check1_CheckInst_3_n57 ), .ZN(\Check1_CheckInst_3_n59 ) );
  NOR2_X1 \Check1_CheckInst_3_U59  ( .A1(\Check1_CheckInst_3_n56 ), .A2(
        \Check1_CheckInst_3_n55 ), .ZN(\Check1_CheckInst_3_n57 ) );
  NAND2_X1 \Check1_CheckInst_3_U58  ( .A1(\Check1_CheckInst_3_n54 ), .A2(
        \Check1_CheckInst_3_n53 ), .ZN(\Check1_CheckInst_3_n55 ) );
  XNOR2_X1 \Check1_CheckInst_3_U57  ( .A(Red_Feedback3[7]), .B(
        Red_SignaltoCheck[199]), .ZN(\Check1_CheckInst_3_n53 ) );
  XNOR2_X1 \Check1_CheckInst_3_U56  ( .A(Red_Feedback3[3]), .B(
        Red_SignaltoCheck[195]), .ZN(\Check1_CheckInst_3_n54 ) );
  NAND2_X1 \Check1_CheckInst_3_U55  ( .A1(\Check1_CheckInst_3_n52 ), .A2(
        \Check1_CheckInst_3_n51 ), .ZN(\Check1_CheckInst_3_n56 ) );
  XNOR2_X1 \Check1_CheckInst_3_U54  ( .A(Red_AddRoundKeyOutput[7]), .B(
        Red_SignaltoCheck[135]), .ZN(\Check1_CheckInst_3_n51 ) );
  XNOR2_X1 \Check1_CheckInst_3_U53  ( .A(Red_AddRoundKeyOutput[3]), .B(
        Red_SignaltoCheck[131]), .ZN(\Check1_CheckInst_3_n52 ) );
  NOR2_X1 \Check1_CheckInst_3_U52  ( .A1(\Check1_CheckInst_3_n50 ), .A2(
        \Check1_CheckInst_3_n49 ), .ZN(\Check1_CheckInst_3_n58 ) );
  XOR2_X1 \Check1_CheckInst_3_U51  ( .A(Red_AddRoundKeyOutput2[55]), .B(
        Red_SignaltoCheck[119]), .Z(\Check1_CheckInst_3_n49 ) );
  XOR2_X1 \Check1_CheckInst_3_U50  ( .A(Red_AddRoundKeyOutput2[63]), .B(
        Red_SignaltoCheck[127]), .Z(\Check1_CheckInst_3_n50 ) );
  NAND2_X1 \Check1_CheckInst_3_U49  ( .A1(\Check1_CheckInst_3_n48 ), .A2(
        \Check1_CheckInst_3_n47 ), .ZN(\Check1_CheckInst_3_n60 ) );
  XNOR2_X1 \Check1_CheckInst_3_U48  ( .A(Red_AddRoundKeyOutput2[47]), .B(
        Red_SignaltoCheck[111]), .ZN(\Check1_CheckInst_3_n47 ) );
  XNOR2_X1 \Check1_CheckInst_3_U47  ( .A(Red_AddRoundKeyOutput2[59]), .B(
        Red_SignaltoCheck[123]), .ZN(\Check1_CheckInst_3_n48 ) );
  NAND2_X1 \Check1_CheckInst_3_U46  ( .A1(\Check1_CheckInst_3_n46 ), .A2(
        \Check1_CheckInst_3_n45 ), .ZN(\Check1_CheckInst_3_n94 ) );
  NOR2_X1 \Check1_CheckInst_3_U45  ( .A1(\Check1_CheckInst_3_n44 ), .A2(
        \Check1_CheckInst_3_n43 ), .ZN(\Check1_CheckInst_3_n45 ) );
  NAND2_X1 \Check1_CheckInst_3_U44  ( .A1(\Check1_CheckInst_3_n42 ), .A2(
        \Check1_CheckInst_3_n41 ), .ZN(\Check1_CheckInst_3_n43 ) );
  NOR2_X1 \Check1_CheckInst_3_U43  ( .A1(\Check1_CheckInst_3_n40 ), .A2(
        \Check1_CheckInst_3_n39 ), .ZN(\Check1_CheckInst_3_n41 ) );
  XOR2_X1 \Check1_CheckInst_3_U42  ( .A(Red_AddRoundKeyOutput[31]), .B(
        Red_SignaltoCheck[159]), .Z(\Check1_CheckInst_3_n39 ) );
  XOR2_X1 \Check1_CheckInst_3_U41  ( .A(Red_AddRoundKeyOutput2[51]), .B(
        Red_SignaltoCheck[115]), .Z(\Check1_CheckInst_3_n40 ) );
  NOR2_X1 \Check1_CheckInst_3_U40  ( .A1(\Check1_CheckInst_3_n38 ), .A2(
        \Check1_CheckInst_3_n37 ), .ZN(\Check1_CheckInst_3_n42 ) );
  XOR2_X1 \Check1_CheckInst_3_U39  ( .A(Red_AddRoundKeyOutput[27]), .B(
        Red_SignaltoCheck[155]), .Z(\Check1_CheckInst_3_n37 ) );
  XOR2_X1 \Check1_CheckInst_3_U38  ( .A(Red_AddRoundKeyOutput[35]), .B(
        Red_SignaltoCheck[163]), .Z(\Check1_CheckInst_3_n38 ) );
  NAND2_X1 \Check1_CheckInst_3_U37  ( .A1(\Check1_CheckInst_3_n36 ), .A2(
        \Check1_CheckInst_3_n35 ), .ZN(\Check1_CheckInst_3_n44 ) );
  XNOR2_X1 \Check1_CheckInst_3_U36  ( .A(Red_AddRoundKeyOutput[23]), .B(
        Red_SignaltoCheck[151]), .ZN(\Check1_CheckInst_3_n35 ) );
  XNOR2_X1 \Check1_CheckInst_3_U35  ( .A(Red_AddRoundKeyOutput[19]), .B(
        Red_SignaltoCheck[147]), .ZN(\Check1_CheckInst_3_n36 ) );
  NOR2_X1 \Check1_CheckInst_3_U34  ( .A1(\Check1_CheckInst_3_n34 ), .A2(
        \Check1_CheckInst_3_n33 ), .ZN(\Check1_CheckInst_3_n46 ) );
  XOR2_X1 \Check1_CheckInst_3_U33  ( .A(Red_AddRoundKeyOutput[15]), .B(
        Red_SignaltoCheck[143]), .Z(\Check1_CheckInst_3_n33 ) );
  XOR2_X1 \Check1_CheckInst_3_U32  ( .A(Red_AddRoundKeyOutput[11]), .B(
        Red_SignaltoCheck[139]), .Z(\Check1_CheckInst_3_n34 ) );
  NAND2_X1 \Check1_CheckInst_3_U31  ( .A1(\Check1_CheckInst_3_n32 ), .A2(
        \Check1_CheckInst_3_n31 ), .ZN(\Check1_CheckInst_3_n224 ) );
  NOR2_X1 \Check1_CheckInst_3_U30  ( .A1(\Check1_CheckInst_3_n30 ), .A2(
        \Check1_CheckInst_3_n29 ), .ZN(\Check1_CheckInst_3_n31 ) );
  NAND2_X1 \Check1_CheckInst_3_U29  ( .A1(\Check1_CheckInst_3_n28 ), .A2(
        \Check1_CheckInst_3_n27 ), .ZN(\Check1_CheckInst_3_n29 ) );
  NOR2_X1 \Check1_CheckInst_3_U28  ( .A1(\Check1_CheckInst_3_n26 ), .A2(
        \Check1_CheckInst_3_n25 ), .ZN(\Check1_CheckInst_3_n27 ) );
  NAND2_X1 \Check1_CheckInst_3_U27  ( .A1(\Check1_CheckInst_3_n24 ), .A2(
        \Check1_CheckInst_3_n23 ), .ZN(\Check1_CheckInst_3_n25 ) );
  XNOR2_X1 \Check1_CheckInst_3_U26  ( .A(Red_StateRegOutput3[31]), .B(
        Red_SignaltoCheck[287]), .ZN(\Check1_CheckInst_3_n23 ) );
  XNOR2_X1 \Check1_CheckInst_3_U25  ( .A(Red_StateRegOutput3[39]), .B(
        Red_SignaltoCheck[295]), .ZN(\Check1_CheckInst_3_n24 ) );
  NAND2_X1 \Check1_CheckInst_3_U24  ( .A1(\Check1_CheckInst_3_n22 ), .A2(
        \Check1_CheckInst_3_n21 ), .ZN(\Check1_CheckInst_3_n26 ) );
  XNOR2_X1 \Check1_CheckInst_3_U23  ( .A(Red_StateRegOutput3[47]), .B(
        Red_SignaltoCheck[303]), .ZN(\Check1_CheckInst_3_n21 ) );
  XNOR2_X1 \Check1_CheckInst_3_U22  ( .A(Red_StateRegOutput3[43]), .B(
        Red_SignaltoCheck[299]), .ZN(\Check1_CheckInst_3_n22 ) );
  NOR2_X1 \Check1_CheckInst_3_U21  ( .A1(\Check1_CheckInst_3_n20 ), .A2(
        \Check1_CheckInst_3_n19 ), .ZN(\Check1_CheckInst_3_n28 ) );
  NAND2_X1 \Check1_CheckInst_3_U20  ( .A1(\Check1_CheckInst_3_n18 ), .A2(
        \Check1_CheckInst_3_n17 ), .ZN(\Check1_CheckInst_3_n19 ) );
  XNOR2_X1 \Check1_CheckInst_3_U19  ( .A(Red_StateRegOutput2[7]), .B(
        Red_SignaltoCheck[327]), .ZN(\Check1_CheckInst_3_n17 ) );
  XNOR2_X1 \Check1_CheckInst_3_U18  ( .A(Red_StateRegOutput3[27]), .B(
        Red_SignaltoCheck[283]), .ZN(\Check1_CheckInst_3_n18 ) );
  NAND2_X1 \Check1_CheckInst_3_U17  ( .A1(\Check1_CheckInst_3_n16 ), .A2(
        \Check1_CheckInst_3_n15 ), .ZN(\Check1_CheckInst_3_n20 ) );
  XNOR2_X1 \Check1_CheckInst_3_U16  ( .A(Red_StateRegOutput3[23]), .B(
        Red_SignaltoCheck[279]), .ZN(\Check1_CheckInst_3_n15 ) );
  XNOR2_X1 \Check1_CheckInst_3_U15  ( .A(Red_StateRegOutput3[35]), .B(
        Red_SignaltoCheck[291]), .ZN(\Check1_CheckInst_3_n16 ) );
  NAND2_X1 \Check1_CheckInst_3_U14  ( .A1(\Check1_CheckInst_3_n14 ), .A2(
        \Check1_CheckInst_3_n13 ), .ZN(\Check1_CheckInst_3_n30 ) );
  NOR2_X1 \Check1_CheckInst_3_U13  ( .A1(\Check1_CheckInst_3_n12 ), .A2(
        \Check1_CheckInst_3_n11 ), .ZN(\Check1_CheckInst_3_n13 ) );
  XOR2_X1 \Check1_CheckInst_3_U12  ( .A(Red_StateRegOutput3[63]), .B(
        Red_SignaltoCheck[319]), .Z(\Check1_CheckInst_3_n11 ) );
  XOR2_X1 \Check1_CheckInst_3_U11  ( .A(Red_StateRegOutput3[59]), .B(
        Red_SignaltoCheck[315]), .Z(\Check1_CheckInst_3_n12 ) );
  NOR2_X1 \Check1_CheckInst_3_U10  ( .A1(\Check1_CheckInst_3_n10 ), .A2(
        \Check1_CheckInst_3_n9 ), .ZN(\Check1_CheckInst_3_n14 ) );
  XOR2_X1 \Check1_CheckInst_3_U9  ( .A(Red_StateRegOutput2[3]), .B(
        Red_SignaltoCheck[323]), .Z(\Check1_CheckInst_3_n9 ) );
  XOR2_X1 \Check1_CheckInst_3_U8  ( .A(Red_StateRegOutput2[11]), .B(
        Red_SignaltoCheck[331]), .Z(\Check1_CheckInst_3_n10 ) );
  NOR2_X1 \Check1_CheckInst_3_U7  ( .A1(\Check1_CheckInst_3_n8 ), .A2(
        \Check1_CheckInst_3_n7 ), .ZN(\Check1_CheckInst_3_n32 ) );
  NAND2_X1 \Check1_CheckInst_3_U6  ( .A1(\Check1_CheckInst_3_n6 ), .A2(
        \Check1_CheckInst_3_n5 ), .ZN(\Check1_CheckInst_3_n7 ) );
  XNOR2_X1 \Check1_CheckInst_3_U5  ( .A(Red_Feedback3[55]), .B(
        Red_SignaltoCheck[247]), .ZN(\Check1_CheckInst_3_n5 ) );
  XNOR2_X1 \Check1_CheckInst_3_U4  ( .A(Red_Feedback3[51]), .B(
        Red_SignaltoCheck[243]), .ZN(\Check1_CheckInst_3_n6 ) );
  NAND2_X1 \Check1_CheckInst_3_U3  ( .A1(\Check1_CheckInst_3_n4 ), .A2(
        \Check1_CheckInst_3_n3 ), .ZN(\Check1_CheckInst_3_n8 ) );
  XNOR2_X1 \Check1_CheckInst_3_U2  ( .A(Red_StateRegOutput3[55]), .B(
        Red_SignaltoCheck[311]), .ZN(\Check1_CheckInst_3_n3 ) );
  XNOR2_X1 \Check1_CheckInst_3_U1  ( .A(Red_StateRegOutput3[51]), .B(
        Red_SignaltoCheck[307]), .ZN(\Check1_CheckInst_3_n4 ) );
endmodule

