
module Cipher ( clk, rst, Input, Key, Output, ErrorFlag );
  input [63:0] Input;
  input [127:0] Key;
  output [63:0] Output;
  (* FIRMER="clock" *)input clk;
  (* FIRMER="control" *)input rst;
  output ErrorFlag;
  wire   MCOutput_63_, MCOutput_62_, MCOutput_61_, MCOutput_60_, MCOutput_59_,
         MCOutput_58_, MCOutput_57_, MCOutput_56_, MCOutput_55_, MCOutput_54_,
         MCOutput_53_, MCOutput_52_, MCOutput_51_, MCOutput_50_, MCOutput_49_,
         MCOutput_48_, MCOutput_47_, MCOutput_46_, MCOutput_45_, MCOutput_44_,
         MCOutput_43_, MCOutput_42_, MCOutput_41_, MCOutput_40_, MCOutput_39_,
         MCOutput_38_, MCOutput_37_, MCOutput_36_, MCOutput_35_, MCOutput_34_,
         MCOutput_33_, MCOutput_32_, Error_0_, MCInst_XOR_r0_Inst_0_n5,
         MCInst_XOR_r0_Inst_1_n5, MCInst_XOR_r0_Inst_2_n5,
         MCInst_XOR_r0_Inst_3_n5, MCInst_XOR_r0_Inst_4_n5,
         MCInst_XOR_r0_Inst_5_n5, MCInst_XOR_r0_Inst_6_n5,
         MCInst_XOR_r0_Inst_7_n5, MCInst_XOR_r0_Inst_8_n5,
         MCInst_XOR_r0_Inst_9_n5, MCInst_XOR_r0_Inst_10_n5,
         MCInst_XOR_r0_Inst_11_n5, MCInst_XOR_r0_Inst_12_n5,
         MCInst_XOR_r0_Inst_13_n5, MCInst_XOR_r0_Inst_14_n5,
         MCInst_XOR_r0_Inst_15_n5, SubCellInst_LFInst_0_LFInst_0_n15,
         SubCellInst_LFInst_0_LFInst_0_n14, SubCellInst_LFInst_0_LFInst_0_n13,
         SubCellInst_LFInst_0_LFInst_0_n12, SubCellInst_LFInst_0_LFInst_0_n11,
         SubCellInst_LFInst_0_LFInst_1_n9, SubCellInst_LFInst_0_LFInst_1_n8,
         SubCellInst_LFInst_0_LFInst_1_n7, SubCellInst_LFInst_0_LFInst_2_n18,
         SubCellInst_LFInst_0_LFInst_2_n17, SubCellInst_LFInst_0_LFInst_2_n16,
         SubCellInst_LFInst_0_LFInst_2_n15, SubCellInst_LFInst_0_LFInst_2_n14,
         SubCellInst_LFInst_0_LFInst_3_n9, SubCellInst_LFInst_0_LFInst_3_n8,
         SubCellInst_LFInst_0_LFInst_3_n7, SubCellInst_LFInst_1_LFInst_0_n15,
         SubCellInst_LFInst_1_LFInst_0_n14, SubCellInst_LFInst_1_LFInst_0_n13,
         SubCellInst_LFInst_1_LFInst_0_n12, SubCellInst_LFInst_1_LFInst_0_n11,
         SubCellInst_LFInst_1_LFInst_1_n9, SubCellInst_LFInst_1_LFInst_1_n8,
         SubCellInst_LFInst_1_LFInst_1_n7, SubCellInst_LFInst_1_LFInst_2_n18,
         SubCellInst_LFInst_1_LFInst_2_n17, SubCellInst_LFInst_1_LFInst_2_n16,
         SubCellInst_LFInst_1_LFInst_2_n15, SubCellInst_LFInst_1_LFInst_2_n14,
         SubCellInst_LFInst_1_LFInst_3_n9, SubCellInst_LFInst_1_LFInst_3_n8,
         SubCellInst_LFInst_1_LFInst_3_n7, SubCellInst_LFInst_2_LFInst_0_n15,
         SubCellInst_LFInst_2_LFInst_0_n14, SubCellInst_LFInst_2_LFInst_0_n13,
         SubCellInst_LFInst_2_LFInst_0_n12, SubCellInst_LFInst_2_LFInst_0_n11,
         SubCellInst_LFInst_2_LFInst_1_n9, SubCellInst_LFInst_2_LFInst_1_n8,
         SubCellInst_LFInst_2_LFInst_1_n7, SubCellInst_LFInst_2_LFInst_2_n18,
         SubCellInst_LFInst_2_LFInst_2_n17, SubCellInst_LFInst_2_LFInst_2_n16,
         SubCellInst_LFInst_2_LFInst_2_n15, SubCellInst_LFInst_2_LFInst_2_n14,
         SubCellInst_LFInst_2_LFInst_3_n9, SubCellInst_LFInst_2_LFInst_3_n8,
         SubCellInst_LFInst_2_LFInst_3_n7, SubCellInst_LFInst_3_LFInst_0_n15,
         SubCellInst_LFInst_3_LFInst_0_n14, SubCellInst_LFInst_3_LFInst_0_n13,
         SubCellInst_LFInst_3_LFInst_0_n12, SubCellInst_LFInst_3_LFInst_0_n11,
         SubCellInst_LFInst_3_LFInst_1_n9, SubCellInst_LFInst_3_LFInst_1_n8,
         SubCellInst_LFInst_3_LFInst_1_n7, SubCellInst_LFInst_3_LFInst_2_n18,
         SubCellInst_LFInst_3_LFInst_2_n17, SubCellInst_LFInst_3_LFInst_2_n16,
         SubCellInst_LFInst_3_LFInst_2_n15, SubCellInst_LFInst_3_LFInst_2_n14,
         SubCellInst_LFInst_3_LFInst_3_n9, SubCellInst_LFInst_3_LFInst_3_n8,
         SubCellInst_LFInst_3_LFInst_3_n7, SubCellInst_LFInst_4_LFInst_0_n15,
         SubCellInst_LFInst_4_LFInst_0_n14, SubCellInst_LFInst_4_LFInst_0_n13,
         SubCellInst_LFInst_4_LFInst_0_n12, SubCellInst_LFInst_4_LFInst_0_n11,
         SubCellInst_LFInst_4_LFInst_1_n9, SubCellInst_LFInst_4_LFInst_1_n8,
         SubCellInst_LFInst_4_LFInst_1_n7, SubCellInst_LFInst_4_LFInst_2_n18,
         SubCellInst_LFInst_4_LFInst_2_n17, SubCellInst_LFInst_4_LFInst_2_n16,
         SubCellInst_LFInst_4_LFInst_2_n15, SubCellInst_LFInst_4_LFInst_2_n14,
         SubCellInst_LFInst_4_LFInst_3_n9, SubCellInst_LFInst_4_LFInst_3_n8,
         SubCellInst_LFInst_4_LFInst_3_n7, SubCellInst_LFInst_5_LFInst_0_n15,
         SubCellInst_LFInst_5_LFInst_0_n14, SubCellInst_LFInst_5_LFInst_0_n13,
         SubCellInst_LFInst_5_LFInst_0_n12, SubCellInst_LFInst_5_LFInst_0_n11,
         SubCellInst_LFInst_5_LFInst_1_n9, SubCellInst_LFInst_5_LFInst_1_n8,
         SubCellInst_LFInst_5_LFInst_1_n7, SubCellInst_LFInst_5_LFInst_2_n18,
         SubCellInst_LFInst_5_LFInst_2_n17, SubCellInst_LFInst_5_LFInst_2_n16,
         SubCellInst_LFInst_5_LFInst_2_n15, SubCellInst_LFInst_5_LFInst_2_n14,
         SubCellInst_LFInst_5_LFInst_3_n9, SubCellInst_LFInst_5_LFInst_3_n8,
         SubCellInst_LFInst_5_LFInst_3_n7, SubCellInst_LFInst_6_LFInst_0_n15,
         SubCellInst_LFInst_6_LFInst_0_n14, SubCellInst_LFInst_6_LFInst_0_n13,
         SubCellInst_LFInst_6_LFInst_0_n12, SubCellInst_LFInst_6_LFInst_0_n11,
         SubCellInst_LFInst_6_LFInst_1_n9, SubCellInst_LFInst_6_LFInst_1_n8,
         SubCellInst_LFInst_6_LFInst_1_n7, SubCellInst_LFInst_6_LFInst_2_n18,
         SubCellInst_LFInst_6_LFInst_2_n17, SubCellInst_LFInst_6_LFInst_2_n16,
         SubCellInst_LFInst_6_LFInst_2_n15, SubCellInst_LFInst_6_LFInst_2_n14,
         SubCellInst_LFInst_6_LFInst_3_n9, SubCellInst_LFInst_6_LFInst_3_n8,
         SubCellInst_LFInst_6_LFInst_3_n7, SubCellInst_LFInst_7_LFInst_0_n15,
         SubCellInst_LFInst_7_LFInst_0_n14, SubCellInst_LFInst_7_LFInst_0_n13,
         SubCellInst_LFInst_7_LFInst_0_n12, SubCellInst_LFInst_7_LFInst_0_n11,
         SubCellInst_LFInst_7_LFInst_1_n9, SubCellInst_LFInst_7_LFInst_1_n8,
         SubCellInst_LFInst_7_LFInst_1_n7, SubCellInst_LFInst_7_LFInst_2_n18,
         SubCellInst_LFInst_7_LFInst_2_n17, SubCellInst_LFInst_7_LFInst_2_n16,
         SubCellInst_LFInst_7_LFInst_2_n15, SubCellInst_LFInst_7_LFInst_2_n14,
         SubCellInst_LFInst_7_LFInst_3_n9, SubCellInst_LFInst_7_LFInst_3_n8,
         SubCellInst_LFInst_7_LFInst_3_n7, SubCellInst_LFInst_8_LFInst_0_n15,
         SubCellInst_LFInst_8_LFInst_0_n14, SubCellInst_LFInst_8_LFInst_0_n13,
         SubCellInst_LFInst_8_LFInst_0_n12, SubCellInst_LFInst_8_LFInst_0_n11,
         SubCellInst_LFInst_8_LFInst_1_n9, SubCellInst_LFInst_8_LFInst_1_n8,
         SubCellInst_LFInst_8_LFInst_1_n7, SubCellInst_LFInst_8_LFInst_2_n18,
         SubCellInst_LFInst_8_LFInst_2_n17, SubCellInst_LFInst_8_LFInst_2_n16,
         SubCellInst_LFInst_8_LFInst_2_n15, SubCellInst_LFInst_8_LFInst_2_n14,
         SubCellInst_LFInst_8_LFInst_3_n9, SubCellInst_LFInst_8_LFInst_3_n8,
         SubCellInst_LFInst_8_LFInst_3_n7, SubCellInst_LFInst_9_LFInst_0_n15,
         SubCellInst_LFInst_9_LFInst_0_n14, SubCellInst_LFInst_9_LFInst_0_n13,
         SubCellInst_LFInst_9_LFInst_0_n12, SubCellInst_LFInst_9_LFInst_0_n11,
         SubCellInst_LFInst_9_LFInst_1_n9, SubCellInst_LFInst_9_LFInst_1_n8,
         SubCellInst_LFInst_9_LFInst_1_n7, SubCellInst_LFInst_9_LFInst_2_n18,
         SubCellInst_LFInst_9_LFInst_2_n17, SubCellInst_LFInst_9_LFInst_2_n16,
         SubCellInst_LFInst_9_LFInst_2_n15, SubCellInst_LFInst_9_LFInst_2_n14,
         SubCellInst_LFInst_9_LFInst_3_n9, SubCellInst_LFInst_9_LFInst_3_n8,
         SubCellInst_LFInst_9_LFInst_3_n7, SubCellInst_LFInst_10_LFInst_0_n15,
         SubCellInst_LFInst_10_LFInst_0_n14,
         SubCellInst_LFInst_10_LFInst_0_n13,
         SubCellInst_LFInst_10_LFInst_0_n12,
         SubCellInst_LFInst_10_LFInst_0_n11, SubCellInst_LFInst_10_LFInst_1_n9,
         SubCellInst_LFInst_10_LFInst_1_n8, SubCellInst_LFInst_10_LFInst_1_n7,
         SubCellInst_LFInst_10_LFInst_2_n18,
         SubCellInst_LFInst_10_LFInst_2_n17,
         SubCellInst_LFInst_10_LFInst_2_n16,
         SubCellInst_LFInst_10_LFInst_2_n15,
         SubCellInst_LFInst_10_LFInst_2_n14, SubCellInst_LFInst_10_LFInst_3_n9,
         SubCellInst_LFInst_10_LFInst_3_n8, SubCellInst_LFInst_10_LFInst_3_n7,
         SubCellInst_LFInst_11_LFInst_0_n15,
         SubCellInst_LFInst_11_LFInst_0_n14,
         SubCellInst_LFInst_11_LFInst_0_n13,
         SubCellInst_LFInst_11_LFInst_0_n12,
         SubCellInst_LFInst_11_LFInst_0_n11, SubCellInst_LFInst_11_LFInst_1_n9,
         SubCellInst_LFInst_11_LFInst_1_n8, SubCellInst_LFInst_11_LFInst_1_n7,
         SubCellInst_LFInst_11_LFInst_2_n18,
         SubCellInst_LFInst_11_LFInst_2_n17,
         SubCellInst_LFInst_11_LFInst_2_n16,
         SubCellInst_LFInst_11_LFInst_2_n15,
         SubCellInst_LFInst_11_LFInst_2_n14, SubCellInst_LFInst_11_LFInst_3_n9,
         SubCellInst_LFInst_11_LFInst_3_n8, SubCellInst_LFInst_11_LFInst_3_n7,
         SubCellInst_LFInst_12_LFInst_0_n15,
         SubCellInst_LFInst_12_LFInst_0_n14,
         SubCellInst_LFInst_12_LFInst_0_n13,
         SubCellInst_LFInst_12_LFInst_0_n12,
         SubCellInst_LFInst_12_LFInst_0_n11, SubCellInst_LFInst_12_LFInst_1_n9,
         SubCellInst_LFInst_12_LFInst_1_n8, SubCellInst_LFInst_12_LFInst_1_n7,
         SubCellInst_LFInst_12_LFInst_2_n18,
         SubCellInst_LFInst_12_LFInst_2_n17,
         SubCellInst_LFInst_12_LFInst_2_n16,
         SubCellInst_LFInst_12_LFInst_2_n15,
         SubCellInst_LFInst_12_LFInst_2_n14, SubCellInst_LFInst_12_LFInst_3_n9,
         SubCellInst_LFInst_12_LFInst_3_n8, SubCellInst_LFInst_12_LFInst_3_n7,
         SubCellInst_LFInst_13_LFInst_0_n15,
         SubCellInst_LFInst_13_LFInst_0_n14,
         SubCellInst_LFInst_13_LFInst_0_n13,
         SubCellInst_LFInst_13_LFInst_0_n12,
         SubCellInst_LFInst_13_LFInst_0_n11, SubCellInst_LFInst_13_LFInst_1_n9,
         SubCellInst_LFInst_13_LFInst_1_n8, SubCellInst_LFInst_13_LFInst_1_n7,
         SubCellInst_LFInst_13_LFInst_2_n18,
         SubCellInst_LFInst_13_LFInst_2_n17,
         SubCellInst_LFInst_13_LFInst_2_n16,
         SubCellInst_LFInst_13_LFInst_2_n15,
         SubCellInst_LFInst_13_LFInst_2_n14, SubCellInst_LFInst_13_LFInst_3_n9,
         SubCellInst_LFInst_13_LFInst_3_n8, SubCellInst_LFInst_13_LFInst_3_n7,
         SubCellInst_LFInst_14_LFInst_0_n15,
         SubCellInst_LFInst_14_LFInst_0_n14,
         SubCellInst_LFInst_14_LFInst_0_n13,
         SubCellInst_LFInst_14_LFInst_0_n12,
         SubCellInst_LFInst_14_LFInst_0_n11, SubCellInst_LFInst_14_LFInst_1_n9,
         SubCellInst_LFInst_14_LFInst_1_n8, SubCellInst_LFInst_14_LFInst_1_n7,
         SubCellInst_LFInst_14_LFInst_2_n18,
         SubCellInst_LFInst_14_LFInst_2_n17,
         SubCellInst_LFInst_14_LFInst_2_n16,
         SubCellInst_LFInst_14_LFInst_2_n15,
         SubCellInst_LFInst_14_LFInst_2_n14, SubCellInst_LFInst_14_LFInst_3_n9,
         SubCellInst_LFInst_14_LFInst_3_n8, SubCellInst_LFInst_14_LFInst_3_n7,
         SubCellInst_LFInst_15_LFInst_0_n15,
         SubCellInst_LFInst_15_LFInst_0_n14,
         SubCellInst_LFInst_15_LFInst_0_n13,
         SubCellInst_LFInst_15_LFInst_0_n12,
         SubCellInst_LFInst_15_LFInst_0_n11, SubCellInst_LFInst_15_LFInst_1_n9,
         SubCellInst_LFInst_15_LFInst_1_n8, SubCellInst_LFInst_15_LFInst_1_n7,
         SubCellInst_LFInst_15_LFInst_2_n18,
         SubCellInst_LFInst_15_LFInst_2_n17,
         SubCellInst_LFInst_15_LFInst_2_n16,
         SubCellInst_LFInst_15_LFInst_2_n15,
         SubCellInst_LFInst_15_LFInst_2_n14, SubCellInst_LFInst_15_LFInst_3_n9,
         SubCellInst_LFInst_15_LFInst_3_n8, SubCellInst_LFInst_15_LFInst_3_n7,
         MCInst2_XOR_r0_Inst_0_n5, MCInst2_XOR_r0_Inst_1_n5,
         MCInst2_XOR_r0_Inst_2_n5, MCInst2_XOR_r0_Inst_3_n5,
         MCInst2_XOR_r0_Inst_4_n5, MCInst2_XOR_r0_Inst_5_n5,
         MCInst2_XOR_r0_Inst_6_n5, MCInst2_XOR_r0_Inst_7_n5,
         MCInst2_XOR_r0_Inst_8_n5, MCInst2_XOR_r0_Inst_9_n5,
         MCInst2_XOR_r0_Inst_10_n5, MCInst2_XOR_r0_Inst_11_n5,
         MCInst2_XOR_r0_Inst_12_n5, MCInst2_XOR_r0_Inst_13_n5,
         MCInst2_XOR_r0_Inst_14_n5, MCInst2_XOR_r0_Inst_15_n5,
         SubCellInst2_LFInst_0_LFInst_0_n15,
         SubCellInst2_LFInst_0_LFInst_0_n14,
         SubCellInst2_LFInst_0_LFInst_0_n13,
         SubCellInst2_LFInst_0_LFInst_0_n12,
         SubCellInst2_LFInst_0_LFInst_0_n11, SubCellInst2_LFInst_0_LFInst_1_n9,
         SubCellInst2_LFInst_0_LFInst_1_n8, SubCellInst2_LFInst_0_LFInst_1_n7,
         SubCellInst2_LFInst_0_LFInst_2_n18,
         SubCellInst2_LFInst_0_LFInst_2_n17,
         SubCellInst2_LFInst_0_LFInst_2_n16,
         SubCellInst2_LFInst_0_LFInst_2_n15,
         SubCellInst2_LFInst_0_LFInst_2_n14, SubCellInst2_LFInst_0_LFInst_3_n9,
         SubCellInst2_LFInst_0_LFInst_3_n8, SubCellInst2_LFInst_0_LFInst_3_n7,
         SubCellInst2_LFInst_1_LFInst_0_n15,
         SubCellInst2_LFInst_1_LFInst_0_n14,
         SubCellInst2_LFInst_1_LFInst_0_n13,
         SubCellInst2_LFInst_1_LFInst_0_n12,
         SubCellInst2_LFInst_1_LFInst_0_n11, SubCellInst2_LFInst_1_LFInst_1_n9,
         SubCellInst2_LFInst_1_LFInst_1_n8, SubCellInst2_LFInst_1_LFInst_1_n7,
         SubCellInst2_LFInst_1_LFInst_2_n18,
         SubCellInst2_LFInst_1_LFInst_2_n17,
         SubCellInst2_LFInst_1_LFInst_2_n16,
         SubCellInst2_LFInst_1_LFInst_2_n15,
         SubCellInst2_LFInst_1_LFInst_2_n14, SubCellInst2_LFInst_1_LFInst_3_n9,
         SubCellInst2_LFInst_1_LFInst_3_n8, SubCellInst2_LFInst_1_LFInst_3_n7,
         SubCellInst2_LFInst_2_LFInst_0_n15,
         SubCellInst2_LFInst_2_LFInst_0_n14,
         SubCellInst2_LFInst_2_LFInst_0_n13,
         SubCellInst2_LFInst_2_LFInst_0_n12,
         SubCellInst2_LFInst_2_LFInst_0_n11, SubCellInst2_LFInst_2_LFInst_1_n9,
         SubCellInst2_LFInst_2_LFInst_1_n8, SubCellInst2_LFInst_2_LFInst_1_n7,
         SubCellInst2_LFInst_2_LFInst_2_n18,
         SubCellInst2_LFInst_2_LFInst_2_n17,
         SubCellInst2_LFInst_2_LFInst_2_n16,
         SubCellInst2_LFInst_2_LFInst_2_n15,
         SubCellInst2_LFInst_2_LFInst_2_n14, SubCellInst2_LFInst_2_LFInst_3_n9,
         SubCellInst2_LFInst_2_LFInst_3_n8, SubCellInst2_LFInst_2_LFInst_3_n7,
         SubCellInst2_LFInst_3_LFInst_0_n15,
         SubCellInst2_LFInst_3_LFInst_0_n14,
         SubCellInst2_LFInst_3_LFInst_0_n13,
         SubCellInst2_LFInst_3_LFInst_0_n12,
         SubCellInst2_LFInst_3_LFInst_0_n11, SubCellInst2_LFInst_3_LFInst_1_n9,
         SubCellInst2_LFInst_3_LFInst_1_n8, SubCellInst2_LFInst_3_LFInst_1_n7,
         SubCellInst2_LFInst_3_LFInst_2_n18,
         SubCellInst2_LFInst_3_LFInst_2_n17,
         SubCellInst2_LFInst_3_LFInst_2_n16,
         SubCellInst2_LFInst_3_LFInst_2_n15,
         SubCellInst2_LFInst_3_LFInst_2_n14, SubCellInst2_LFInst_3_LFInst_3_n9,
         SubCellInst2_LFInst_3_LFInst_3_n8, SubCellInst2_LFInst_3_LFInst_3_n7,
         SubCellInst2_LFInst_4_LFInst_0_n15,
         SubCellInst2_LFInst_4_LFInst_0_n14,
         SubCellInst2_LFInst_4_LFInst_0_n13,
         SubCellInst2_LFInst_4_LFInst_0_n12,
         SubCellInst2_LFInst_4_LFInst_0_n11, SubCellInst2_LFInst_4_LFInst_1_n9,
         SubCellInst2_LFInst_4_LFInst_1_n8, SubCellInst2_LFInst_4_LFInst_1_n7,
         SubCellInst2_LFInst_4_LFInst_2_n18,
         SubCellInst2_LFInst_4_LFInst_2_n17,
         SubCellInst2_LFInst_4_LFInst_2_n16,
         SubCellInst2_LFInst_4_LFInst_2_n15,
         SubCellInst2_LFInst_4_LFInst_2_n14, SubCellInst2_LFInst_4_LFInst_3_n9,
         SubCellInst2_LFInst_4_LFInst_3_n8, SubCellInst2_LFInst_4_LFInst_3_n7,
         SubCellInst2_LFInst_5_LFInst_0_n15,
         SubCellInst2_LFInst_5_LFInst_0_n14,
         SubCellInst2_LFInst_5_LFInst_0_n13,
         SubCellInst2_LFInst_5_LFInst_0_n12,
         SubCellInst2_LFInst_5_LFInst_0_n11, SubCellInst2_LFInst_5_LFInst_1_n9,
         SubCellInst2_LFInst_5_LFInst_1_n8, SubCellInst2_LFInst_5_LFInst_1_n7,
         SubCellInst2_LFInst_5_LFInst_2_n18,
         SubCellInst2_LFInst_5_LFInst_2_n17,
         SubCellInst2_LFInst_5_LFInst_2_n16,
         SubCellInst2_LFInst_5_LFInst_2_n15,
         SubCellInst2_LFInst_5_LFInst_2_n14, SubCellInst2_LFInst_5_LFInst_3_n9,
         SubCellInst2_LFInst_5_LFInst_3_n8, SubCellInst2_LFInst_5_LFInst_3_n7,
         SubCellInst2_LFInst_6_LFInst_0_n15,
         SubCellInst2_LFInst_6_LFInst_0_n14,
         SubCellInst2_LFInst_6_LFInst_0_n13,
         SubCellInst2_LFInst_6_LFInst_0_n12,
         SubCellInst2_LFInst_6_LFInst_0_n11, SubCellInst2_LFInst_6_LFInst_1_n9,
         SubCellInst2_LFInst_6_LFInst_1_n8, SubCellInst2_LFInst_6_LFInst_1_n7,
         SubCellInst2_LFInst_6_LFInst_2_n18,
         SubCellInst2_LFInst_6_LFInst_2_n17,
         SubCellInst2_LFInst_6_LFInst_2_n16,
         SubCellInst2_LFInst_6_LFInst_2_n15,
         SubCellInst2_LFInst_6_LFInst_2_n14, SubCellInst2_LFInst_6_LFInst_3_n9,
         SubCellInst2_LFInst_6_LFInst_3_n8, SubCellInst2_LFInst_6_LFInst_3_n7,
         SubCellInst2_LFInst_7_LFInst_0_n15,
         SubCellInst2_LFInst_7_LFInst_0_n14,
         SubCellInst2_LFInst_7_LFInst_0_n13,
         SubCellInst2_LFInst_7_LFInst_0_n12,
         SubCellInst2_LFInst_7_LFInst_0_n11, SubCellInst2_LFInst_7_LFInst_1_n9,
         SubCellInst2_LFInst_7_LFInst_1_n8, SubCellInst2_LFInst_7_LFInst_1_n7,
         SubCellInst2_LFInst_7_LFInst_2_n18,
         SubCellInst2_LFInst_7_LFInst_2_n17,
         SubCellInst2_LFInst_7_LFInst_2_n16,
         SubCellInst2_LFInst_7_LFInst_2_n15,
         SubCellInst2_LFInst_7_LFInst_2_n14, SubCellInst2_LFInst_7_LFInst_3_n9,
         SubCellInst2_LFInst_7_LFInst_3_n8, SubCellInst2_LFInst_7_LFInst_3_n7,
         SubCellInst2_LFInst_8_LFInst_0_n15,
         SubCellInst2_LFInst_8_LFInst_0_n14,
         SubCellInst2_LFInst_8_LFInst_0_n13,
         SubCellInst2_LFInst_8_LFInst_0_n12,
         SubCellInst2_LFInst_8_LFInst_0_n11, SubCellInst2_LFInst_8_LFInst_1_n9,
         SubCellInst2_LFInst_8_LFInst_1_n8, SubCellInst2_LFInst_8_LFInst_1_n7,
         SubCellInst2_LFInst_8_LFInst_2_n18,
         SubCellInst2_LFInst_8_LFInst_2_n17,
         SubCellInst2_LFInst_8_LFInst_2_n16,
         SubCellInst2_LFInst_8_LFInst_2_n15,
         SubCellInst2_LFInst_8_LFInst_2_n14, SubCellInst2_LFInst_8_LFInst_3_n9,
         SubCellInst2_LFInst_8_LFInst_3_n8, SubCellInst2_LFInst_8_LFInst_3_n7,
         SubCellInst2_LFInst_9_LFInst_0_n15,
         SubCellInst2_LFInst_9_LFInst_0_n14,
         SubCellInst2_LFInst_9_LFInst_0_n13,
         SubCellInst2_LFInst_9_LFInst_0_n12,
         SubCellInst2_LFInst_9_LFInst_0_n11, SubCellInst2_LFInst_9_LFInst_1_n9,
         SubCellInst2_LFInst_9_LFInst_1_n8, SubCellInst2_LFInst_9_LFInst_1_n7,
         SubCellInst2_LFInst_9_LFInst_2_n18,
         SubCellInst2_LFInst_9_LFInst_2_n17,
         SubCellInst2_LFInst_9_LFInst_2_n16,
         SubCellInst2_LFInst_9_LFInst_2_n15,
         SubCellInst2_LFInst_9_LFInst_2_n14, SubCellInst2_LFInst_9_LFInst_3_n9,
         SubCellInst2_LFInst_9_LFInst_3_n8, SubCellInst2_LFInst_9_LFInst_3_n7,
         SubCellInst2_LFInst_10_LFInst_0_n15,
         SubCellInst2_LFInst_10_LFInst_0_n14,
         SubCellInst2_LFInst_10_LFInst_0_n13,
         SubCellInst2_LFInst_10_LFInst_0_n12,
         SubCellInst2_LFInst_10_LFInst_0_n11,
         SubCellInst2_LFInst_10_LFInst_1_n9,
         SubCellInst2_LFInst_10_LFInst_1_n8,
         SubCellInst2_LFInst_10_LFInst_1_n7,
         SubCellInst2_LFInst_10_LFInst_2_n18,
         SubCellInst2_LFInst_10_LFInst_2_n17,
         SubCellInst2_LFInst_10_LFInst_2_n16,
         SubCellInst2_LFInst_10_LFInst_2_n15,
         SubCellInst2_LFInst_10_LFInst_2_n14,
         SubCellInst2_LFInst_10_LFInst_3_n9,
         SubCellInst2_LFInst_10_LFInst_3_n8,
         SubCellInst2_LFInst_10_LFInst_3_n7,
         SubCellInst2_LFInst_11_LFInst_0_n15,
         SubCellInst2_LFInst_11_LFInst_0_n14,
         SubCellInst2_LFInst_11_LFInst_0_n13,
         SubCellInst2_LFInst_11_LFInst_0_n12,
         SubCellInst2_LFInst_11_LFInst_0_n11,
         SubCellInst2_LFInst_11_LFInst_1_n9,
         SubCellInst2_LFInst_11_LFInst_1_n8,
         SubCellInst2_LFInst_11_LFInst_1_n7,
         SubCellInst2_LFInst_11_LFInst_2_n18,
         SubCellInst2_LFInst_11_LFInst_2_n17,
         SubCellInst2_LFInst_11_LFInst_2_n16,
         SubCellInst2_LFInst_11_LFInst_2_n15,
         SubCellInst2_LFInst_11_LFInst_2_n14,
         SubCellInst2_LFInst_11_LFInst_3_n9,
         SubCellInst2_LFInst_11_LFInst_3_n8,
         SubCellInst2_LFInst_11_LFInst_3_n7,
         SubCellInst2_LFInst_12_LFInst_0_n15,
         SubCellInst2_LFInst_12_LFInst_0_n14,
         SubCellInst2_LFInst_12_LFInst_0_n13,
         SubCellInst2_LFInst_12_LFInst_0_n12,
         SubCellInst2_LFInst_12_LFInst_0_n11,
         SubCellInst2_LFInst_12_LFInst_1_n9,
         SubCellInst2_LFInst_12_LFInst_1_n8,
         SubCellInst2_LFInst_12_LFInst_1_n7,
         SubCellInst2_LFInst_12_LFInst_2_n18,
         SubCellInst2_LFInst_12_LFInst_2_n17,
         SubCellInst2_LFInst_12_LFInst_2_n16,
         SubCellInst2_LFInst_12_LFInst_2_n15,
         SubCellInst2_LFInst_12_LFInst_2_n14,
         SubCellInst2_LFInst_12_LFInst_3_n9,
         SubCellInst2_LFInst_12_LFInst_3_n8,
         SubCellInst2_LFInst_12_LFInst_3_n7,
         SubCellInst2_LFInst_13_LFInst_0_n15,
         SubCellInst2_LFInst_13_LFInst_0_n14,
         SubCellInst2_LFInst_13_LFInst_0_n13,
         SubCellInst2_LFInst_13_LFInst_0_n12,
         SubCellInst2_LFInst_13_LFInst_0_n11,
         SubCellInst2_LFInst_13_LFInst_1_n9,
         SubCellInst2_LFInst_13_LFInst_1_n8,
         SubCellInst2_LFInst_13_LFInst_1_n7,
         SubCellInst2_LFInst_13_LFInst_2_n18,
         SubCellInst2_LFInst_13_LFInst_2_n17,
         SubCellInst2_LFInst_13_LFInst_2_n16,
         SubCellInst2_LFInst_13_LFInst_2_n15,
         SubCellInst2_LFInst_13_LFInst_2_n14,
         SubCellInst2_LFInst_13_LFInst_3_n9,
         SubCellInst2_LFInst_13_LFInst_3_n8,
         SubCellInst2_LFInst_13_LFInst_3_n7,
         SubCellInst2_LFInst_14_LFInst_0_n15,
         SubCellInst2_LFInst_14_LFInst_0_n14,
         SubCellInst2_LFInst_14_LFInst_0_n13,
         SubCellInst2_LFInst_14_LFInst_0_n12,
         SubCellInst2_LFInst_14_LFInst_0_n11,
         SubCellInst2_LFInst_14_LFInst_1_n9,
         SubCellInst2_LFInst_14_LFInst_1_n8,
         SubCellInst2_LFInst_14_LFInst_1_n7,
         SubCellInst2_LFInst_14_LFInst_2_n18,
         SubCellInst2_LFInst_14_LFInst_2_n17,
         SubCellInst2_LFInst_14_LFInst_2_n16,
         SubCellInst2_LFInst_14_LFInst_2_n15,
         SubCellInst2_LFInst_14_LFInst_2_n14,
         SubCellInst2_LFInst_14_LFInst_3_n9,
         SubCellInst2_LFInst_14_LFInst_3_n8,
         SubCellInst2_LFInst_14_LFInst_3_n7,
         SubCellInst2_LFInst_15_LFInst_0_n15,
         SubCellInst2_LFInst_15_LFInst_0_n14,
         SubCellInst2_LFInst_15_LFInst_0_n13,
         SubCellInst2_LFInst_15_LFInst_0_n12,
         SubCellInst2_LFInst_15_LFInst_0_n11,
         SubCellInst2_LFInst_15_LFInst_1_n9,
         SubCellInst2_LFInst_15_LFInst_1_n8,
         SubCellInst2_LFInst_15_LFInst_1_n7,
         SubCellInst2_LFInst_15_LFInst_2_n18,
         SubCellInst2_LFInst_15_LFInst_2_n17,
         SubCellInst2_LFInst_15_LFInst_2_n16,
         SubCellInst2_LFInst_15_LFInst_2_n15,
         SubCellInst2_LFInst_15_LFInst_2_n14,
         SubCellInst2_LFInst_15_LFInst_3_n9,
         SubCellInst2_LFInst_15_LFInst_3_n8,
         SubCellInst2_LFInst_15_LFInst_3_n7,
         Red_PlaintextInst_LFInst_0_LFInst_0_n6,
         Red_PlaintextInst_LFInst_0_LFInst_0_n5,
         Red_PlaintextInst_LFInst_1_LFInst_0_n6,
         Red_PlaintextInst_LFInst_1_LFInst_0_n5,
         Red_PlaintextInst_LFInst_2_LFInst_0_n6,
         Red_PlaintextInst_LFInst_2_LFInst_0_n5,
         Red_PlaintextInst_LFInst_3_LFInst_0_n6,
         Red_PlaintextInst_LFInst_3_LFInst_0_n5,
         Red_PlaintextInst_LFInst_4_LFInst_0_n6,
         Red_PlaintextInst_LFInst_4_LFInst_0_n5,
         Red_PlaintextInst_LFInst_5_LFInst_0_n6,
         Red_PlaintextInst_LFInst_5_LFInst_0_n5,
         Red_PlaintextInst_LFInst_6_LFInst_0_n6,
         Red_PlaintextInst_LFInst_6_LFInst_0_n5,
         Red_PlaintextInst_LFInst_7_LFInst_0_n6,
         Red_PlaintextInst_LFInst_7_LFInst_0_n5,
         Red_PlaintextInst_LFInst_8_LFInst_0_n6,
         Red_PlaintextInst_LFInst_8_LFInst_0_n5,
         Red_PlaintextInst_LFInst_9_LFInst_0_n6,
         Red_PlaintextInst_LFInst_9_LFInst_0_n5,
         Red_PlaintextInst_LFInst_10_LFInst_0_n6,
         Red_PlaintextInst_LFInst_10_LFInst_0_n5,
         Red_PlaintextInst_LFInst_11_LFInst_0_n6,
         Red_PlaintextInst_LFInst_11_LFInst_0_n5,
         Red_PlaintextInst_LFInst_12_LFInst_0_n6,
         Red_PlaintextInst_LFInst_12_LFInst_0_n5,
         Red_PlaintextInst_LFInst_13_LFInst_0_n6,
         Red_PlaintextInst_LFInst_13_LFInst_0_n5,
         Red_PlaintextInst_LFInst_14_LFInst_0_n6,
         Red_PlaintextInst_LFInst_14_LFInst_0_n5,
         Red_PlaintextInst_LFInst_15_LFInst_0_n6,
         Red_PlaintextInst_LFInst_15_LFInst_0_n5, Red_MCInst_XOR_r0_Inst_0_n5,
         Red_MCInst_XOR_r0_Inst_1_n5, Red_MCInst_XOR_r0_Inst_2_n5,
         Red_MCInst_XOR_r0_Inst_3_n5, Red_SubCellInst_LFInst_0_LFInst_0_n22,
         Red_SubCellInst_LFInst_0_LFInst_0_n21,
         Red_SubCellInst_LFInst_0_LFInst_0_n20,
         Red_SubCellInst_LFInst_0_LFInst_0_n19,
         Red_SubCellInst_LFInst_0_LFInst_0_n18,
         Red_SubCellInst_LFInst_0_LFInst_0_n17,
         Red_SubCellInst_LFInst_0_LFInst_0_n16,
         Red_SubCellInst_LFInst_0_LFInst_0_n15,
         Red_SubCellInst_LFInst_0_LFInst_0_n14,
         Red_SubCellInst_LFInst_1_LFInst_0_n22,
         Red_SubCellInst_LFInst_1_LFInst_0_n21,
         Red_SubCellInst_LFInst_1_LFInst_0_n20,
         Red_SubCellInst_LFInst_1_LFInst_0_n19,
         Red_SubCellInst_LFInst_1_LFInst_0_n18,
         Red_SubCellInst_LFInst_1_LFInst_0_n17,
         Red_SubCellInst_LFInst_1_LFInst_0_n16,
         Red_SubCellInst_LFInst_1_LFInst_0_n15,
         Red_SubCellInst_LFInst_1_LFInst_0_n14,
         Red_SubCellInst_LFInst_2_LFInst_0_n22,
         Red_SubCellInst_LFInst_2_LFInst_0_n21,
         Red_SubCellInst_LFInst_2_LFInst_0_n20,
         Red_SubCellInst_LFInst_2_LFInst_0_n19,
         Red_SubCellInst_LFInst_2_LFInst_0_n18,
         Red_SubCellInst_LFInst_2_LFInst_0_n17,
         Red_SubCellInst_LFInst_2_LFInst_0_n16,
         Red_SubCellInst_LFInst_2_LFInst_0_n15,
         Red_SubCellInst_LFInst_2_LFInst_0_n14,
         Red_SubCellInst_LFInst_3_LFInst_0_n22,
         Red_SubCellInst_LFInst_3_LFInst_0_n21,
         Red_SubCellInst_LFInst_3_LFInst_0_n20,
         Red_SubCellInst_LFInst_3_LFInst_0_n19,
         Red_SubCellInst_LFInst_3_LFInst_0_n18,
         Red_SubCellInst_LFInst_3_LFInst_0_n17,
         Red_SubCellInst_LFInst_3_LFInst_0_n16,
         Red_SubCellInst_LFInst_3_LFInst_0_n15,
         Red_SubCellInst_LFInst_3_LFInst_0_n14,
         Red_SubCellInst_LFInst_4_LFInst_0_n19,
         Red_SubCellInst_LFInst_4_LFInst_0_n18,
         Red_SubCellInst_LFInst_4_LFInst_0_n17,
         Red_SubCellInst_LFInst_4_LFInst_0_n16,
         Red_SubCellInst_LFInst_4_LFInst_0_n15,
         Red_SubCellInst_LFInst_4_LFInst_0_n14,
         Red_SubCellInst_LFInst_5_LFInst_0_n19,
         Red_SubCellInst_LFInst_5_LFInst_0_n18,
         Red_SubCellInst_LFInst_5_LFInst_0_n17,
         Red_SubCellInst_LFInst_5_LFInst_0_n16,
         Red_SubCellInst_LFInst_5_LFInst_0_n15,
         Red_SubCellInst_LFInst_5_LFInst_0_n14,
         Red_SubCellInst_LFInst_6_LFInst_0_n19,
         Red_SubCellInst_LFInst_6_LFInst_0_n18,
         Red_SubCellInst_LFInst_6_LFInst_0_n17,
         Red_SubCellInst_LFInst_6_LFInst_0_n16,
         Red_SubCellInst_LFInst_6_LFInst_0_n15,
         Red_SubCellInst_LFInst_6_LFInst_0_n14,
         Red_SubCellInst_LFInst_7_LFInst_0_n19,
         Red_SubCellInst_LFInst_7_LFInst_0_n18,
         Red_SubCellInst_LFInst_7_LFInst_0_n17,
         Red_SubCellInst_LFInst_7_LFInst_0_n16,
         Red_SubCellInst_LFInst_7_LFInst_0_n15,
         Red_SubCellInst_LFInst_7_LFInst_0_n14,
         Red_SubCellInst_LFInst_8_LFInst_0_n22,
         Red_SubCellInst_LFInst_8_LFInst_0_n21,
         Red_SubCellInst_LFInst_8_LFInst_0_n20,
         Red_SubCellInst_LFInst_8_LFInst_0_n19,
         Red_SubCellInst_LFInst_8_LFInst_0_n18,
         Red_SubCellInst_LFInst_8_LFInst_0_n17,
         Red_SubCellInst_LFInst_8_LFInst_0_n16,
         Red_SubCellInst_LFInst_8_LFInst_0_n15,
         Red_SubCellInst_LFInst_8_LFInst_0_n14,
         Red_SubCellInst_LFInst_9_LFInst_0_n22,
         Red_SubCellInst_LFInst_9_LFInst_0_n21,
         Red_SubCellInst_LFInst_9_LFInst_0_n20,
         Red_SubCellInst_LFInst_9_LFInst_0_n19,
         Red_SubCellInst_LFInst_9_LFInst_0_n18,
         Red_SubCellInst_LFInst_9_LFInst_0_n17,
         Red_SubCellInst_LFInst_9_LFInst_0_n16,
         Red_SubCellInst_LFInst_9_LFInst_0_n15,
         Red_SubCellInst_LFInst_9_LFInst_0_n14,
         Red_SubCellInst_LFInst_10_LFInst_0_n22,
         Red_SubCellInst_LFInst_10_LFInst_0_n21,
         Red_SubCellInst_LFInst_10_LFInst_0_n20,
         Red_SubCellInst_LFInst_10_LFInst_0_n19,
         Red_SubCellInst_LFInst_10_LFInst_0_n18,
         Red_SubCellInst_LFInst_10_LFInst_0_n17,
         Red_SubCellInst_LFInst_10_LFInst_0_n16,
         Red_SubCellInst_LFInst_10_LFInst_0_n15,
         Red_SubCellInst_LFInst_10_LFInst_0_n14,
         Red_SubCellInst_LFInst_11_LFInst_0_n22,
         Red_SubCellInst_LFInst_11_LFInst_0_n21,
         Red_SubCellInst_LFInst_11_LFInst_0_n20,
         Red_SubCellInst_LFInst_11_LFInst_0_n19,
         Red_SubCellInst_LFInst_11_LFInst_0_n18,
         Red_SubCellInst_LFInst_11_LFInst_0_n17,
         Red_SubCellInst_LFInst_11_LFInst_0_n16,
         Red_SubCellInst_LFInst_11_LFInst_0_n15,
         Red_SubCellInst_LFInst_11_LFInst_0_n14,
         Red_SubCellInst_LFInst_12_LFInst_0_n22,
         Red_SubCellInst_LFInst_12_LFInst_0_n21,
         Red_SubCellInst_LFInst_12_LFInst_0_n20,
         Red_SubCellInst_LFInst_12_LFInst_0_n19,
         Red_SubCellInst_LFInst_12_LFInst_0_n18,
         Red_SubCellInst_LFInst_12_LFInst_0_n17,
         Red_SubCellInst_LFInst_12_LFInst_0_n16,
         Red_SubCellInst_LFInst_12_LFInst_0_n15,
         Red_SubCellInst_LFInst_12_LFInst_0_n14,
         Red_SubCellInst_LFInst_13_LFInst_0_n22,
         Red_SubCellInst_LFInst_13_LFInst_0_n21,
         Red_SubCellInst_LFInst_13_LFInst_0_n20,
         Red_SubCellInst_LFInst_13_LFInst_0_n19,
         Red_SubCellInst_LFInst_13_LFInst_0_n18,
         Red_SubCellInst_LFInst_13_LFInst_0_n17,
         Red_SubCellInst_LFInst_13_LFInst_0_n16,
         Red_SubCellInst_LFInst_13_LFInst_0_n15,
         Red_SubCellInst_LFInst_13_LFInst_0_n14,
         Red_SubCellInst_LFInst_14_LFInst_0_n22,
         Red_SubCellInst_LFInst_14_LFInst_0_n21,
         Red_SubCellInst_LFInst_14_LFInst_0_n20,
         Red_SubCellInst_LFInst_14_LFInst_0_n19,
         Red_SubCellInst_LFInst_14_LFInst_0_n18,
         Red_SubCellInst_LFInst_14_LFInst_0_n17,
         Red_SubCellInst_LFInst_14_LFInst_0_n16,
         Red_SubCellInst_LFInst_14_LFInst_0_n15,
         Red_SubCellInst_LFInst_14_LFInst_0_n14,
         Red_SubCellInst_LFInst_15_LFInst_0_n22,
         Red_SubCellInst_LFInst_15_LFInst_0_n21,
         Red_SubCellInst_LFInst_15_LFInst_0_n20,
         Red_SubCellInst_LFInst_15_LFInst_0_n19,
         Red_SubCellInst_LFInst_15_LFInst_0_n18,
         Red_SubCellInst_LFInst_15_LFInst_0_n17,
         Red_SubCellInst_LFInst_15_LFInst_0_n16,
         Red_SubCellInst_LFInst_15_LFInst_0_n15,
         Red_SubCellInst_LFInst_15_LFInst_0_n14, Red_MCInst2_XOR_r0_Inst_0_n5,
         Red_MCInst2_XOR_r0_Inst_1_n5, Red_MCInst2_XOR_r0_Inst_2_n5,
         Red_MCInst2_XOR_r0_Inst_3_n5, Red_SubCellInst2_LFInst_0_LFInst_0_n17,
         Red_SubCellInst2_LFInst_0_LFInst_0_n16,
         Red_SubCellInst2_LFInst_0_LFInst_0_n15,
         Red_SubCellInst2_LFInst_0_LFInst_0_n14,
         Red_SubCellInst2_LFInst_1_LFInst_0_n21,
         Red_SubCellInst2_LFInst_1_LFInst_0_n20,
         Red_SubCellInst2_LFInst_1_LFInst_0_n19,
         Red_SubCellInst2_LFInst_1_LFInst_0_n18,
         Red_SubCellInst2_LFInst_1_LFInst_0_n17,
         Red_SubCellInst2_LFInst_1_LFInst_0_n16,
         Red_SubCellInst2_LFInst_2_LFInst_0_n17,
         Red_SubCellInst2_LFInst_2_LFInst_0_n16,
         Red_SubCellInst2_LFInst_2_LFInst_0_n15,
         Red_SubCellInst2_LFInst_2_LFInst_0_n14,
         Red_SubCellInst2_LFInst_3_LFInst_0_n17,
         Red_SubCellInst2_LFInst_3_LFInst_0_n16,
         Red_SubCellInst2_LFInst_3_LFInst_0_n15,
         Red_SubCellInst2_LFInst_3_LFInst_0_n14,
         Red_SubCellInst2_LFInst_4_LFInst_0_n22,
         Red_SubCellInst2_LFInst_4_LFInst_0_n21,
         Red_SubCellInst2_LFInst_4_LFInst_0_n20,
         Red_SubCellInst2_LFInst_4_LFInst_0_n19,
         Red_SubCellInst2_LFInst_4_LFInst_0_n18,
         Red_SubCellInst2_LFInst_4_LFInst_0_n17,
         Red_SubCellInst2_LFInst_4_LFInst_0_n16,
         Red_SubCellInst2_LFInst_4_LFInst_0_n15,
         Red_SubCellInst2_LFInst_4_LFInst_0_n14,
         Red_SubCellInst2_LFInst_5_LFInst_0_n17,
         Red_SubCellInst2_LFInst_5_LFInst_0_n16,
         Red_SubCellInst2_LFInst_5_LFInst_0_n15,
         Red_SubCellInst2_LFInst_5_LFInst_0_n14,
         Red_SubCellInst2_LFInst_6_LFInst_0_n22,
         Red_SubCellInst2_LFInst_6_LFInst_0_n21,
         Red_SubCellInst2_LFInst_6_LFInst_0_n20,
         Red_SubCellInst2_LFInst_6_LFInst_0_n19,
         Red_SubCellInst2_LFInst_6_LFInst_0_n18,
         Red_SubCellInst2_LFInst_6_LFInst_0_n17,
         Red_SubCellInst2_LFInst_6_LFInst_0_n16,
         Red_SubCellInst2_LFInst_6_LFInst_0_n15,
         Red_SubCellInst2_LFInst_6_LFInst_0_n14,
         Red_SubCellInst2_LFInst_7_LFInst_0_n22,
         Red_SubCellInst2_LFInst_7_LFInst_0_n21,
         Red_SubCellInst2_LFInst_7_LFInst_0_n20,
         Red_SubCellInst2_LFInst_7_LFInst_0_n19,
         Red_SubCellInst2_LFInst_7_LFInst_0_n18,
         Red_SubCellInst2_LFInst_7_LFInst_0_n17,
         Red_SubCellInst2_LFInst_7_LFInst_0_n16,
         Red_SubCellInst2_LFInst_7_LFInst_0_n15,
         Red_SubCellInst2_LFInst_7_LFInst_0_n14,
         Red_SubCellInst2_LFInst_8_LFInst_0_n17,
         Red_SubCellInst2_LFInst_8_LFInst_0_n16,
         Red_SubCellInst2_LFInst_8_LFInst_0_n15,
         Red_SubCellInst2_LFInst_8_LFInst_0_n14,
         Red_SubCellInst2_LFInst_9_LFInst_0_n17,
         Red_SubCellInst2_LFInst_9_LFInst_0_n16,
         Red_SubCellInst2_LFInst_9_LFInst_0_n15,
         Red_SubCellInst2_LFInst_9_LFInst_0_n14,
         Red_SubCellInst2_LFInst_10_LFInst_0_n22,
         Red_SubCellInst2_LFInst_10_LFInst_0_n21,
         Red_SubCellInst2_LFInst_10_LFInst_0_n20,
         Red_SubCellInst2_LFInst_10_LFInst_0_n19,
         Red_SubCellInst2_LFInst_10_LFInst_0_n18,
         Red_SubCellInst2_LFInst_10_LFInst_0_n17,
         Red_SubCellInst2_LFInst_10_LFInst_0_n16,
         Red_SubCellInst2_LFInst_10_LFInst_0_n15,
         Red_SubCellInst2_LFInst_10_LFInst_0_n14,
         Red_SubCellInst2_LFInst_11_LFInst_0_n17,
         Red_SubCellInst2_LFInst_11_LFInst_0_n16,
         Red_SubCellInst2_LFInst_11_LFInst_0_n15,
         Red_SubCellInst2_LFInst_11_LFInst_0_n14,
         Red_SubCellInst2_LFInst_12_LFInst_0_n21,
         Red_SubCellInst2_LFInst_12_LFInst_0_n20,
         Red_SubCellInst2_LFInst_12_LFInst_0_n19,
         Red_SubCellInst2_LFInst_12_LFInst_0_n18,
         Red_SubCellInst2_LFInst_12_LFInst_0_n17,
         Red_SubCellInst2_LFInst_12_LFInst_0_n16,
         Red_SubCellInst2_LFInst_13_LFInst_0_n17,
         Red_SubCellInst2_LFInst_13_LFInst_0_n16,
         Red_SubCellInst2_LFInst_13_LFInst_0_n15,
         Red_SubCellInst2_LFInst_13_LFInst_0_n14,
         Red_SubCellInst2_LFInst_14_LFInst_0_n21,
         Red_SubCellInst2_LFInst_14_LFInst_0_n20,
         Red_SubCellInst2_LFInst_14_LFInst_0_n19,
         Red_SubCellInst2_LFInst_14_LFInst_0_n18,
         Red_SubCellInst2_LFInst_14_LFInst_0_n17,
         Red_SubCellInst2_LFInst_14_LFInst_0_n16,
         Red_SubCellInst2_LFInst_15_LFInst_0_n21,
         Red_SubCellInst2_LFInst_15_LFInst_0_n20,
         Red_SubCellInst2_LFInst_15_LFInst_0_n19,
         Red_SubCellInst2_LFInst_15_LFInst_0_n18,
         Red_SubCellInst2_LFInst_15_LFInst_0_n17,
         Red_SubCellInst2_LFInst_15_LFInst_0_n16,
         Red_K0Inst_LFInst_0_LFInst_0_n6, Red_K0Inst_LFInst_0_LFInst_0_n5,
         Red_K0Inst_LFInst_1_LFInst_0_n6, Red_K0Inst_LFInst_1_LFInst_0_n5,
         Red_K0Inst_LFInst_2_LFInst_0_n6, Red_K0Inst_LFInst_2_LFInst_0_n5,
         Red_K0Inst_LFInst_3_LFInst_0_n6, Red_K0Inst_LFInst_3_LFInst_0_n5,
         Red_K0Inst_LFInst_4_LFInst_0_n6, Red_K0Inst_LFInst_4_LFInst_0_n5,
         Red_K0Inst_LFInst_5_LFInst_0_n6, Red_K0Inst_LFInst_5_LFInst_0_n5,
         Red_K0Inst_LFInst_6_LFInst_0_n6, Red_K0Inst_LFInst_6_LFInst_0_n5,
         Red_K0Inst_LFInst_7_LFInst_0_n6, Red_K0Inst_LFInst_7_LFInst_0_n5,
         Red_K0Inst_LFInst_8_LFInst_0_n6, Red_K0Inst_LFInst_8_LFInst_0_n5,
         Red_K0Inst_LFInst_9_LFInst_0_n6, Red_K0Inst_LFInst_9_LFInst_0_n5,
         Red_K0Inst_LFInst_10_LFInst_0_n6, Red_K0Inst_LFInst_10_LFInst_0_n5,
         Red_K0Inst_LFInst_11_LFInst_0_n6, Red_K0Inst_LFInst_11_LFInst_0_n5,
         Red_K0Inst_LFInst_12_LFInst_0_n6, Red_K0Inst_LFInst_12_LFInst_0_n5,
         Red_K0Inst_LFInst_13_LFInst_0_n6, Red_K0Inst_LFInst_13_LFInst_0_n5,
         Red_K0Inst_LFInst_14_LFInst_0_n6, Red_K0Inst_LFInst_14_LFInst_0_n5,
         Red_K0Inst_LFInst_15_LFInst_0_n6, Red_K0Inst_LFInst_15_LFInst_0_n5,
         Red_K1Inst_LFInst_0_LFInst_0_n6, Red_K1Inst_LFInst_0_LFInst_0_n5,
         Red_K1Inst_LFInst_1_LFInst_0_n6, Red_K1Inst_LFInst_1_LFInst_0_n5,
         Red_K1Inst_LFInst_2_LFInst_0_n6, Red_K1Inst_LFInst_2_LFInst_0_n5,
         Red_K1Inst_LFInst_3_LFInst_0_n6, Red_K1Inst_LFInst_3_LFInst_0_n5,
         Red_K1Inst_LFInst_4_LFInst_0_n6, Red_K1Inst_LFInst_4_LFInst_0_n5,
         Red_K1Inst_LFInst_5_LFInst_0_n6, Red_K1Inst_LFInst_5_LFInst_0_n5,
         Red_K1Inst_LFInst_6_LFInst_0_n6, Red_K1Inst_LFInst_6_LFInst_0_n5,
         Red_K1Inst_LFInst_7_LFInst_0_n6, Red_K1Inst_LFInst_7_LFInst_0_n5,
         Red_K1Inst_LFInst_8_LFInst_0_n6, Red_K1Inst_LFInst_8_LFInst_0_n5,
         Red_K1Inst_LFInst_9_LFInst_0_n6, Red_K1Inst_LFInst_9_LFInst_0_n5,
         Red_K1Inst_LFInst_10_LFInst_0_n6, Red_K1Inst_LFInst_10_LFInst_0_n5,
         Red_K1Inst_LFInst_11_LFInst_0_n6, Red_K1Inst_LFInst_11_LFInst_0_n5,
         Red_K1Inst_LFInst_12_LFInst_0_n6, Red_K1Inst_LFInst_12_LFInst_0_n5,
         Red_K1Inst_LFInst_13_LFInst_0_n6, Red_K1Inst_LFInst_13_LFInst_0_n5,
         Red_K1Inst_LFInst_14_LFInst_0_n6, Red_K1Inst_LFInst_14_LFInst_0_n5,
         Red_K1Inst_LFInst_15_LFInst_0_n6, Red_K1Inst_LFInst_15_LFInst_0_n5,
         Red_ToCheckInst_LFInst_0_LFInst_0_n6,
         Red_ToCheckInst_LFInst_0_LFInst_0_n5,
         Red_ToCheckInst_LFInst_1_LFInst_0_n6,
         Red_ToCheckInst_LFInst_1_LFInst_0_n5,
         Red_ToCheckInst_LFInst_2_LFInst_0_n6,
         Red_ToCheckInst_LFInst_2_LFInst_0_n5,
         Red_ToCheckInst_LFInst_3_LFInst_0_n6,
         Red_ToCheckInst_LFInst_3_LFInst_0_n5,
         Red_ToCheckInst_LFInst_4_LFInst_0_n6,
         Red_ToCheckInst_LFInst_4_LFInst_0_n5,
         Red_ToCheckInst_LFInst_5_LFInst_0_n6,
         Red_ToCheckInst_LFInst_5_LFInst_0_n5,
         Red_ToCheckInst_LFInst_6_LFInst_0_n6,
         Red_ToCheckInst_LFInst_6_LFInst_0_n5,
         Red_ToCheckInst_LFInst_7_LFInst_0_n6,
         Red_ToCheckInst_LFInst_7_LFInst_0_n5,
         Red_ToCheckInst_LFInst_8_LFInst_0_n6,
         Red_ToCheckInst_LFInst_8_LFInst_0_n5,
         Red_ToCheckInst_LFInst_9_LFInst_0_n6,
         Red_ToCheckInst_LFInst_9_LFInst_0_n5,
         Red_ToCheckInst_LFInst_10_LFInst_0_n6,
         Red_ToCheckInst_LFInst_10_LFInst_0_n5,
         Red_ToCheckInst_LFInst_11_LFInst_0_n6,
         Red_ToCheckInst_LFInst_11_LFInst_0_n5,
         Red_ToCheckInst_LFInst_12_LFInst_0_n6,
         Red_ToCheckInst_LFInst_12_LFInst_0_n5,
         Red_ToCheckInst_LFInst_13_LFInst_0_n6,
         Red_ToCheckInst_LFInst_13_LFInst_0_n5,
         Red_ToCheckInst_LFInst_14_LFInst_0_n6,
         Red_ToCheckInst_LFInst_14_LFInst_0_n5,
         Red_ToCheckInst_LFInst_15_LFInst_0_n6,
         Red_ToCheckInst_LFInst_15_LFInst_0_n5,
         Red_ToCheckInst_LFInst_16_LFInst_0_n6,
         Red_ToCheckInst_LFInst_16_LFInst_0_n5,
         Red_ToCheckInst_LFInst_17_LFInst_0_n6,
         Red_ToCheckInst_LFInst_17_LFInst_0_n5,
         Red_ToCheckInst_LFInst_18_LFInst_0_n6,
         Red_ToCheckInst_LFInst_18_LFInst_0_n5,
         Red_ToCheckInst_LFInst_19_LFInst_0_n6,
         Red_ToCheckInst_LFInst_19_LFInst_0_n5,
         Red_ToCheckInst_LFInst_20_LFInst_0_n6,
         Red_ToCheckInst_LFInst_20_LFInst_0_n5,
         Red_ToCheckInst_LFInst_21_LFInst_0_n6,
         Red_ToCheckInst_LFInst_21_LFInst_0_n5,
         Red_ToCheckInst_LFInst_22_LFInst_0_n6,
         Red_ToCheckInst_LFInst_22_LFInst_0_n5,
         Red_ToCheckInst_LFInst_23_LFInst_0_n6,
         Red_ToCheckInst_LFInst_23_LFInst_0_n5,
         Red_ToCheckInst_LFInst_24_LFInst_0_n6,
         Red_ToCheckInst_LFInst_24_LFInst_0_n5,
         Red_ToCheckInst_LFInst_25_LFInst_0_n6,
         Red_ToCheckInst_LFInst_25_LFInst_0_n5,
         Red_ToCheckInst_LFInst_26_LFInst_0_n6,
         Red_ToCheckInst_LFInst_26_LFInst_0_n5,
         Red_ToCheckInst_LFInst_27_LFInst_0_n6,
         Red_ToCheckInst_LFInst_27_LFInst_0_n5,
         Red_ToCheckInst_LFInst_28_LFInst_0_n6,
         Red_ToCheckInst_LFInst_28_LFInst_0_n5,
         Red_ToCheckInst_LFInst_29_LFInst_0_n6,
         Red_ToCheckInst_LFInst_29_LFInst_0_n5,
         Red_ToCheckInst_LFInst_30_LFInst_0_n6,
         Red_ToCheckInst_LFInst_30_LFInst_0_n5,
         Red_ToCheckInst_LFInst_31_LFInst_0_n6,
         Red_ToCheckInst_LFInst_31_LFInst_0_n5,
         Red_ToCheckInst_LFInst_32_LFInst_0_n6,
         Red_ToCheckInst_LFInst_32_LFInst_0_n5,
         Red_ToCheckInst_LFInst_33_LFInst_0_n6,
         Red_ToCheckInst_LFInst_33_LFInst_0_n5,
         Red_ToCheckInst_LFInst_34_LFInst_0_n6,
         Red_ToCheckInst_LFInst_34_LFInst_0_n5,
         Red_ToCheckInst_LFInst_35_LFInst_0_n6,
         Red_ToCheckInst_LFInst_35_LFInst_0_n5,
         Red_ToCheckInst_LFInst_36_LFInst_0_n6,
         Red_ToCheckInst_LFInst_36_LFInst_0_n5,
         Red_ToCheckInst_LFInst_37_LFInst_0_n6,
         Red_ToCheckInst_LFInst_37_LFInst_0_n5,
         Red_ToCheckInst_LFInst_38_LFInst_0_n6,
         Red_ToCheckInst_LFInst_38_LFInst_0_n5,
         Red_ToCheckInst_LFInst_39_LFInst_0_n6,
         Red_ToCheckInst_LFInst_39_LFInst_0_n5,
         Red_ToCheckInst_LFInst_40_LFInst_0_n6,
         Red_ToCheckInst_LFInst_40_LFInst_0_n5,
         Red_ToCheckInst_LFInst_41_LFInst_0_n6,
         Red_ToCheckInst_LFInst_41_LFInst_0_n5,
         Red_ToCheckInst_LFInst_42_LFInst_0_n6,
         Red_ToCheckInst_LFInst_42_LFInst_0_n5,
         Red_ToCheckInst_LFInst_43_LFInst_0_n6,
         Red_ToCheckInst_LFInst_43_LFInst_0_n5,
         Red_ToCheckInst_LFInst_44_LFInst_0_n6,
         Red_ToCheckInst_LFInst_44_LFInst_0_n5,
         Red_ToCheckInst_LFInst_45_LFInst_0_n6,
         Red_ToCheckInst_LFInst_45_LFInst_0_n5,
         Red_ToCheckInst_LFInst_46_LFInst_0_n6,
         Red_ToCheckInst_LFInst_46_LFInst_0_n5,
         Red_ToCheckInst_LFInst_47_LFInst_0_n6,
         Red_ToCheckInst_LFInst_47_LFInst_0_n5,
         Red_ToCheckInst_LFInst_48_LFInst_0_n6,
         Red_ToCheckInst_LFInst_48_LFInst_0_n5,
         Red_ToCheckInst_LFInst_49_LFInst_0_n6,
         Red_ToCheckInst_LFInst_49_LFInst_0_n5,
         Red_ToCheckInst_LFInst_50_LFInst_0_n6,
         Red_ToCheckInst_LFInst_50_LFInst_0_n5,
         Red_ToCheckInst_LFInst_51_LFInst_0_n6,
         Red_ToCheckInst_LFInst_51_LFInst_0_n5,
         Red_ToCheckInst_LFInst_52_LFInst_0_n6,
         Red_ToCheckInst_LFInst_52_LFInst_0_n5,
         Red_ToCheckInst_LFInst_53_LFInst_0_n6,
         Red_ToCheckInst_LFInst_53_LFInst_0_n5,
         Red_ToCheckInst_LFInst_54_LFInst_0_n6,
         Red_ToCheckInst_LFInst_54_LFInst_0_n5,
         Red_ToCheckInst_LFInst_55_LFInst_0_n6,
         Red_ToCheckInst_LFInst_55_LFInst_0_n5,
         Red_ToCheckInst_LFInst_56_LFInst_0_n6,
         Red_ToCheckInst_LFInst_56_LFInst_0_n5,
         Red_ToCheckInst_LFInst_57_LFInst_0_n6,
         Red_ToCheckInst_LFInst_57_LFInst_0_n5,
         Red_ToCheckInst_LFInst_58_LFInst_0_n6,
         Red_ToCheckInst_LFInst_58_LFInst_0_n5,
         Red_ToCheckInst_LFInst_59_LFInst_0_n6,
         Red_ToCheckInst_LFInst_59_LFInst_0_n5,
         Red_ToCheckInst_LFInst_60_LFInst_0_n6,
         Red_ToCheckInst_LFInst_60_LFInst_0_n5,
         Red_ToCheckInst_LFInst_61_LFInst_0_n6,
         Red_ToCheckInst_LFInst_61_LFInst_0_n5,
         Red_ToCheckInst_LFInst_62_LFInst_0_n6,
         Red_ToCheckInst_LFInst_62_LFInst_0_n5,
         Red_ToCheckInst_LFInst_63_LFInst_0_n6,
         Red_ToCheckInst_LFInst_63_LFInst_0_n5,
         Red_ToCheckInst_LFInst_64_LFInst_0_n6,
         Red_ToCheckInst_LFInst_64_LFInst_0_n5,
         Red_ToCheckInst_LFInst_65_LFInst_0_n6,
         Red_ToCheckInst_LFInst_65_LFInst_0_n5,
         Red_ToCheckInst_LFInst_66_LFInst_0_n6,
         Red_ToCheckInst_LFInst_66_LFInst_0_n5,
         Red_ToCheckInst_LFInst_67_LFInst_0_n6,
         Red_ToCheckInst_LFInst_67_LFInst_0_n5,
         Red_ToCheckInst_LFInst_68_LFInst_0_n6,
         Red_ToCheckInst_LFInst_68_LFInst_0_n5,
         Red_ToCheckInst_LFInst_69_LFInst_0_n6,
         Red_ToCheckInst_LFInst_69_LFInst_0_n5,
         Red_ToCheckInst_LFInst_70_LFInst_0_n6,
         Red_ToCheckInst_LFInst_70_LFInst_0_n5,
         Red_ToCheckInst_LFInst_71_LFInst_0_n6,
         Red_ToCheckInst_LFInst_71_LFInst_0_n5,
         Red_ToCheckInst_LFInst_72_LFInst_0_n6,
         Red_ToCheckInst_LFInst_72_LFInst_0_n5,
         Red_ToCheckInst_LFInst_73_LFInst_0_n6,
         Red_ToCheckInst_LFInst_73_LFInst_0_n5,
         Red_ToCheckInst_LFInst_74_LFInst_0_n6,
         Red_ToCheckInst_LFInst_74_LFInst_0_n5,
         Red_ToCheckInst_LFInst_75_LFInst_0_n6,
         Red_ToCheckInst_LFInst_75_LFInst_0_n5,
         Red_ToCheckInst_LFInst_76_LFInst_0_n6,
         Red_ToCheckInst_LFInst_76_LFInst_0_n5,
         Red_ToCheckInst_LFInst_77_LFInst_0_n6,
         Red_ToCheckInst_LFInst_77_LFInst_0_n5,
         Red_ToCheckInst_LFInst_78_LFInst_0_n6,
         Red_ToCheckInst_LFInst_78_LFInst_0_n5,
         Red_ToCheckInst_LFInst_79_LFInst_0_n6,
         Red_ToCheckInst_LFInst_79_LFInst_0_n5, Check1_CheckInst_0_n158,
         Check1_CheckInst_0_n157, Check1_CheckInst_0_n156,
         Check1_CheckInst_0_n155, Check1_CheckInst_0_n154,
         Check1_CheckInst_0_n153, Check1_CheckInst_0_n152,
         Check1_CheckInst_0_n151, Check1_CheckInst_0_n150,
         Check1_CheckInst_0_n149, Check1_CheckInst_0_n148,
         Check1_CheckInst_0_n147, Check1_CheckInst_0_n146,
         Check1_CheckInst_0_n145, Check1_CheckInst_0_n144,
         Check1_CheckInst_0_n143, Check1_CheckInst_0_n142,
         Check1_CheckInst_0_n141, Check1_CheckInst_0_n140,
         Check1_CheckInst_0_n139, Check1_CheckInst_0_n138,
         Check1_CheckInst_0_n137, Check1_CheckInst_0_n136,
         Check1_CheckInst_0_n135, Check1_CheckInst_0_n134,
         Check1_CheckInst_0_n133, Check1_CheckInst_0_n132,
         Check1_CheckInst_0_n131, Check1_CheckInst_0_n130,
         Check1_CheckInst_0_n129, Check1_CheckInst_0_n128,
         Check1_CheckInst_0_n127, Check1_CheckInst_0_n126,
         Check1_CheckInst_0_n125, Check1_CheckInst_0_n124,
         Check1_CheckInst_0_n123, Check1_CheckInst_0_n122,
         Check1_CheckInst_0_n121, Check1_CheckInst_0_n120,
         Check1_CheckInst_0_n119, Check1_CheckInst_0_n118,
         Check1_CheckInst_0_n117, Check1_CheckInst_0_n116,
         Check1_CheckInst_0_n115, Check1_CheckInst_0_n114,
         Check1_CheckInst_0_n113, Check1_CheckInst_0_n112,
         Check1_CheckInst_0_n111, Check1_CheckInst_0_n110,
         Check1_CheckInst_0_n109, Check1_CheckInst_0_n108,
         Check1_CheckInst_0_n107, Check1_CheckInst_0_n106,
         Check1_CheckInst_0_n105, Check1_CheckInst_0_n104,
         Check1_CheckInst_0_n103, Check1_CheckInst_0_n102,
         Check1_CheckInst_0_n101, Check1_CheckInst_0_n100,
         Check1_CheckInst_0_n99, Check1_CheckInst_0_n98,
         Check1_CheckInst_0_n97, Check1_CheckInst_0_n96,
         Check1_CheckInst_0_n95, Check1_CheckInst_0_n94,
         Check1_CheckInst_0_n93, Check1_CheckInst_0_n92,
         Check1_CheckInst_0_n91, Check1_CheckInst_0_n90,
         Check1_CheckInst_0_n89, Check1_CheckInst_0_n88,
         Check1_CheckInst_0_n87, Check1_CheckInst_0_n86,
         Check1_CheckInst_0_n85, Check1_CheckInst_0_n84,
         Check1_CheckInst_0_n83, Check1_CheckInst_0_n82,
         Check1_CheckInst_0_n81, Check1_CheckInst_0_n80,
         Check1_CheckInst_0_n79, Check1_CheckInst_0_n78,
         Check1_CheckInst_0_n77, Check1_CheckInst_0_n76,
         Check1_CheckInst_0_n75, Check1_CheckInst_0_n74,
         Check1_CheckInst_0_n73, Check1_CheckInst_0_n72,
         Check1_CheckInst_0_n71, Check1_CheckInst_0_n70,
         Check1_CheckInst_0_n69, Check1_CheckInst_0_n68,
         Check1_CheckInst_0_n67, Check1_CheckInst_0_n66,
         Check1_CheckInst_0_n65, Check1_CheckInst_0_n64,
         Check1_CheckInst_0_n63, Check1_CheckInst_0_n62,
         Check1_CheckInst_0_n61, Check1_CheckInst_0_n60,
         Check1_CheckInst_0_n59, Check1_CheckInst_0_n58,
         Check1_CheckInst_0_n57, Check1_CheckInst_0_n56,
         Check1_CheckInst_0_n55, Check1_CheckInst_0_n54,
         Check1_CheckInst_0_n53, Check1_CheckInst_0_n52,
         Check1_CheckInst_0_n51, Check1_CheckInst_0_n50,
         Check1_CheckInst_0_n49, Check1_CheckInst_0_n48,
         Check1_CheckInst_0_n47, Check1_CheckInst_0_n46,
         Check1_CheckInst_0_n45, Check1_CheckInst_0_n44,
         Check1_CheckInst_0_n43, Check1_CheckInst_0_n42,
         Check1_CheckInst_0_n41, Check1_CheckInst_0_n40,
         Check1_CheckInst_0_n39, Check1_CheckInst_0_n38,
         Check1_CheckInst_0_n37, Check1_CheckInst_0_n36,
         Check1_CheckInst_0_n35, Check1_CheckInst_0_n34,
         Check1_CheckInst_0_n33, Check1_CheckInst_0_n32,
         Check1_CheckInst_0_n31, Check1_CheckInst_0_n30,
         Check1_CheckInst_0_n29, Check1_CheckInst_0_n28,
         Check1_CheckInst_0_n27, Check1_CheckInst_0_n26,
         Check1_CheckInst_0_n25, Check1_CheckInst_0_n24,
         Check1_CheckInst_0_n23, Check1_CheckInst_0_n22,
         Check1_CheckInst_0_n21, Check1_CheckInst_0_n20,
         Check1_CheckInst_0_n19, Check1_CheckInst_0_n18,
         Check1_CheckInst_0_n17, Check1_CheckInst_0_n16,
         Check1_CheckInst_0_n15, Check1_CheckInst_0_n14,
         Check1_CheckInst_0_n13, Check1_CheckInst_0_n12,
         Check1_CheckInst_0_n11, Check1_CheckInst_0_n10, Check1_CheckInst_0_n9,
         Check1_CheckInst_0_n8, Check1_CheckInst_0_n7, Check1_CheckInst_0_n6,
         Check1_CheckInst_0_n5, Check1_CheckInst_0_n4, Check1_CheckInst_0_n3,
         Check1_CheckInst_0_n2, Check1_CheckInst_0_n1;
  wire   [63:0] AddRoundKeyOutput;
  wire   [63:0] PermutationOutput;
  wire   [63:32] SboxOut;
  wire   [63:0] MCOutput2;
  wire   [63:0] AddRoundKeyOutput2;
  wire   [63:0] PermutationOutput2;
  wire   [15:8] Red_Input;
  wire   [15:0] Red_MCOutput;
  wire   [15:0] Red_K0;
  wire   [15:0] Red_StateRegOutput;
  wire   [15:8] Red_SboxOut;
  wire   [15:0] Red_MCOutput2;
  wire   [15:0] Red_K1;
  wire   [15:0] Red_StateRegOutput2;
  wire   [15:0] Red_Feedback;
  wire   [31:0] Red_final;
  wire   [79:0] Red_SignaltoCheck;

  INV_X1 U4 ( .A(Error_0_), .ZN(ErrorFlag) );
  XNOR2_X1 MCInst_XOR_r0_Inst_0_U2 ( .A(MCInst_XOR_r0_Inst_0_n5), .B(Input[16]), .ZN(MCOutput_48_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_0_U1 ( .A(Input[0]), .B(Input[48]), .ZN(
        MCInst_XOR_r0_Inst_0_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_0_U1 ( .A(Input[32]), .B(Input[0]), .Z(
        MCOutput_32_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_1_U2 ( .A(MCInst_XOR_r0_Inst_1_n5), .B(Input[17]), .ZN(MCOutput_49_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_1_U1 ( .A(Input[1]), .B(Input[49]), .ZN(
        MCInst_XOR_r0_Inst_1_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_1_U1 ( .A(Input[33]), .B(Input[1]), .Z(
        MCOutput_33_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_2_U2 ( .A(MCInst_XOR_r0_Inst_2_n5), .B(Input[18]), .ZN(MCOutput_50_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_2_U1 ( .A(Input[2]), .B(Input[50]), .ZN(
        MCInst_XOR_r0_Inst_2_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_2_U1 ( .A(Input[34]), .B(Input[2]), .Z(
        MCOutput_34_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_3_U2 ( .A(MCInst_XOR_r0_Inst_3_n5), .B(Input[19]), .ZN(MCOutput_51_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_3_U1 ( .A(Input[3]), .B(Input[51]), .ZN(
        MCInst_XOR_r0_Inst_3_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_3_U1 ( .A(Input[35]), .B(Input[3]), .Z(
        MCOutput_35_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_4_U2 ( .A(MCInst_XOR_r0_Inst_4_n5), .B(Input[20]), .ZN(MCOutput_52_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_4_U1 ( .A(Input[4]), .B(Input[52]), .ZN(
        MCInst_XOR_r0_Inst_4_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_4_U1 ( .A(Input[36]), .B(Input[4]), .Z(
        MCOutput_36_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_5_U2 ( .A(MCInst_XOR_r0_Inst_5_n5), .B(Input[21]), .ZN(MCOutput_53_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_5_U1 ( .A(Input[5]), .B(Input[53]), .ZN(
        MCInst_XOR_r0_Inst_5_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_5_U1 ( .A(Input[37]), .B(Input[5]), .Z(
        MCOutput_37_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_6_U2 ( .A(MCInst_XOR_r0_Inst_6_n5), .B(Input[22]), .ZN(MCOutput_54_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_6_U1 ( .A(Input[6]), .B(Input[54]), .ZN(
        MCInst_XOR_r0_Inst_6_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_6_U1 ( .A(Input[38]), .B(Input[6]), .Z(
        MCOutput_38_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_7_U2 ( .A(MCInst_XOR_r0_Inst_7_n5), .B(Input[23]), .ZN(MCOutput_55_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_7_U1 ( .A(Input[7]), .B(Input[55]), .ZN(
        MCInst_XOR_r0_Inst_7_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_7_U1 ( .A(Input[39]), .B(Input[7]), .Z(
        MCOutput_39_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_8_U2 ( .A(MCInst_XOR_r0_Inst_8_n5), .B(Input[24]), .ZN(MCOutput_56_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_8_U1 ( .A(Input[8]), .B(Input[56]), .ZN(
        MCInst_XOR_r0_Inst_8_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_8_U1 ( .A(Input[40]), .B(Input[8]), .Z(
        MCOutput_40_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_9_U2 ( .A(MCInst_XOR_r0_Inst_9_n5), .B(Input[25]), .ZN(MCOutput_57_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_9_U1 ( .A(Input[9]), .B(Input[57]), .ZN(
        MCInst_XOR_r0_Inst_9_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_9_U1 ( .A(Input[41]), .B(Input[9]), .Z(
        MCOutput_41_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_10_U2 ( .A(MCInst_XOR_r0_Inst_10_n5), .B(
        Input[26]), .ZN(MCOutput_58_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_10_U1 ( .A(Input[10]), .B(Input[58]), .ZN(
        MCInst_XOR_r0_Inst_10_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_10_U1 ( .A(Input[42]), .B(Input[10]), .Z(
        MCOutput_42_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_11_U2 ( .A(MCInst_XOR_r0_Inst_11_n5), .B(
        Input[27]), .ZN(MCOutput_59_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_11_U1 ( .A(Input[11]), .B(Input[59]), .ZN(
        MCInst_XOR_r0_Inst_11_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_11_U1 ( .A(Input[43]), .B(Input[11]), .Z(
        MCOutput_43_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_12_U2 ( .A(MCInst_XOR_r0_Inst_12_n5), .B(
        Input[28]), .ZN(MCOutput_60_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_12_U1 ( .A(Input[12]), .B(Input[60]), .ZN(
        MCInst_XOR_r0_Inst_12_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_12_U1 ( .A(Input[44]), .B(Input[12]), .Z(
        MCOutput_44_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_13_U2 ( .A(MCInst_XOR_r0_Inst_13_n5), .B(
        Input[29]), .ZN(MCOutput_61_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_13_U1 ( .A(Input[13]), .B(Input[61]), .ZN(
        MCInst_XOR_r0_Inst_13_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_13_U1 ( .A(Input[45]), .B(Input[13]), .Z(
        MCOutput_45_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_14_U2 ( .A(MCInst_XOR_r0_Inst_14_n5), .B(
        Input[30]), .ZN(MCOutput_62_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_14_U1 ( .A(Input[14]), .B(Input[62]), .ZN(
        MCInst_XOR_r0_Inst_14_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_14_U1 ( .A(Input[46]), .B(Input[14]), .Z(
        MCOutput_46_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_15_U2 ( .A(MCInst_XOR_r0_Inst_15_n5), .B(
        Input[31]), .ZN(MCOutput_63_) );
  XNOR2_X1 MCInst_XOR_r0_Inst_15_U1 ( .A(Input[15]), .B(Input[63]), .ZN(
        MCInst_XOR_r0_Inst_15_n5) );
  XOR2_X1 MCInst_XOR_r1_Inst_15_U1 ( .A(Input[47]), .B(Input[15]), .Z(
        MCOutput_47_) );
  XOR2_X1 AddKeyXOR1_XORInst_0_0_U1 ( .A(MCOutput_48_), .B(Key[112]), .Z(
        AddRoundKeyOutput[48]) );
  XOR2_X1 AddKeyXOR1_XORInst_0_1_U1 ( .A(MCOutput_49_), .B(Key[113]), .Z(
        AddRoundKeyOutput[49]) );
  XOR2_X1 AddKeyXOR1_XORInst_0_2_U1 ( .A(MCOutput_50_), .B(Key[114]), .Z(
        AddRoundKeyOutput[50]) );
  XOR2_X1 AddKeyXOR1_XORInst_0_3_U1 ( .A(MCOutput_51_), .B(Key[115]), .Z(
        AddRoundKeyOutput[51]) );
  XOR2_X1 AddKeyXOR1_XORInst_1_0_U1 ( .A(MCOutput_52_), .B(Key[116]), .Z(
        AddRoundKeyOutput[52]) );
  XOR2_X1 AddKeyXOR1_XORInst_1_1_U1 ( .A(MCOutput_53_), .B(Key[117]), .Z(
        AddRoundKeyOutput[53]) );
  XOR2_X1 AddKeyXOR1_XORInst_1_2_U1 ( .A(MCOutput_54_), .B(Key[118]), .Z(
        AddRoundKeyOutput[54]) );
  XOR2_X1 AddKeyXOR1_XORInst_1_3_U1 ( .A(MCOutput_55_), .B(Key[119]), .Z(
        AddRoundKeyOutput[55]) );
  XOR2_X1 AddKeyXOR1_XORInst_2_0_U1 ( .A(MCOutput_56_), .B(Key[120]), .Z(
        AddRoundKeyOutput[56]) );
  XOR2_X1 AddKeyXOR1_XORInst_2_1_U1 ( .A(MCOutput_57_), .B(Key[121]), .Z(
        AddRoundKeyOutput[57]) );
  XOR2_X1 AddKeyXOR1_XORInst_2_2_U1 ( .A(MCOutput_58_), .B(Key[122]), .Z(
        AddRoundKeyOutput[58]) );
  XOR2_X1 AddKeyXOR1_XORInst_2_3_U1 ( .A(MCOutput_59_), .B(Key[123]), .Z(
        AddRoundKeyOutput[59]) );
  XOR2_X1 AddKeyXOR1_XORInst_3_0_U1 ( .A(MCOutput_60_), .B(Key[124]), .Z(
        AddRoundKeyOutput[60]) );
  XOR2_X1 AddKeyXOR1_XORInst_3_1_U1 ( .A(MCOutput_61_), .B(Key[125]), .Z(
        AddRoundKeyOutput[61]) );
  XOR2_X1 AddKeyXOR1_XORInst_3_2_U1 ( .A(MCOutput_62_), .B(Key[126]), .Z(
        AddRoundKeyOutput[62]) );
  XOR2_X1 AddKeyXOR1_XORInst_3_3_U1 ( .A(MCOutput_63_), .B(Key[127]), .Z(
        AddRoundKeyOutput[63]) );
  XOR2_X1 AddKeyConstXOR_XORInst_0_0_U1 ( .A(MCOutput_40_), .B(Key[104]), .Z(
        AddRoundKeyOutput[40]) );
  XOR2_X1 AddKeyConstXOR_XORInst_0_1_U1 ( .A(MCOutput_41_), .B(Key[105]), .Z(
        AddRoundKeyOutput[41]) );
  XOR2_X1 AddKeyConstXOR_XORInst_0_2_U1 ( .A(MCOutput_42_), .B(Key[106]), .Z(
        AddRoundKeyOutput[42]) );
  XOR2_X1 AddKeyConstXOR_XORInst_0_3_U1 ( .A(MCOutput_43_), .B(Key[107]), .Z(
        AddRoundKeyOutput[43]) );
  XOR2_X1 AddKeyConstXOR_XORInst_1_0_U1 ( .A(MCOutput_44_), .B(Key[108]), .Z(
        AddRoundKeyOutput[44]) );
  XOR2_X1 AddKeyConstXOR_XORInst_1_1_U1 ( .A(MCOutput_45_), .B(Key[109]), .Z(
        AddRoundKeyOutput[45]) );
  XOR2_X1 AddKeyConstXOR_XORInst_1_2_U1 ( .A(MCOutput_46_), .B(Key[110]), .Z(
        AddRoundKeyOutput[46]) );
  XOR2_X1 AddKeyConstXOR_XORInst_1_3_U1 ( .A(MCOutput_47_), .B(Key[111]), .Z(
        AddRoundKeyOutput[47]) );
  XOR2_X1 AddKeyXOR2_XORInst_0_0_U1 ( .A(Input[0]), .B(Key[64]), .Z(
        AddRoundKeyOutput[0]) );
  XOR2_X1 AddKeyXOR2_XORInst_0_1_U1 ( .A(Input[1]), .B(Key[65]), .Z(
        AddRoundKeyOutput[1]) );
  XOR2_X1 AddKeyXOR2_XORInst_0_2_U1 ( .A(Input[2]), .B(Key[66]), .Z(
        AddRoundKeyOutput[2]) );
  XOR2_X1 AddKeyXOR2_XORInst_0_3_U1 ( .A(Input[3]), .B(Key[67]), .Z(
        AddRoundKeyOutput[3]) );
  XOR2_X1 AddKeyXOR2_XORInst_1_0_U1 ( .A(Input[4]), .B(Key[68]), .Z(
        AddRoundKeyOutput[4]) );
  XOR2_X1 AddKeyXOR2_XORInst_1_1_U1 ( .A(Input[5]), .B(Key[69]), .Z(
        AddRoundKeyOutput[5]) );
  XOR2_X1 AddKeyXOR2_XORInst_1_2_U1 ( .A(Input[6]), .B(Key[70]), .Z(
        AddRoundKeyOutput[6]) );
  XOR2_X1 AddKeyXOR2_XORInst_1_3_U1 ( .A(Input[7]), .B(Key[71]), .Z(
        AddRoundKeyOutput[7]) );
  XOR2_X1 AddKeyXOR2_XORInst_2_0_U1 ( .A(Input[8]), .B(Key[72]), .Z(
        AddRoundKeyOutput[8]) );
  XOR2_X1 AddKeyXOR2_XORInst_2_1_U1 ( .A(Input[9]), .B(Key[73]), .Z(
        AddRoundKeyOutput[9]) );
  XOR2_X1 AddKeyXOR2_XORInst_2_2_U1 ( .A(Input[10]), .B(Key[74]), .Z(
        AddRoundKeyOutput[10]) );
  XOR2_X1 AddKeyXOR2_XORInst_2_3_U1 ( .A(Input[11]), .B(Key[75]), .Z(
        AddRoundKeyOutput[11]) );
  XOR2_X1 AddKeyXOR2_XORInst_3_0_U1 ( .A(Input[12]), .B(Key[76]), .Z(
        AddRoundKeyOutput[12]) );
  XOR2_X1 AddKeyXOR2_XORInst_3_1_U1 ( .A(Input[13]), .B(Key[77]), .Z(
        AddRoundKeyOutput[13]) );
  XOR2_X1 AddKeyXOR2_XORInst_3_2_U1 ( .A(Input[14]), .B(Key[78]), .Z(
        AddRoundKeyOutput[14]) );
  XOR2_X1 AddKeyXOR2_XORInst_3_3_U1 ( .A(Input[15]), .B(Key[79]), .Z(
        AddRoundKeyOutput[15]) );
  XOR2_X1 AddKeyXOR2_XORInst_4_0_U1 ( .A(Input[16]), .B(Key[80]), .Z(
        AddRoundKeyOutput[16]) );
  XOR2_X1 AddKeyXOR2_XORInst_4_1_U1 ( .A(Input[17]), .B(Key[81]), .Z(
        AddRoundKeyOutput[17]) );
  XOR2_X1 AddKeyXOR2_XORInst_4_2_U1 ( .A(Input[18]), .B(Key[82]), .Z(
        AddRoundKeyOutput[18]) );
  XOR2_X1 AddKeyXOR2_XORInst_4_3_U1 ( .A(Input[19]), .B(Key[83]), .Z(
        AddRoundKeyOutput[19]) );
  XOR2_X1 AddKeyXOR2_XORInst_5_0_U1 ( .A(Input[20]), .B(Key[84]), .Z(
        AddRoundKeyOutput[20]) );
  XOR2_X1 AddKeyXOR2_XORInst_5_1_U1 ( .A(Input[21]), .B(Key[85]), .Z(
        AddRoundKeyOutput[21]) );
  XOR2_X1 AddKeyXOR2_XORInst_5_2_U1 ( .A(Input[22]), .B(Key[86]), .Z(
        AddRoundKeyOutput[22]) );
  XOR2_X1 AddKeyXOR2_XORInst_5_3_U1 ( .A(Input[23]), .B(Key[87]), .Z(
        AddRoundKeyOutput[23]) );
  XOR2_X1 AddKeyXOR2_XORInst_6_0_U1 ( .A(Input[24]), .B(Key[88]), .Z(
        AddRoundKeyOutput[24]) );
  XOR2_X1 AddKeyXOR2_XORInst_6_1_U1 ( .A(Input[25]), .B(Key[89]), .Z(
        AddRoundKeyOutput[25]) );
  XOR2_X1 AddKeyXOR2_XORInst_6_2_U1 ( .A(Input[26]), .B(Key[90]), .Z(
        AddRoundKeyOutput[26]) );
  XOR2_X1 AddKeyXOR2_XORInst_6_3_U1 ( .A(Input[27]), .B(Key[91]), .Z(
        AddRoundKeyOutput[27]) );
  XOR2_X1 AddKeyXOR2_XORInst_7_0_U1 ( .A(Input[28]), .B(Key[92]), .Z(
        AddRoundKeyOutput[28]) );
  XOR2_X1 AddKeyXOR2_XORInst_7_1_U1 ( .A(Input[29]), .B(Key[93]), .Z(
        AddRoundKeyOutput[29]) );
  XOR2_X1 AddKeyXOR2_XORInst_7_2_U1 ( .A(Input[30]), .B(Key[94]), .Z(
        AddRoundKeyOutput[30]) );
  XOR2_X1 AddKeyXOR2_XORInst_7_3_U1 ( .A(Input[31]), .B(Key[95]), .Z(
        AddRoundKeyOutput[31]) );
  XOR2_X1 AddKeyXOR2_XORInst_8_0_U1 ( .A(MCOutput_32_), .B(Key[96]), .Z(
        AddRoundKeyOutput[32]) );
  XOR2_X1 AddKeyXOR2_XORInst_8_1_U1 ( .A(MCOutput_33_), .B(Key[97]), .Z(
        AddRoundKeyOutput[33]) );
  XOR2_X1 AddKeyXOR2_XORInst_8_2_U1 ( .A(MCOutput_34_), .B(Key[98]), .Z(
        AddRoundKeyOutput[34]) );
  XOR2_X1 AddKeyXOR2_XORInst_8_3_U1 ( .A(MCOutput_35_), .B(Key[99]), .Z(
        AddRoundKeyOutput[35]) );
  XOR2_X1 AddKeyXOR2_XORInst_9_0_U1 ( .A(MCOutput_36_), .B(Key[100]), .Z(
        AddRoundKeyOutput[36]) );
  XOR2_X1 AddKeyXOR2_XORInst_9_1_U1 ( .A(MCOutput_37_), .B(Key[101]), .Z(
        AddRoundKeyOutput[37]) );
  XOR2_X1 AddKeyXOR2_XORInst_9_2_U1 ( .A(MCOutput_38_), .B(Key[102]), .Z(
        AddRoundKeyOutput[38]) );
  XOR2_X1 AddKeyXOR2_XORInst_9_3_U1 ( .A(MCOutput_39_), .B(Key[103]), .Z(
        AddRoundKeyOutput[39]) );
  DFF_X1 StateReg_s_current_state_reg_0_ ( .D(AddRoundKeyOutput[0]), .CK(clk), 
        .Q(PermutationOutput[60]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_1_ ( .D(AddRoundKeyOutput[1]), .CK(clk), 
        .Q(PermutationOutput[61]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_2_ ( .D(AddRoundKeyOutput[2]), .CK(clk), 
        .Q(PermutationOutput[62]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_3_ ( .D(AddRoundKeyOutput[3]), .CK(clk), 
        .Q(PermutationOutput[63]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_4_ ( .D(AddRoundKeyOutput[4]), .CK(clk), 
        .Q(PermutationOutput[48]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_5_ ( .D(AddRoundKeyOutput[5]), .CK(clk), 
        .Q(PermutationOutput[49]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_6_ ( .D(AddRoundKeyOutput[6]), .CK(clk), 
        .Q(PermutationOutput[50]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_7_ ( .D(AddRoundKeyOutput[7]), .CK(clk), 
        .Q(PermutationOutput[51]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_8_ ( .D(AddRoundKeyOutput[8]), .CK(clk), 
        .Q(PermutationOutput[52]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_9_ ( .D(AddRoundKeyOutput[9]), .CK(clk), 
        .Q(PermutationOutput[53]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_10_ ( .D(AddRoundKeyOutput[10]), .CK(clk), .Q(PermutationOutput[54]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_11_ ( .D(AddRoundKeyOutput[11]), .CK(clk), .Q(PermutationOutput[55]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_12_ ( .D(AddRoundKeyOutput[12]), .CK(clk), .Q(PermutationOutput[56]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_13_ ( .D(AddRoundKeyOutput[13]), .CK(clk), .Q(PermutationOutput[57]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_14_ ( .D(AddRoundKeyOutput[14]), .CK(clk), .Q(PermutationOutput[58]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_15_ ( .D(AddRoundKeyOutput[15]), .CK(clk), .Q(PermutationOutput[59]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_16_ ( .D(AddRoundKeyOutput[16]), .CK(clk), .Q(PermutationOutput[32]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_17_ ( .D(AddRoundKeyOutput[17]), .CK(clk), .Q(PermutationOutput[33]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_18_ ( .D(AddRoundKeyOutput[18]), .CK(clk), .Q(PermutationOutput[34]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_19_ ( .D(AddRoundKeyOutput[19]), .CK(clk), .Q(PermutationOutput[35]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_20_ ( .D(AddRoundKeyOutput[20]), .CK(clk), .Q(PermutationOutput[44]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_21_ ( .D(AddRoundKeyOutput[21]), .CK(clk), .Q(PermutationOutput[45]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_22_ ( .D(AddRoundKeyOutput[22]), .CK(clk), .Q(PermutationOutput[46]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_23_ ( .D(AddRoundKeyOutput[23]), .CK(clk), .Q(PermutationOutput[47]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_24_ ( .D(AddRoundKeyOutput[24]), .CK(clk), .Q(PermutationOutput[40]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_25_ ( .D(AddRoundKeyOutput[25]), .CK(clk), .Q(PermutationOutput[41]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_26_ ( .D(AddRoundKeyOutput[26]), .CK(clk), .Q(PermutationOutput[42]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_27_ ( .D(AddRoundKeyOutput[27]), .CK(clk), .Q(PermutationOutput[43]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_28_ ( .D(AddRoundKeyOutput[28]), .CK(clk), .Q(PermutationOutput[36]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_29_ ( .D(AddRoundKeyOutput[29]), .CK(clk), .Q(PermutationOutput[37]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_30_ ( .D(AddRoundKeyOutput[30]), .CK(clk), .Q(PermutationOutput[38]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_31_ ( .D(AddRoundKeyOutput[31]), .CK(clk), .Q(PermutationOutput[39]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_32_ ( .D(AddRoundKeyOutput[32]), .CK(clk), .Q(PermutationOutput[16]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_33_ ( .D(AddRoundKeyOutput[33]), .CK(clk), .Q(PermutationOutput[17]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_34_ ( .D(AddRoundKeyOutput[34]), .CK(clk), .Q(PermutationOutput[18]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_35_ ( .D(AddRoundKeyOutput[35]), .CK(clk), .Q(PermutationOutput[19]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_36_ ( .D(AddRoundKeyOutput[36]), .CK(clk), .Q(PermutationOutput[28]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_37_ ( .D(AddRoundKeyOutput[37]), .CK(clk), .Q(PermutationOutput[29]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_38_ ( .D(AddRoundKeyOutput[38]), .CK(clk), .Q(PermutationOutput[30]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_39_ ( .D(AddRoundKeyOutput[39]), .CK(clk), .Q(PermutationOutput[31]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_40_ ( .D(AddRoundKeyOutput[40]), .CK(clk), .Q(PermutationOutput[24]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_41_ ( .D(AddRoundKeyOutput[41]), .CK(clk), .Q(PermutationOutput[25]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_42_ ( .D(AddRoundKeyOutput[42]), .CK(clk), .Q(PermutationOutput[26]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_43_ ( .D(AddRoundKeyOutput[43]), .CK(clk), .Q(PermutationOutput[27]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_44_ ( .D(AddRoundKeyOutput[44]), .CK(clk), .Q(PermutationOutput[20]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_45_ ( .D(AddRoundKeyOutput[45]), .CK(clk), .Q(PermutationOutput[21]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_46_ ( .D(AddRoundKeyOutput[46]), .CK(clk), .Q(PermutationOutput[22]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_47_ ( .D(AddRoundKeyOutput[47]), .CK(clk), .Q(PermutationOutput[23]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_48_ ( .D(AddRoundKeyOutput[48]), .CK(clk), .Q(PermutationOutput[4]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_49_ ( .D(AddRoundKeyOutput[49]), .CK(clk), .Q(PermutationOutput[5]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_50_ ( .D(AddRoundKeyOutput[50]), .CK(clk), .Q(PermutationOutput[6]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_51_ ( .D(AddRoundKeyOutput[51]), .CK(clk), .Q(PermutationOutput[7]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_52_ ( .D(AddRoundKeyOutput[52]), .CK(clk), .Q(PermutationOutput[8]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_53_ ( .D(AddRoundKeyOutput[53]), .CK(clk), .Q(PermutationOutput[9]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_54_ ( .D(AddRoundKeyOutput[54]), .CK(clk), .Q(PermutationOutput[10]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_55_ ( .D(AddRoundKeyOutput[55]), .CK(clk), .Q(PermutationOutput[11]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_56_ ( .D(AddRoundKeyOutput[56]), .CK(clk), .Q(PermutationOutput[12]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_57_ ( .D(AddRoundKeyOutput[57]), .CK(clk), .Q(PermutationOutput[13]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_58_ ( .D(AddRoundKeyOutput[58]), .CK(clk), .Q(PermutationOutput[14]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_59_ ( .D(AddRoundKeyOutput[59]), .CK(clk), .Q(PermutationOutput[15]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_60_ ( .D(AddRoundKeyOutput[60]), .CK(clk), .Q(PermutationOutput[0]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_61_ ( .D(AddRoundKeyOutput[61]), .CK(clk), .Q(PermutationOutput[1]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_62_ ( .D(AddRoundKeyOutput[62]), .CK(clk), .Q(PermutationOutput[2]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_63_ ( .D(AddRoundKeyOutput[63]), .CK(clk), .Q(PermutationOutput[3]), .QN() );
  NOR2_X1 SubCellInst_LFInst_0_LFInst_0_U6 ( .A1(
        SubCellInst_LFInst_0_LFInst_0_n15), .A2(
        SubCellInst_LFInst_0_LFInst_0_n14), .ZN(MCOutput2[0]) );
  AND2_X1 SubCellInst_LFInst_0_LFInst_0_U5 ( .A1(PermutationOutput[3]), .A2(
        PermutationOutput[2]), .ZN(SubCellInst_LFInst_0_LFInst_0_n14) );
  NOR2_X1 SubCellInst_LFInst_0_LFInst_0_U4 ( .A1(PermutationOutput[1]), .A2(
        SubCellInst_LFInst_0_LFInst_0_n13), .ZN(
        SubCellInst_LFInst_0_LFInst_0_n15) );
  NOR2_X1 SubCellInst_LFInst_0_LFInst_0_U3 ( .A1(
        SubCellInst_LFInst_0_LFInst_0_n12), .A2(
        SubCellInst_LFInst_0_LFInst_0_n11), .ZN(
        SubCellInst_LFInst_0_LFInst_0_n13) );
  NOR2_X1 SubCellInst_LFInst_0_LFInst_0_U2 ( .A1(PermutationOutput[3]), .A2(
        PermutationOutput[2]), .ZN(SubCellInst_LFInst_0_LFInst_0_n11) );
  INV_X1 SubCellInst_LFInst_0_LFInst_0_U1 ( .A(PermutationOutput[0]), .ZN(
        SubCellInst_LFInst_0_LFInst_0_n12) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_1_U4 ( .A1(
        SubCellInst_LFInst_0_LFInst_1_n9), .A2(
        SubCellInst_LFInst_0_LFInst_1_n8), .ZN(MCOutput2[1]) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_1_U3 ( .A1(PermutationOutput[0]), .A2(
        PermutationOutput[2]), .ZN(SubCellInst_LFInst_0_LFInst_1_n8) );
  OR2_X1 SubCellInst_LFInst_0_LFInst_1_U2 ( .A1(PermutationOutput[3]), .A2(
        SubCellInst_LFInst_0_LFInst_1_n7), .ZN(
        SubCellInst_LFInst_0_LFInst_1_n9) );
  NOR2_X1 SubCellInst_LFInst_0_LFInst_1_U1 ( .A1(PermutationOutput[0]), .A2(
        PermutationOutput[2]), .ZN(SubCellInst_LFInst_0_LFInst_1_n7) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_2_U6 ( .A1(
        SubCellInst_LFInst_0_LFInst_2_n18), .A2(
        SubCellInst_LFInst_0_LFInst_2_n17), .ZN(MCOutput2[2]) );
  OR2_X1 SubCellInst_LFInst_0_LFInst_2_U5 ( .A1(PermutationOutput[0]), .A2(
        PermutationOutput[3]), .ZN(SubCellInst_LFInst_0_LFInst_2_n17) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_2_U4 ( .A1(PermutationOutput[1]), .A2(
        SubCellInst_LFInst_0_LFInst_2_n16), .ZN(
        SubCellInst_LFInst_0_LFInst_2_n18) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_2_U3 ( .A1(
        SubCellInst_LFInst_0_LFInst_2_n15), .A2(
        SubCellInst_LFInst_0_LFInst_2_n14), .ZN(
        SubCellInst_LFInst_0_LFInst_2_n16) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_2_U2 ( .A1(PermutationOutput[0]), .A2(
        PermutationOutput[3]), .ZN(SubCellInst_LFInst_0_LFInst_2_n14) );
  INV_X1 SubCellInst_LFInst_0_LFInst_2_U1 ( .A(PermutationOutput[2]), .ZN(
        SubCellInst_LFInst_0_LFInst_2_n15) );
  NOR2_X1 SubCellInst_LFInst_0_LFInst_3_U4 ( .A1(PermutationOutput[1]), .A2(
        PermutationOutput[2]), .ZN(SubCellInst_LFInst_0_LFInst_3_n8) );
  NOR2_X1 SubCellInst_LFInst_0_LFInst_3_U3 ( .A1(PermutationOutput[3]), .A2(
        SubCellInst_LFInst_0_LFInst_3_n7), .ZN(
        SubCellInst_LFInst_0_LFInst_3_n9) );
  AND2_X1 SubCellInst_LFInst_0_LFInst_3_U2 ( .A1(PermutationOutput[1]), .A2(
        PermutationOutput[0]), .ZN(SubCellInst_LFInst_0_LFInst_3_n7) );
  OR2_X1 SubCellInst_LFInst_0_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_0_LFInst_3_n9), .A2(
        SubCellInst_LFInst_0_LFInst_3_n8), .ZN(MCOutput2[3]) );
  NOR2_X1 SubCellInst_LFInst_1_LFInst_0_U6 ( .A1(
        SubCellInst_LFInst_1_LFInst_0_n15), .A2(
        SubCellInst_LFInst_1_LFInst_0_n14), .ZN(MCOutput2[4]) );
  AND2_X1 SubCellInst_LFInst_1_LFInst_0_U5 ( .A1(PermutationOutput[7]), .A2(
        PermutationOutput[6]), .ZN(SubCellInst_LFInst_1_LFInst_0_n14) );
  NOR2_X1 SubCellInst_LFInst_1_LFInst_0_U4 ( .A1(PermutationOutput[5]), .A2(
        SubCellInst_LFInst_1_LFInst_0_n13), .ZN(
        SubCellInst_LFInst_1_LFInst_0_n15) );
  NOR2_X1 SubCellInst_LFInst_1_LFInst_0_U3 ( .A1(
        SubCellInst_LFInst_1_LFInst_0_n12), .A2(
        SubCellInst_LFInst_1_LFInst_0_n11), .ZN(
        SubCellInst_LFInst_1_LFInst_0_n13) );
  NOR2_X1 SubCellInst_LFInst_1_LFInst_0_U2 ( .A1(PermutationOutput[7]), .A2(
        PermutationOutput[6]), .ZN(SubCellInst_LFInst_1_LFInst_0_n11) );
  INV_X1 SubCellInst_LFInst_1_LFInst_0_U1 ( .A(PermutationOutput[4]), .ZN(
        SubCellInst_LFInst_1_LFInst_0_n12) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_1_U4 ( .A1(
        SubCellInst_LFInst_1_LFInst_1_n9), .A2(
        SubCellInst_LFInst_1_LFInst_1_n8), .ZN(MCOutput2[5]) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_1_U3 ( .A1(PermutationOutput[4]), .A2(
        PermutationOutput[6]), .ZN(SubCellInst_LFInst_1_LFInst_1_n8) );
  OR2_X1 SubCellInst_LFInst_1_LFInst_1_U2 ( .A1(PermutationOutput[7]), .A2(
        SubCellInst_LFInst_1_LFInst_1_n7), .ZN(
        SubCellInst_LFInst_1_LFInst_1_n9) );
  NOR2_X1 SubCellInst_LFInst_1_LFInst_1_U1 ( .A1(PermutationOutput[4]), .A2(
        PermutationOutput[6]), .ZN(SubCellInst_LFInst_1_LFInst_1_n7) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_2_U6 ( .A1(
        SubCellInst_LFInst_1_LFInst_2_n18), .A2(
        SubCellInst_LFInst_1_LFInst_2_n17), .ZN(MCOutput2[6]) );
  OR2_X1 SubCellInst_LFInst_1_LFInst_2_U5 ( .A1(PermutationOutput[4]), .A2(
        PermutationOutput[7]), .ZN(SubCellInst_LFInst_1_LFInst_2_n17) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_2_U4 ( .A1(PermutationOutput[5]), .A2(
        SubCellInst_LFInst_1_LFInst_2_n16), .ZN(
        SubCellInst_LFInst_1_LFInst_2_n18) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_2_U3 ( .A1(
        SubCellInst_LFInst_1_LFInst_2_n15), .A2(
        SubCellInst_LFInst_1_LFInst_2_n14), .ZN(
        SubCellInst_LFInst_1_LFInst_2_n16) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_2_U2 ( .A1(PermutationOutput[4]), .A2(
        PermutationOutput[7]), .ZN(SubCellInst_LFInst_1_LFInst_2_n14) );
  INV_X1 SubCellInst_LFInst_1_LFInst_2_U1 ( .A(PermutationOutput[6]), .ZN(
        SubCellInst_LFInst_1_LFInst_2_n15) );
  NOR2_X1 SubCellInst_LFInst_1_LFInst_3_U4 ( .A1(PermutationOutput[5]), .A2(
        PermutationOutput[6]), .ZN(SubCellInst_LFInst_1_LFInst_3_n8) );
  NOR2_X1 SubCellInst_LFInst_1_LFInst_3_U3 ( .A1(PermutationOutput[7]), .A2(
        SubCellInst_LFInst_1_LFInst_3_n7), .ZN(
        SubCellInst_LFInst_1_LFInst_3_n9) );
  AND2_X1 SubCellInst_LFInst_1_LFInst_3_U2 ( .A1(PermutationOutput[5]), .A2(
        PermutationOutput[4]), .ZN(SubCellInst_LFInst_1_LFInst_3_n7) );
  OR2_X1 SubCellInst_LFInst_1_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_1_LFInst_3_n9), .A2(
        SubCellInst_LFInst_1_LFInst_3_n8), .ZN(MCOutput2[7]) );
  NOR2_X1 SubCellInst_LFInst_2_LFInst_0_U6 ( .A1(
        SubCellInst_LFInst_2_LFInst_0_n15), .A2(
        SubCellInst_LFInst_2_LFInst_0_n14), .ZN(MCOutput2[8]) );
  AND2_X1 SubCellInst_LFInst_2_LFInst_0_U5 ( .A1(PermutationOutput[11]), .A2(
        PermutationOutput[10]), .ZN(SubCellInst_LFInst_2_LFInst_0_n14) );
  NOR2_X1 SubCellInst_LFInst_2_LFInst_0_U4 ( .A1(PermutationOutput[9]), .A2(
        SubCellInst_LFInst_2_LFInst_0_n13), .ZN(
        SubCellInst_LFInst_2_LFInst_0_n15) );
  NOR2_X1 SubCellInst_LFInst_2_LFInst_0_U3 ( .A1(
        SubCellInst_LFInst_2_LFInst_0_n12), .A2(
        SubCellInst_LFInst_2_LFInst_0_n11), .ZN(
        SubCellInst_LFInst_2_LFInst_0_n13) );
  NOR2_X1 SubCellInst_LFInst_2_LFInst_0_U2 ( .A1(PermutationOutput[11]), .A2(
        PermutationOutput[10]), .ZN(SubCellInst_LFInst_2_LFInst_0_n11) );
  INV_X1 SubCellInst_LFInst_2_LFInst_0_U1 ( .A(PermutationOutput[8]), .ZN(
        SubCellInst_LFInst_2_LFInst_0_n12) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_1_U4 ( .A1(
        SubCellInst_LFInst_2_LFInst_1_n9), .A2(
        SubCellInst_LFInst_2_LFInst_1_n8), .ZN(MCOutput2[9]) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_1_U3 ( .A1(PermutationOutput[8]), .A2(
        PermutationOutput[10]), .ZN(SubCellInst_LFInst_2_LFInst_1_n8) );
  OR2_X1 SubCellInst_LFInst_2_LFInst_1_U2 ( .A1(PermutationOutput[11]), .A2(
        SubCellInst_LFInst_2_LFInst_1_n7), .ZN(
        SubCellInst_LFInst_2_LFInst_1_n9) );
  NOR2_X1 SubCellInst_LFInst_2_LFInst_1_U1 ( .A1(PermutationOutput[8]), .A2(
        PermutationOutput[10]), .ZN(SubCellInst_LFInst_2_LFInst_1_n7) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_2_U6 ( .A1(
        SubCellInst_LFInst_2_LFInst_2_n18), .A2(
        SubCellInst_LFInst_2_LFInst_2_n17), .ZN(MCOutput2[10]) );
  OR2_X1 SubCellInst_LFInst_2_LFInst_2_U5 ( .A1(PermutationOutput[8]), .A2(
        PermutationOutput[11]), .ZN(SubCellInst_LFInst_2_LFInst_2_n17) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_2_U4 ( .A1(PermutationOutput[9]), .A2(
        SubCellInst_LFInst_2_LFInst_2_n16), .ZN(
        SubCellInst_LFInst_2_LFInst_2_n18) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_2_U3 ( .A1(
        SubCellInst_LFInst_2_LFInst_2_n15), .A2(
        SubCellInst_LFInst_2_LFInst_2_n14), .ZN(
        SubCellInst_LFInst_2_LFInst_2_n16) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_2_U2 ( .A1(PermutationOutput[8]), .A2(
        PermutationOutput[11]), .ZN(SubCellInst_LFInst_2_LFInst_2_n14) );
  INV_X1 SubCellInst_LFInst_2_LFInst_2_U1 ( .A(PermutationOutput[10]), .ZN(
        SubCellInst_LFInst_2_LFInst_2_n15) );
  NOR2_X1 SubCellInst_LFInst_2_LFInst_3_U4 ( .A1(PermutationOutput[9]), .A2(
        PermutationOutput[10]), .ZN(SubCellInst_LFInst_2_LFInst_3_n8) );
  NOR2_X1 SubCellInst_LFInst_2_LFInst_3_U3 ( .A1(PermutationOutput[11]), .A2(
        SubCellInst_LFInst_2_LFInst_3_n7), .ZN(
        SubCellInst_LFInst_2_LFInst_3_n9) );
  AND2_X1 SubCellInst_LFInst_2_LFInst_3_U2 ( .A1(PermutationOutput[9]), .A2(
        PermutationOutput[8]), .ZN(SubCellInst_LFInst_2_LFInst_3_n7) );
  OR2_X1 SubCellInst_LFInst_2_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_2_LFInst_3_n9), .A2(
        SubCellInst_LFInst_2_LFInst_3_n8), .ZN(MCOutput2[11]) );
  NOR2_X1 SubCellInst_LFInst_3_LFInst_0_U6 ( .A1(
        SubCellInst_LFInst_3_LFInst_0_n15), .A2(
        SubCellInst_LFInst_3_LFInst_0_n14), .ZN(MCOutput2[12]) );
  AND2_X1 SubCellInst_LFInst_3_LFInst_0_U5 ( .A1(PermutationOutput[15]), .A2(
        PermutationOutput[14]), .ZN(SubCellInst_LFInst_3_LFInst_0_n14) );
  NOR2_X1 SubCellInst_LFInst_3_LFInst_0_U4 ( .A1(PermutationOutput[13]), .A2(
        SubCellInst_LFInst_3_LFInst_0_n13), .ZN(
        SubCellInst_LFInst_3_LFInst_0_n15) );
  NOR2_X1 SubCellInst_LFInst_3_LFInst_0_U3 ( .A1(
        SubCellInst_LFInst_3_LFInst_0_n12), .A2(
        SubCellInst_LFInst_3_LFInst_0_n11), .ZN(
        SubCellInst_LFInst_3_LFInst_0_n13) );
  NOR2_X1 SubCellInst_LFInst_3_LFInst_0_U2 ( .A1(PermutationOutput[15]), .A2(
        PermutationOutput[14]), .ZN(SubCellInst_LFInst_3_LFInst_0_n11) );
  INV_X1 SubCellInst_LFInst_3_LFInst_0_U1 ( .A(PermutationOutput[12]), .ZN(
        SubCellInst_LFInst_3_LFInst_0_n12) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_1_U4 ( .A1(
        SubCellInst_LFInst_3_LFInst_1_n9), .A2(
        SubCellInst_LFInst_3_LFInst_1_n8), .ZN(MCOutput2[13]) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_1_U3 ( .A1(PermutationOutput[12]), .A2(
        PermutationOutput[14]), .ZN(SubCellInst_LFInst_3_LFInst_1_n8) );
  OR2_X1 SubCellInst_LFInst_3_LFInst_1_U2 ( .A1(PermutationOutput[15]), .A2(
        SubCellInst_LFInst_3_LFInst_1_n7), .ZN(
        SubCellInst_LFInst_3_LFInst_1_n9) );
  NOR2_X1 SubCellInst_LFInst_3_LFInst_1_U1 ( .A1(PermutationOutput[12]), .A2(
        PermutationOutput[14]), .ZN(SubCellInst_LFInst_3_LFInst_1_n7) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_2_U6 ( .A1(
        SubCellInst_LFInst_3_LFInst_2_n18), .A2(
        SubCellInst_LFInst_3_LFInst_2_n17), .ZN(MCOutput2[14]) );
  OR2_X1 SubCellInst_LFInst_3_LFInst_2_U5 ( .A1(PermutationOutput[12]), .A2(
        PermutationOutput[15]), .ZN(SubCellInst_LFInst_3_LFInst_2_n17) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_2_U4 ( .A1(PermutationOutput[13]), .A2(
        SubCellInst_LFInst_3_LFInst_2_n16), .ZN(
        SubCellInst_LFInst_3_LFInst_2_n18) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_2_U3 ( .A1(
        SubCellInst_LFInst_3_LFInst_2_n15), .A2(
        SubCellInst_LFInst_3_LFInst_2_n14), .ZN(
        SubCellInst_LFInst_3_LFInst_2_n16) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_2_U2 ( .A1(PermutationOutput[12]), .A2(
        PermutationOutput[15]), .ZN(SubCellInst_LFInst_3_LFInst_2_n14) );
  INV_X1 SubCellInst_LFInst_3_LFInst_2_U1 ( .A(PermutationOutput[14]), .ZN(
        SubCellInst_LFInst_3_LFInst_2_n15) );
  NOR2_X1 SubCellInst_LFInst_3_LFInst_3_U4 ( .A1(PermutationOutput[13]), .A2(
        PermutationOutput[14]), .ZN(SubCellInst_LFInst_3_LFInst_3_n8) );
  NOR2_X1 SubCellInst_LFInst_3_LFInst_3_U3 ( .A1(PermutationOutput[15]), .A2(
        SubCellInst_LFInst_3_LFInst_3_n7), .ZN(
        SubCellInst_LFInst_3_LFInst_3_n9) );
  AND2_X1 SubCellInst_LFInst_3_LFInst_3_U2 ( .A1(PermutationOutput[13]), .A2(
        PermutationOutput[12]), .ZN(SubCellInst_LFInst_3_LFInst_3_n7) );
  OR2_X1 SubCellInst_LFInst_3_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_3_LFInst_3_n9), .A2(
        SubCellInst_LFInst_3_LFInst_3_n8), .ZN(MCOutput2[15]) );
  NOR2_X1 SubCellInst_LFInst_4_LFInst_0_U6 ( .A1(
        SubCellInst_LFInst_4_LFInst_0_n15), .A2(
        SubCellInst_LFInst_4_LFInst_0_n14), .ZN(MCOutput2[16]) );
  AND2_X1 SubCellInst_LFInst_4_LFInst_0_U5 ( .A1(PermutationOutput[19]), .A2(
        PermutationOutput[18]), .ZN(SubCellInst_LFInst_4_LFInst_0_n14) );
  NOR2_X1 SubCellInst_LFInst_4_LFInst_0_U4 ( .A1(PermutationOutput[17]), .A2(
        SubCellInst_LFInst_4_LFInst_0_n13), .ZN(
        SubCellInst_LFInst_4_LFInst_0_n15) );
  NOR2_X1 SubCellInst_LFInst_4_LFInst_0_U3 ( .A1(
        SubCellInst_LFInst_4_LFInst_0_n12), .A2(
        SubCellInst_LFInst_4_LFInst_0_n11), .ZN(
        SubCellInst_LFInst_4_LFInst_0_n13) );
  NOR2_X1 SubCellInst_LFInst_4_LFInst_0_U2 ( .A1(PermutationOutput[19]), .A2(
        PermutationOutput[18]), .ZN(SubCellInst_LFInst_4_LFInst_0_n11) );
  INV_X1 SubCellInst_LFInst_4_LFInst_0_U1 ( .A(PermutationOutput[16]), .ZN(
        SubCellInst_LFInst_4_LFInst_0_n12) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_1_U4 ( .A1(
        SubCellInst_LFInst_4_LFInst_1_n9), .A2(
        SubCellInst_LFInst_4_LFInst_1_n8), .ZN(MCOutput2[17]) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_1_U3 ( .A1(PermutationOutput[16]), .A2(
        PermutationOutput[18]), .ZN(SubCellInst_LFInst_4_LFInst_1_n8) );
  OR2_X1 SubCellInst_LFInst_4_LFInst_1_U2 ( .A1(PermutationOutput[19]), .A2(
        SubCellInst_LFInst_4_LFInst_1_n7), .ZN(
        SubCellInst_LFInst_4_LFInst_1_n9) );
  NOR2_X1 SubCellInst_LFInst_4_LFInst_1_U1 ( .A1(PermutationOutput[16]), .A2(
        PermutationOutput[18]), .ZN(SubCellInst_LFInst_4_LFInst_1_n7) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_2_U6 ( .A1(
        SubCellInst_LFInst_4_LFInst_2_n18), .A2(
        SubCellInst_LFInst_4_LFInst_2_n17), .ZN(MCOutput2[18]) );
  OR2_X1 SubCellInst_LFInst_4_LFInst_2_U5 ( .A1(PermutationOutput[16]), .A2(
        PermutationOutput[19]), .ZN(SubCellInst_LFInst_4_LFInst_2_n17) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_2_U4 ( .A1(PermutationOutput[17]), .A2(
        SubCellInst_LFInst_4_LFInst_2_n16), .ZN(
        SubCellInst_LFInst_4_LFInst_2_n18) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_2_U3 ( .A1(
        SubCellInst_LFInst_4_LFInst_2_n15), .A2(
        SubCellInst_LFInst_4_LFInst_2_n14), .ZN(
        SubCellInst_LFInst_4_LFInst_2_n16) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_2_U2 ( .A1(PermutationOutput[16]), .A2(
        PermutationOutput[19]), .ZN(SubCellInst_LFInst_4_LFInst_2_n14) );
  INV_X1 SubCellInst_LFInst_4_LFInst_2_U1 ( .A(PermutationOutput[18]), .ZN(
        SubCellInst_LFInst_4_LFInst_2_n15) );
  NOR2_X1 SubCellInst_LFInst_4_LFInst_3_U4 ( .A1(PermutationOutput[17]), .A2(
        PermutationOutput[18]), .ZN(SubCellInst_LFInst_4_LFInst_3_n8) );
  NOR2_X1 SubCellInst_LFInst_4_LFInst_3_U3 ( .A1(PermutationOutput[19]), .A2(
        SubCellInst_LFInst_4_LFInst_3_n7), .ZN(
        SubCellInst_LFInst_4_LFInst_3_n9) );
  AND2_X1 SubCellInst_LFInst_4_LFInst_3_U2 ( .A1(PermutationOutput[17]), .A2(
        PermutationOutput[16]), .ZN(SubCellInst_LFInst_4_LFInst_3_n7) );
  OR2_X1 SubCellInst_LFInst_4_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_4_LFInst_3_n9), .A2(
        SubCellInst_LFInst_4_LFInst_3_n8), .ZN(MCOutput2[19]) );
  NOR2_X1 SubCellInst_LFInst_5_LFInst_0_U6 ( .A1(
        SubCellInst_LFInst_5_LFInst_0_n15), .A2(
        SubCellInst_LFInst_5_LFInst_0_n14), .ZN(MCOutput2[20]) );
  AND2_X1 SubCellInst_LFInst_5_LFInst_0_U5 ( .A1(PermutationOutput[23]), .A2(
        PermutationOutput[22]), .ZN(SubCellInst_LFInst_5_LFInst_0_n14) );
  NOR2_X1 SubCellInst_LFInst_5_LFInst_0_U4 ( .A1(PermutationOutput[21]), .A2(
        SubCellInst_LFInst_5_LFInst_0_n13), .ZN(
        SubCellInst_LFInst_5_LFInst_0_n15) );
  NOR2_X1 SubCellInst_LFInst_5_LFInst_0_U3 ( .A1(
        SubCellInst_LFInst_5_LFInst_0_n12), .A2(
        SubCellInst_LFInst_5_LFInst_0_n11), .ZN(
        SubCellInst_LFInst_5_LFInst_0_n13) );
  NOR2_X1 SubCellInst_LFInst_5_LFInst_0_U2 ( .A1(PermutationOutput[23]), .A2(
        PermutationOutput[22]), .ZN(SubCellInst_LFInst_5_LFInst_0_n11) );
  INV_X1 SubCellInst_LFInst_5_LFInst_0_U1 ( .A(PermutationOutput[20]), .ZN(
        SubCellInst_LFInst_5_LFInst_0_n12) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_1_U4 ( .A1(
        SubCellInst_LFInst_5_LFInst_1_n9), .A2(
        SubCellInst_LFInst_5_LFInst_1_n8), .ZN(MCOutput2[21]) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_1_U3 ( .A1(PermutationOutput[20]), .A2(
        PermutationOutput[22]), .ZN(SubCellInst_LFInst_5_LFInst_1_n8) );
  OR2_X1 SubCellInst_LFInst_5_LFInst_1_U2 ( .A1(PermutationOutput[23]), .A2(
        SubCellInst_LFInst_5_LFInst_1_n7), .ZN(
        SubCellInst_LFInst_5_LFInst_1_n9) );
  NOR2_X1 SubCellInst_LFInst_5_LFInst_1_U1 ( .A1(PermutationOutput[20]), .A2(
        PermutationOutput[22]), .ZN(SubCellInst_LFInst_5_LFInst_1_n7) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_2_U6 ( .A1(
        SubCellInst_LFInst_5_LFInst_2_n18), .A2(
        SubCellInst_LFInst_5_LFInst_2_n17), .ZN(MCOutput2[22]) );
  OR2_X1 SubCellInst_LFInst_5_LFInst_2_U5 ( .A1(PermutationOutput[20]), .A2(
        PermutationOutput[23]), .ZN(SubCellInst_LFInst_5_LFInst_2_n17) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_2_U4 ( .A1(PermutationOutput[21]), .A2(
        SubCellInst_LFInst_5_LFInst_2_n16), .ZN(
        SubCellInst_LFInst_5_LFInst_2_n18) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_2_U3 ( .A1(
        SubCellInst_LFInst_5_LFInst_2_n15), .A2(
        SubCellInst_LFInst_5_LFInst_2_n14), .ZN(
        SubCellInst_LFInst_5_LFInst_2_n16) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_2_U2 ( .A1(PermutationOutput[20]), .A2(
        PermutationOutput[23]), .ZN(SubCellInst_LFInst_5_LFInst_2_n14) );
  INV_X1 SubCellInst_LFInst_5_LFInst_2_U1 ( .A(PermutationOutput[22]), .ZN(
        SubCellInst_LFInst_5_LFInst_2_n15) );
  NOR2_X1 SubCellInst_LFInst_5_LFInst_3_U4 ( .A1(PermutationOutput[21]), .A2(
        PermutationOutput[22]), .ZN(SubCellInst_LFInst_5_LFInst_3_n8) );
  NOR2_X1 SubCellInst_LFInst_5_LFInst_3_U3 ( .A1(PermutationOutput[23]), .A2(
        SubCellInst_LFInst_5_LFInst_3_n7), .ZN(
        SubCellInst_LFInst_5_LFInst_3_n9) );
  AND2_X1 SubCellInst_LFInst_5_LFInst_3_U2 ( .A1(PermutationOutput[21]), .A2(
        PermutationOutput[20]), .ZN(SubCellInst_LFInst_5_LFInst_3_n7) );
  OR2_X1 SubCellInst_LFInst_5_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_5_LFInst_3_n9), .A2(
        SubCellInst_LFInst_5_LFInst_3_n8), .ZN(MCOutput2[23]) );
  NOR2_X1 SubCellInst_LFInst_6_LFInst_0_U6 ( .A1(
        SubCellInst_LFInst_6_LFInst_0_n15), .A2(
        SubCellInst_LFInst_6_LFInst_0_n14), .ZN(MCOutput2[24]) );
  AND2_X1 SubCellInst_LFInst_6_LFInst_0_U5 ( .A1(PermutationOutput[27]), .A2(
        PermutationOutput[26]), .ZN(SubCellInst_LFInst_6_LFInst_0_n14) );
  NOR2_X1 SubCellInst_LFInst_6_LFInst_0_U4 ( .A1(PermutationOutput[25]), .A2(
        SubCellInst_LFInst_6_LFInst_0_n13), .ZN(
        SubCellInst_LFInst_6_LFInst_0_n15) );
  NOR2_X1 SubCellInst_LFInst_6_LFInst_0_U3 ( .A1(
        SubCellInst_LFInst_6_LFInst_0_n12), .A2(
        SubCellInst_LFInst_6_LFInst_0_n11), .ZN(
        SubCellInst_LFInst_6_LFInst_0_n13) );
  NOR2_X1 SubCellInst_LFInst_6_LFInst_0_U2 ( .A1(PermutationOutput[27]), .A2(
        PermutationOutput[26]), .ZN(SubCellInst_LFInst_6_LFInst_0_n11) );
  INV_X1 SubCellInst_LFInst_6_LFInst_0_U1 ( .A(PermutationOutput[24]), .ZN(
        SubCellInst_LFInst_6_LFInst_0_n12) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_1_U4 ( .A1(
        SubCellInst_LFInst_6_LFInst_1_n9), .A2(
        SubCellInst_LFInst_6_LFInst_1_n8), .ZN(MCOutput2[25]) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_1_U3 ( .A1(PermutationOutput[24]), .A2(
        PermutationOutput[26]), .ZN(SubCellInst_LFInst_6_LFInst_1_n8) );
  OR2_X1 SubCellInst_LFInst_6_LFInst_1_U2 ( .A1(PermutationOutput[27]), .A2(
        SubCellInst_LFInst_6_LFInst_1_n7), .ZN(
        SubCellInst_LFInst_6_LFInst_1_n9) );
  NOR2_X1 SubCellInst_LFInst_6_LFInst_1_U1 ( .A1(PermutationOutput[24]), .A2(
        PermutationOutput[26]), .ZN(SubCellInst_LFInst_6_LFInst_1_n7) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_2_U6 ( .A1(
        SubCellInst_LFInst_6_LFInst_2_n18), .A2(
        SubCellInst_LFInst_6_LFInst_2_n17), .ZN(MCOutput2[26]) );
  OR2_X1 SubCellInst_LFInst_6_LFInst_2_U5 ( .A1(PermutationOutput[24]), .A2(
        PermutationOutput[27]), .ZN(SubCellInst_LFInst_6_LFInst_2_n17) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_2_U4 ( .A1(PermutationOutput[25]), .A2(
        SubCellInst_LFInst_6_LFInst_2_n16), .ZN(
        SubCellInst_LFInst_6_LFInst_2_n18) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_2_U3 ( .A1(
        SubCellInst_LFInst_6_LFInst_2_n15), .A2(
        SubCellInst_LFInst_6_LFInst_2_n14), .ZN(
        SubCellInst_LFInst_6_LFInst_2_n16) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_2_U2 ( .A1(PermutationOutput[24]), .A2(
        PermutationOutput[27]), .ZN(SubCellInst_LFInst_6_LFInst_2_n14) );
  INV_X1 SubCellInst_LFInst_6_LFInst_2_U1 ( .A(PermutationOutput[26]), .ZN(
        SubCellInst_LFInst_6_LFInst_2_n15) );
  NOR2_X1 SubCellInst_LFInst_6_LFInst_3_U4 ( .A1(PermutationOutput[25]), .A2(
        PermutationOutput[26]), .ZN(SubCellInst_LFInst_6_LFInst_3_n8) );
  NOR2_X1 SubCellInst_LFInst_6_LFInst_3_U3 ( .A1(PermutationOutput[27]), .A2(
        SubCellInst_LFInst_6_LFInst_3_n7), .ZN(
        SubCellInst_LFInst_6_LFInst_3_n9) );
  AND2_X1 SubCellInst_LFInst_6_LFInst_3_U2 ( .A1(PermutationOutput[25]), .A2(
        PermutationOutput[24]), .ZN(SubCellInst_LFInst_6_LFInst_3_n7) );
  OR2_X1 SubCellInst_LFInst_6_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_6_LFInst_3_n9), .A2(
        SubCellInst_LFInst_6_LFInst_3_n8), .ZN(MCOutput2[27]) );
  NOR2_X1 SubCellInst_LFInst_7_LFInst_0_U6 ( .A1(
        SubCellInst_LFInst_7_LFInst_0_n15), .A2(
        SubCellInst_LFInst_7_LFInst_0_n14), .ZN(MCOutput2[28]) );
  AND2_X1 SubCellInst_LFInst_7_LFInst_0_U5 ( .A1(PermutationOutput[31]), .A2(
        PermutationOutput[30]), .ZN(SubCellInst_LFInst_7_LFInst_0_n14) );
  NOR2_X1 SubCellInst_LFInst_7_LFInst_0_U4 ( .A1(PermutationOutput[29]), .A2(
        SubCellInst_LFInst_7_LFInst_0_n13), .ZN(
        SubCellInst_LFInst_7_LFInst_0_n15) );
  NOR2_X1 SubCellInst_LFInst_7_LFInst_0_U3 ( .A1(
        SubCellInst_LFInst_7_LFInst_0_n12), .A2(
        SubCellInst_LFInst_7_LFInst_0_n11), .ZN(
        SubCellInst_LFInst_7_LFInst_0_n13) );
  NOR2_X1 SubCellInst_LFInst_7_LFInst_0_U2 ( .A1(PermutationOutput[31]), .A2(
        PermutationOutput[30]), .ZN(SubCellInst_LFInst_7_LFInst_0_n11) );
  INV_X1 SubCellInst_LFInst_7_LFInst_0_U1 ( .A(PermutationOutput[28]), .ZN(
        SubCellInst_LFInst_7_LFInst_0_n12) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_1_U4 ( .A1(
        SubCellInst_LFInst_7_LFInst_1_n9), .A2(
        SubCellInst_LFInst_7_LFInst_1_n8), .ZN(MCOutput2[29]) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_1_U3 ( .A1(PermutationOutput[28]), .A2(
        PermutationOutput[30]), .ZN(SubCellInst_LFInst_7_LFInst_1_n8) );
  OR2_X1 SubCellInst_LFInst_7_LFInst_1_U2 ( .A1(PermutationOutput[31]), .A2(
        SubCellInst_LFInst_7_LFInst_1_n7), .ZN(
        SubCellInst_LFInst_7_LFInst_1_n9) );
  NOR2_X1 SubCellInst_LFInst_7_LFInst_1_U1 ( .A1(PermutationOutput[28]), .A2(
        PermutationOutput[30]), .ZN(SubCellInst_LFInst_7_LFInst_1_n7) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_2_U6 ( .A1(
        SubCellInst_LFInst_7_LFInst_2_n18), .A2(
        SubCellInst_LFInst_7_LFInst_2_n17), .ZN(MCOutput2[30]) );
  OR2_X1 SubCellInst_LFInst_7_LFInst_2_U5 ( .A1(PermutationOutput[28]), .A2(
        PermutationOutput[31]), .ZN(SubCellInst_LFInst_7_LFInst_2_n17) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_2_U4 ( .A1(PermutationOutput[29]), .A2(
        SubCellInst_LFInst_7_LFInst_2_n16), .ZN(
        SubCellInst_LFInst_7_LFInst_2_n18) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_2_U3 ( .A1(
        SubCellInst_LFInst_7_LFInst_2_n15), .A2(
        SubCellInst_LFInst_7_LFInst_2_n14), .ZN(
        SubCellInst_LFInst_7_LFInst_2_n16) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_2_U2 ( .A1(PermutationOutput[28]), .A2(
        PermutationOutput[31]), .ZN(SubCellInst_LFInst_7_LFInst_2_n14) );
  INV_X1 SubCellInst_LFInst_7_LFInst_2_U1 ( .A(PermutationOutput[30]), .ZN(
        SubCellInst_LFInst_7_LFInst_2_n15) );
  NOR2_X1 SubCellInst_LFInst_7_LFInst_3_U4 ( .A1(PermutationOutput[29]), .A2(
        PermutationOutput[30]), .ZN(SubCellInst_LFInst_7_LFInst_3_n8) );
  NOR2_X1 SubCellInst_LFInst_7_LFInst_3_U3 ( .A1(PermutationOutput[31]), .A2(
        SubCellInst_LFInst_7_LFInst_3_n7), .ZN(
        SubCellInst_LFInst_7_LFInst_3_n9) );
  AND2_X1 SubCellInst_LFInst_7_LFInst_3_U2 ( .A1(PermutationOutput[29]), .A2(
        PermutationOutput[28]), .ZN(SubCellInst_LFInst_7_LFInst_3_n7) );
  OR2_X1 SubCellInst_LFInst_7_LFInst_3_U1 ( .A1(
        SubCellInst_LFInst_7_LFInst_3_n9), .A2(
        SubCellInst_LFInst_7_LFInst_3_n8), .ZN(MCOutput2[31]) );
  NOR2_X1 SubCellInst_LFInst_8_LFInst_0_U6 ( .A1(
        SubCellInst_LFInst_8_LFInst_0_n15), .A2(
        SubCellInst_LFInst_8_LFInst_0_n14), .ZN(SboxOut[32]) );
  AND2_X1 SubCellInst_LFInst_8_LFInst_0_U5 ( .A1(PermutationOutput[35]), .A2(
        PermutationOutput[34]), .ZN(SubCellInst_LFInst_8_LFInst_0_n14) );
  NOR2_X1 SubCellInst_LFInst_8_LFInst_0_U4 ( .A1(PermutationOutput[33]), .A2(
        SubCellInst_LFInst_8_LFInst_0_n13), .ZN(
        SubCellInst_LFInst_8_LFInst_0_n15) );
  NOR2_X1 SubCellInst_LFInst_8_LFInst_0_U3 ( .A1(
        SubCellInst_LFInst_8_LFInst_0_n12), .A2(
        SubCellInst_LFInst_8_LFInst_0_n11), .ZN(
        SubCellInst_LFInst_8_LFInst_0_n13) );
  NOR2_X1 SubCellInst_LFInst_8_LFInst_0_U2 ( .A1(PermutationOutput[35]), .A2(
        PermutationOutput[34]), .ZN(SubCellInst_LFInst_8_LFInst_0_n11) );
  INV_X1 SubCellInst_LFInst_8_LFInst_0_U1 ( .A(PermutationOutput[32]), .ZN(
        SubCellInst_LFInst_8_LFInst_0_n12) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_1_U4 ( .A1(
        SubCellInst_LFInst_8_LFInst_1_n9), .A2(
        SubCellInst_LFInst_8_LFInst_1_n8), .ZN(SboxOut[33]) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_1_U3 ( .A1(PermutationOutput[32]), .A2(
        PermutationOutput[34]), .ZN(SubCellInst_LFInst_8_LFInst_1_n8) );
  OR2_X1 SubCellInst_LFInst_8_LFInst_1_U2 ( .A1(PermutationOutput[35]), .A2(
        SubCellInst_LFInst_8_LFInst_1_n7), .ZN(
        SubCellInst_LFInst_8_LFInst_1_n9) );
  NOR2_X1 SubCellInst_LFInst_8_LFInst_1_U1 ( .A1(PermutationOutput[32]), .A2(
        PermutationOutput[34]), .ZN(SubCellInst_LFInst_8_LFInst_1_n7) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_2_U6 ( .A1(
        SubCellInst_LFInst_8_LFInst_2_n18), .A2(
        SubCellInst_LFInst_8_LFInst_2_n17), .ZN(SboxOut[34]) );
  OR2_X1 SubCellInst_LFInst_8_LFInst_2_U5 ( .A1(PermutationOutput[32]), .A2(
        PermutationOutput[35]), .ZN(SubCellInst_LFInst_8_LFInst_2_n17) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_2_U4 ( .A1(PermutationOutput[33]), .A2(
        SubCellInst_LFInst_8_LFInst_2_n16), .ZN(
        SubCellInst_LFInst_8_LFInst_2_n18) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_2_U3 ( .A1(
        SubCellInst_LFInst_8_LFInst_2_n15), .A2(
        SubCellInst_LFInst_8_LFInst_2_n14), .ZN(
        SubCellInst_LFInst_8_LFInst_2_n16) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_2_U2 ( .A1(PermutationOutput[32]), .A2(
        PermutationOutput[35]), .ZN(SubCellInst_LFInst_8_LFInst_2_n14) );
  INV_X1 SubCellInst_LFInst_8_LFInst_2_U1 ( .A(PermutationOutput[34]), .ZN(
        SubCellInst_LFInst_8_LFInst_2_n15) );
  OR2_X1 SubCellInst_LFInst_8_LFInst_3_U4 ( .A1(
        SubCellInst_LFInst_8_LFInst_3_n9), .A2(
        SubCellInst_LFInst_8_LFInst_3_n8), .ZN(SboxOut[35]) );
  NOR2_X1 SubCellInst_LFInst_8_LFInst_3_U3 ( .A1(PermutationOutput[33]), .A2(
        PermutationOutput[34]), .ZN(SubCellInst_LFInst_8_LFInst_3_n8) );
  NOR2_X1 SubCellInst_LFInst_8_LFInst_3_U2 ( .A1(PermutationOutput[35]), .A2(
        SubCellInst_LFInst_8_LFInst_3_n7), .ZN(
        SubCellInst_LFInst_8_LFInst_3_n9) );
  AND2_X1 SubCellInst_LFInst_8_LFInst_3_U1 ( .A1(PermutationOutput[33]), .A2(
        PermutationOutput[32]), .ZN(SubCellInst_LFInst_8_LFInst_3_n7) );
  NOR2_X1 SubCellInst_LFInst_9_LFInst_0_U6 ( .A1(
        SubCellInst_LFInst_9_LFInst_0_n15), .A2(
        SubCellInst_LFInst_9_LFInst_0_n14), .ZN(SboxOut[36]) );
  AND2_X1 SubCellInst_LFInst_9_LFInst_0_U5 ( .A1(PermutationOutput[39]), .A2(
        PermutationOutput[38]), .ZN(SubCellInst_LFInst_9_LFInst_0_n14) );
  NOR2_X1 SubCellInst_LFInst_9_LFInst_0_U4 ( .A1(PermutationOutput[37]), .A2(
        SubCellInst_LFInst_9_LFInst_0_n13), .ZN(
        SubCellInst_LFInst_9_LFInst_0_n15) );
  NOR2_X1 SubCellInst_LFInst_9_LFInst_0_U3 ( .A1(
        SubCellInst_LFInst_9_LFInst_0_n12), .A2(
        SubCellInst_LFInst_9_LFInst_0_n11), .ZN(
        SubCellInst_LFInst_9_LFInst_0_n13) );
  NOR2_X1 SubCellInst_LFInst_9_LFInst_0_U2 ( .A1(PermutationOutput[39]), .A2(
        PermutationOutput[38]), .ZN(SubCellInst_LFInst_9_LFInst_0_n11) );
  INV_X1 SubCellInst_LFInst_9_LFInst_0_U1 ( .A(PermutationOutput[36]), .ZN(
        SubCellInst_LFInst_9_LFInst_0_n12) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_1_U4 ( .A1(
        SubCellInst_LFInst_9_LFInst_1_n9), .A2(
        SubCellInst_LFInst_9_LFInst_1_n8), .ZN(SboxOut[37]) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_1_U3 ( .A1(PermutationOutput[36]), .A2(
        PermutationOutput[38]), .ZN(SubCellInst_LFInst_9_LFInst_1_n8) );
  OR2_X1 SubCellInst_LFInst_9_LFInst_1_U2 ( .A1(PermutationOutput[39]), .A2(
        SubCellInst_LFInst_9_LFInst_1_n7), .ZN(
        SubCellInst_LFInst_9_LFInst_1_n9) );
  NOR2_X1 SubCellInst_LFInst_9_LFInst_1_U1 ( .A1(PermutationOutput[36]), .A2(
        PermutationOutput[38]), .ZN(SubCellInst_LFInst_9_LFInst_1_n7) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_2_U6 ( .A1(
        SubCellInst_LFInst_9_LFInst_2_n18), .A2(
        SubCellInst_LFInst_9_LFInst_2_n17), .ZN(SboxOut[38]) );
  OR2_X1 SubCellInst_LFInst_9_LFInst_2_U5 ( .A1(PermutationOutput[36]), .A2(
        PermutationOutput[39]), .ZN(SubCellInst_LFInst_9_LFInst_2_n17) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_2_U4 ( .A1(PermutationOutput[37]), .A2(
        SubCellInst_LFInst_9_LFInst_2_n16), .ZN(
        SubCellInst_LFInst_9_LFInst_2_n18) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_2_U3 ( .A1(
        SubCellInst_LFInst_9_LFInst_2_n15), .A2(
        SubCellInst_LFInst_9_LFInst_2_n14), .ZN(
        SubCellInst_LFInst_9_LFInst_2_n16) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_2_U2 ( .A1(PermutationOutput[36]), .A2(
        PermutationOutput[39]), .ZN(SubCellInst_LFInst_9_LFInst_2_n14) );
  INV_X1 SubCellInst_LFInst_9_LFInst_2_U1 ( .A(PermutationOutput[38]), .ZN(
        SubCellInst_LFInst_9_LFInst_2_n15) );
  OR2_X1 SubCellInst_LFInst_9_LFInst_3_U4 ( .A1(
        SubCellInst_LFInst_9_LFInst_3_n9), .A2(
        SubCellInst_LFInst_9_LFInst_3_n8), .ZN(SboxOut[39]) );
  NOR2_X1 SubCellInst_LFInst_9_LFInst_3_U3 ( .A1(PermutationOutput[37]), .A2(
        PermutationOutput[38]), .ZN(SubCellInst_LFInst_9_LFInst_3_n8) );
  NOR2_X1 SubCellInst_LFInst_9_LFInst_3_U2 ( .A1(PermutationOutput[39]), .A2(
        SubCellInst_LFInst_9_LFInst_3_n7), .ZN(
        SubCellInst_LFInst_9_LFInst_3_n9) );
  AND2_X1 SubCellInst_LFInst_9_LFInst_3_U1 ( .A1(PermutationOutput[37]), .A2(
        PermutationOutput[36]), .ZN(SubCellInst_LFInst_9_LFInst_3_n7) );
  NOR2_X1 SubCellInst_LFInst_10_LFInst_0_U6 ( .A1(
        SubCellInst_LFInst_10_LFInst_0_n15), .A2(
        SubCellInst_LFInst_10_LFInst_0_n14), .ZN(SboxOut[40]) );
  AND2_X1 SubCellInst_LFInst_10_LFInst_0_U5 ( .A1(PermutationOutput[43]), .A2(
        PermutationOutput[42]), .ZN(SubCellInst_LFInst_10_LFInst_0_n14) );
  NOR2_X1 SubCellInst_LFInst_10_LFInst_0_U4 ( .A1(PermutationOutput[41]), .A2(
        SubCellInst_LFInst_10_LFInst_0_n13), .ZN(
        SubCellInst_LFInst_10_LFInst_0_n15) );
  NOR2_X1 SubCellInst_LFInst_10_LFInst_0_U3 ( .A1(
        SubCellInst_LFInst_10_LFInst_0_n12), .A2(
        SubCellInst_LFInst_10_LFInst_0_n11), .ZN(
        SubCellInst_LFInst_10_LFInst_0_n13) );
  NOR2_X1 SubCellInst_LFInst_10_LFInst_0_U2 ( .A1(PermutationOutput[43]), .A2(
        PermutationOutput[42]), .ZN(SubCellInst_LFInst_10_LFInst_0_n11) );
  INV_X1 SubCellInst_LFInst_10_LFInst_0_U1 ( .A(PermutationOutput[40]), .ZN(
        SubCellInst_LFInst_10_LFInst_0_n12) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_1_U4 ( .A1(
        SubCellInst_LFInst_10_LFInst_1_n9), .A2(
        SubCellInst_LFInst_10_LFInst_1_n8), .ZN(SboxOut[41]) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_1_U3 ( .A1(PermutationOutput[40]), 
        .A2(PermutationOutput[42]), .ZN(SubCellInst_LFInst_10_LFInst_1_n8) );
  OR2_X1 SubCellInst_LFInst_10_LFInst_1_U2 ( .A1(PermutationOutput[43]), .A2(
        SubCellInst_LFInst_10_LFInst_1_n7), .ZN(
        SubCellInst_LFInst_10_LFInst_1_n9) );
  NOR2_X1 SubCellInst_LFInst_10_LFInst_1_U1 ( .A1(PermutationOutput[40]), .A2(
        PermutationOutput[42]), .ZN(SubCellInst_LFInst_10_LFInst_1_n7) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_2_U6 ( .A1(
        SubCellInst_LFInst_10_LFInst_2_n18), .A2(
        SubCellInst_LFInst_10_LFInst_2_n17), .ZN(SboxOut[42]) );
  OR2_X1 SubCellInst_LFInst_10_LFInst_2_U5 ( .A1(PermutationOutput[40]), .A2(
        PermutationOutput[43]), .ZN(SubCellInst_LFInst_10_LFInst_2_n17) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_2_U4 ( .A1(PermutationOutput[41]), 
        .A2(SubCellInst_LFInst_10_LFInst_2_n16), .ZN(
        SubCellInst_LFInst_10_LFInst_2_n18) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_2_U3 ( .A1(
        SubCellInst_LFInst_10_LFInst_2_n15), .A2(
        SubCellInst_LFInst_10_LFInst_2_n14), .ZN(
        SubCellInst_LFInst_10_LFInst_2_n16) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_2_U2 ( .A1(PermutationOutput[40]), 
        .A2(PermutationOutput[43]), .ZN(SubCellInst_LFInst_10_LFInst_2_n14) );
  INV_X1 SubCellInst_LFInst_10_LFInst_2_U1 ( .A(PermutationOutput[42]), .ZN(
        SubCellInst_LFInst_10_LFInst_2_n15) );
  OR2_X1 SubCellInst_LFInst_10_LFInst_3_U4 ( .A1(
        SubCellInst_LFInst_10_LFInst_3_n9), .A2(
        SubCellInst_LFInst_10_LFInst_3_n8), .ZN(SboxOut[43]) );
  NOR2_X1 SubCellInst_LFInst_10_LFInst_3_U3 ( .A1(PermutationOutput[41]), .A2(
        PermutationOutput[42]), .ZN(SubCellInst_LFInst_10_LFInst_3_n8) );
  NOR2_X1 SubCellInst_LFInst_10_LFInst_3_U2 ( .A1(PermutationOutput[43]), .A2(
        SubCellInst_LFInst_10_LFInst_3_n7), .ZN(
        SubCellInst_LFInst_10_LFInst_3_n9) );
  AND2_X1 SubCellInst_LFInst_10_LFInst_3_U1 ( .A1(PermutationOutput[41]), .A2(
        PermutationOutput[40]), .ZN(SubCellInst_LFInst_10_LFInst_3_n7) );
  NOR2_X1 SubCellInst_LFInst_11_LFInst_0_U6 ( .A1(
        SubCellInst_LFInst_11_LFInst_0_n15), .A2(
        SubCellInst_LFInst_11_LFInst_0_n14), .ZN(SboxOut[44]) );
  AND2_X1 SubCellInst_LFInst_11_LFInst_0_U5 ( .A1(PermutationOutput[47]), .A2(
        PermutationOutput[46]), .ZN(SubCellInst_LFInst_11_LFInst_0_n14) );
  NOR2_X1 SubCellInst_LFInst_11_LFInst_0_U4 ( .A1(PermutationOutput[45]), .A2(
        SubCellInst_LFInst_11_LFInst_0_n13), .ZN(
        SubCellInst_LFInst_11_LFInst_0_n15) );
  NOR2_X1 SubCellInst_LFInst_11_LFInst_0_U3 ( .A1(
        SubCellInst_LFInst_11_LFInst_0_n12), .A2(
        SubCellInst_LFInst_11_LFInst_0_n11), .ZN(
        SubCellInst_LFInst_11_LFInst_0_n13) );
  NOR2_X1 SubCellInst_LFInst_11_LFInst_0_U2 ( .A1(PermutationOutput[47]), .A2(
        PermutationOutput[46]), .ZN(SubCellInst_LFInst_11_LFInst_0_n11) );
  INV_X1 SubCellInst_LFInst_11_LFInst_0_U1 ( .A(PermutationOutput[44]), .ZN(
        SubCellInst_LFInst_11_LFInst_0_n12) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_1_U4 ( .A1(
        SubCellInst_LFInst_11_LFInst_1_n9), .A2(
        SubCellInst_LFInst_11_LFInst_1_n8), .ZN(SboxOut[45]) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_1_U3 ( .A1(PermutationOutput[44]), 
        .A2(PermutationOutput[46]), .ZN(SubCellInst_LFInst_11_LFInst_1_n8) );
  OR2_X1 SubCellInst_LFInst_11_LFInst_1_U2 ( .A1(PermutationOutput[47]), .A2(
        SubCellInst_LFInst_11_LFInst_1_n7), .ZN(
        SubCellInst_LFInst_11_LFInst_1_n9) );
  NOR2_X1 SubCellInst_LFInst_11_LFInst_1_U1 ( .A1(PermutationOutput[44]), .A2(
        PermutationOutput[46]), .ZN(SubCellInst_LFInst_11_LFInst_1_n7) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_2_U6 ( .A1(
        SubCellInst_LFInst_11_LFInst_2_n18), .A2(
        SubCellInst_LFInst_11_LFInst_2_n17), .ZN(SboxOut[46]) );
  OR2_X1 SubCellInst_LFInst_11_LFInst_2_U5 ( .A1(PermutationOutput[44]), .A2(
        PermutationOutput[47]), .ZN(SubCellInst_LFInst_11_LFInst_2_n17) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_2_U4 ( .A1(PermutationOutput[45]), 
        .A2(SubCellInst_LFInst_11_LFInst_2_n16), .ZN(
        SubCellInst_LFInst_11_LFInst_2_n18) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_2_U3 ( .A1(
        SubCellInst_LFInst_11_LFInst_2_n15), .A2(
        SubCellInst_LFInst_11_LFInst_2_n14), .ZN(
        SubCellInst_LFInst_11_LFInst_2_n16) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_2_U2 ( .A1(PermutationOutput[44]), 
        .A2(PermutationOutput[47]), .ZN(SubCellInst_LFInst_11_LFInst_2_n14) );
  INV_X1 SubCellInst_LFInst_11_LFInst_2_U1 ( .A(PermutationOutput[46]), .ZN(
        SubCellInst_LFInst_11_LFInst_2_n15) );
  OR2_X1 SubCellInst_LFInst_11_LFInst_3_U4 ( .A1(
        SubCellInst_LFInst_11_LFInst_3_n9), .A2(
        SubCellInst_LFInst_11_LFInst_3_n8), .ZN(SboxOut[47]) );
  NOR2_X1 SubCellInst_LFInst_11_LFInst_3_U3 ( .A1(PermutationOutput[45]), .A2(
        PermutationOutput[46]), .ZN(SubCellInst_LFInst_11_LFInst_3_n8) );
  NOR2_X1 SubCellInst_LFInst_11_LFInst_3_U2 ( .A1(PermutationOutput[47]), .A2(
        SubCellInst_LFInst_11_LFInst_3_n7), .ZN(
        SubCellInst_LFInst_11_LFInst_3_n9) );
  AND2_X1 SubCellInst_LFInst_11_LFInst_3_U1 ( .A1(PermutationOutput[45]), .A2(
        PermutationOutput[44]), .ZN(SubCellInst_LFInst_11_LFInst_3_n7) );
  NOR2_X1 SubCellInst_LFInst_12_LFInst_0_U6 ( .A1(
        SubCellInst_LFInst_12_LFInst_0_n15), .A2(
        SubCellInst_LFInst_12_LFInst_0_n14), .ZN(SboxOut[48]) );
  AND2_X1 SubCellInst_LFInst_12_LFInst_0_U5 ( .A1(PermutationOutput[51]), .A2(
        PermutationOutput[50]), .ZN(SubCellInst_LFInst_12_LFInst_0_n14) );
  NOR2_X1 SubCellInst_LFInst_12_LFInst_0_U4 ( .A1(PermutationOutput[49]), .A2(
        SubCellInst_LFInst_12_LFInst_0_n13), .ZN(
        SubCellInst_LFInst_12_LFInst_0_n15) );
  NOR2_X1 SubCellInst_LFInst_12_LFInst_0_U3 ( .A1(
        SubCellInst_LFInst_12_LFInst_0_n12), .A2(
        SubCellInst_LFInst_12_LFInst_0_n11), .ZN(
        SubCellInst_LFInst_12_LFInst_0_n13) );
  NOR2_X1 SubCellInst_LFInst_12_LFInst_0_U2 ( .A1(PermutationOutput[51]), .A2(
        PermutationOutput[50]), .ZN(SubCellInst_LFInst_12_LFInst_0_n11) );
  INV_X1 SubCellInst_LFInst_12_LFInst_0_U1 ( .A(PermutationOutput[48]), .ZN(
        SubCellInst_LFInst_12_LFInst_0_n12) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_1_U4 ( .A1(
        SubCellInst_LFInst_12_LFInst_1_n9), .A2(
        SubCellInst_LFInst_12_LFInst_1_n8), .ZN(SboxOut[49]) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_1_U3 ( .A1(PermutationOutput[48]), 
        .A2(PermutationOutput[50]), .ZN(SubCellInst_LFInst_12_LFInst_1_n8) );
  OR2_X1 SubCellInst_LFInst_12_LFInst_1_U2 ( .A1(PermutationOutput[51]), .A2(
        SubCellInst_LFInst_12_LFInst_1_n7), .ZN(
        SubCellInst_LFInst_12_LFInst_1_n9) );
  NOR2_X1 SubCellInst_LFInst_12_LFInst_1_U1 ( .A1(PermutationOutput[48]), .A2(
        PermutationOutput[50]), .ZN(SubCellInst_LFInst_12_LFInst_1_n7) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_2_U6 ( .A1(
        SubCellInst_LFInst_12_LFInst_2_n18), .A2(
        SubCellInst_LFInst_12_LFInst_2_n17), .ZN(SboxOut[50]) );
  OR2_X1 SubCellInst_LFInst_12_LFInst_2_U5 ( .A1(PermutationOutput[48]), .A2(
        PermutationOutput[51]), .ZN(SubCellInst_LFInst_12_LFInst_2_n17) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_2_U4 ( .A1(PermutationOutput[49]), 
        .A2(SubCellInst_LFInst_12_LFInst_2_n16), .ZN(
        SubCellInst_LFInst_12_LFInst_2_n18) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_2_U3 ( .A1(
        SubCellInst_LFInst_12_LFInst_2_n15), .A2(
        SubCellInst_LFInst_12_LFInst_2_n14), .ZN(
        SubCellInst_LFInst_12_LFInst_2_n16) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_2_U2 ( .A1(PermutationOutput[48]), 
        .A2(PermutationOutput[51]), .ZN(SubCellInst_LFInst_12_LFInst_2_n14) );
  INV_X1 SubCellInst_LFInst_12_LFInst_2_U1 ( .A(PermutationOutput[50]), .ZN(
        SubCellInst_LFInst_12_LFInst_2_n15) );
  OR2_X1 SubCellInst_LFInst_12_LFInst_3_U4 ( .A1(
        SubCellInst_LFInst_12_LFInst_3_n9), .A2(
        SubCellInst_LFInst_12_LFInst_3_n8), .ZN(SboxOut[51]) );
  NOR2_X1 SubCellInst_LFInst_12_LFInst_3_U3 ( .A1(PermutationOutput[49]), .A2(
        PermutationOutput[50]), .ZN(SubCellInst_LFInst_12_LFInst_3_n8) );
  NOR2_X1 SubCellInst_LFInst_12_LFInst_3_U2 ( .A1(PermutationOutput[51]), .A2(
        SubCellInst_LFInst_12_LFInst_3_n7), .ZN(
        SubCellInst_LFInst_12_LFInst_3_n9) );
  AND2_X1 SubCellInst_LFInst_12_LFInst_3_U1 ( .A1(PermutationOutput[49]), .A2(
        PermutationOutput[48]), .ZN(SubCellInst_LFInst_12_LFInst_3_n7) );
  NOR2_X1 SubCellInst_LFInst_13_LFInst_0_U6 ( .A1(
        SubCellInst_LFInst_13_LFInst_0_n15), .A2(
        SubCellInst_LFInst_13_LFInst_0_n14), .ZN(SboxOut[52]) );
  AND2_X1 SubCellInst_LFInst_13_LFInst_0_U5 ( .A1(PermutationOutput[55]), .A2(
        PermutationOutput[54]), .ZN(SubCellInst_LFInst_13_LFInst_0_n14) );
  NOR2_X1 SubCellInst_LFInst_13_LFInst_0_U4 ( .A1(PermutationOutput[53]), .A2(
        SubCellInst_LFInst_13_LFInst_0_n13), .ZN(
        SubCellInst_LFInst_13_LFInst_0_n15) );
  NOR2_X1 SubCellInst_LFInst_13_LFInst_0_U3 ( .A1(
        SubCellInst_LFInst_13_LFInst_0_n12), .A2(
        SubCellInst_LFInst_13_LFInst_0_n11), .ZN(
        SubCellInst_LFInst_13_LFInst_0_n13) );
  NOR2_X1 SubCellInst_LFInst_13_LFInst_0_U2 ( .A1(PermutationOutput[55]), .A2(
        PermutationOutput[54]), .ZN(SubCellInst_LFInst_13_LFInst_0_n11) );
  INV_X1 SubCellInst_LFInst_13_LFInst_0_U1 ( .A(PermutationOutput[52]), .ZN(
        SubCellInst_LFInst_13_LFInst_0_n12) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_1_U4 ( .A1(
        SubCellInst_LFInst_13_LFInst_1_n9), .A2(
        SubCellInst_LFInst_13_LFInst_1_n8), .ZN(SboxOut[53]) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_1_U3 ( .A1(PermutationOutput[52]), 
        .A2(PermutationOutput[54]), .ZN(SubCellInst_LFInst_13_LFInst_1_n8) );
  OR2_X1 SubCellInst_LFInst_13_LFInst_1_U2 ( .A1(PermutationOutput[55]), .A2(
        SubCellInst_LFInst_13_LFInst_1_n7), .ZN(
        SubCellInst_LFInst_13_LFInst_1_n9) );
  NOR2_X1 SubCellInst_LFInst_13_LFInst_1_U1 ( .A1(PermutationOutput[52]), .A2(
        PermutationOutput[54]), .ZN(SubCellInst_LFInst_13_LFInst_1_n7) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_2_U6 ( .A1(
        SubCellInst_LFInst_13_LFInst_2_n18), .A2(
        SubCellInst_LFInst_13_LFInst_2_n17), .ZN(SboxOut[54]) );
  OR2_X1 SubCellInst_LFInst_13_LFInst_2_U5 ( .A1(PermutationOutput[52]), .A2(
        PermutationOutput[55]), .ZN(SubCellInst_LFInst_13_LFInst_2_n17) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_2_U4 ( .A1(PermutationOutput[53]), 
        .A2(SubCellInst_LFInst_13_LFInst_2_n16), .ZN(
        SubCellInst_LFInst_13_LFInst_2_n18) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_2_U3 ( .A1(
        SubCellInst_LFInst_13_LFInst_2_n15), .A2(
        SubCellInst_LFInst_13_LFInst_2_n14), .ZN(
        SubCellInst_LFInst_13_LFInst_2_n16) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_2_U2 ( .A1(PermutationOutput[52]), 
        .A2(PermutationOutput[55]), .ZN(SubCellInst_LFInst_13_LFInst_2_n14) );
  INV_X1 SubCellInst_LFInst_13_LFInst_2_U1 ( .A(PermutationOutput[54]), .ZN(
        SubCellInst_LFInst_13_LFInst_2_n15) );
  OR2_X1 SubCellInst_LFInst_13_LFInst_3_U4 ( .A1(
        SubCellInst_LFInst_13_LFInst_3_n9), .A2(
        SubCellInst_LFInst_13_LFInst_3_n8), .ZN(SboxOut[55]) );
  NOR2_X1 SubCellInst_LFInst_13_LFInst_3_U3 ( .A1(PermutationOutput[53]), .A2(
        PermutationOutput[54]), .ZN(SubCellInst_LFInst_13_LFInst_3_n8) );
  NOR2_X1 SubCellInst_LFInst_13_LFInst_3_U2 ( .A1(PermutationOutput[55]), .A2(
        SubCellInst_LFInst_13_LFInst_3_n7), .ZN(
        SubCellInst_LFInst_13_LFInst_3_n9) );
  AND2_X1 SubCellInst_LFInst_13_LFInst_3_U1 ( .A1(PermutationOutput[53]), .A2(
        PermutationOutput[52]), .ZN(SubCellInst_LFInst_13_LFInst_3_n7) );
  NOR2_X1 SubCellInst_LFInst_14_LFInst_0_U6 ( .A1(
        SubCellInst_LFInst_14_LFInst_0_n15), .A2(
        SubCellInst_LFInst_14_LFInst_0_n14), .ZN(SboxOut[56]) );
  AND2_X1 SubCellInst_LFInst_14_LFInst_0_U5 ( .A1(PermutationOutput[59]), .A2(
        PermutationOutput[58]), .ZN(SubCellInst_LFInst_14_LFInst_0_n14) );
  NOR2_X1 SubCellInst_LFInst_14_LFInst_0_U4 ( .A1(PermutationOutput[57]), .A2(
        SubCellInst_LFInst_14_LFInst_0_n13), .ZN(
        SubCellInst_LFInst_14_LFInst_0_n15) );
  NOR2_X1 SubCellInst_LFInst_14_LFInst_0_U3 ( .A1(
        SubCellInst_LFInst_14_LFInst_0_n12), .A2(
        SubCellInst_LFInst_14_LFInst_0_n11), .ZN(
        SubCellInst_LFInst_14_LFInst_0_n13) );
  NOR2_X1 SubCellInst_LFInst_14_LFInst_0_U2 ( .A1(PermutationOutput[59]), .A2(
        PermutationOutput[58]), .ZN(SubCellInst_LFInst_14_LFInst_0_n11) );
  INV_X1 SubCellInst_LFInst_14_LFInst_0_U1 ( .A(PermutationOutput[56]), .ZN(
        SubCellInst_LFInst_14_LFInst_0_n12) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_1_U4 ( .A1(
        SubCellInst_LFInst_14_LFInst_1_n9), .A2(
        SubCellInst_LFInst_14_LFInst_1_n8), .ZN(SboxOut[57]) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_1_U3 ( .A1(PermutationOutput[56]), 
        .A2(PermutationOutput[58]), .ZN(SubCellInst_LFInst_14_LFInst_1_n8) );
  OR2_X1 SubCellInst_LFInst_14_LFInst_1_U2 ( .A1(PermutationOutput[59]), .A2(
        SubCellInst_LFInst_14_LFInst_1_n7), .ZN(
        SubCellInst_LFInst_14_LFInst_1_n9) );
  NOR2_X1 SubCellInst_LFInst_14_LFInst_1_U1 ( .A1(PermutationOutput[56]), .A2(
        PermutationOutput[58]), .ZN(SubCellInst_LFInst_14_LFInst_1_n7) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_2_U6 ( .A1(
        SubCellInst_LFInst_14_LFInst_2_n18), .A2(
        SubCellInst_LFInst_14_LFInst_2_n17), .ZN(SboxOut[58]) );
  OR2_X1 SubCellInst_LFInst_14_LFInst_2_U5 ( .A1(PermutationOutput[56]), .A2(
        PermutationOutput[59]), .ZN(SubCellInst_LFInst_14_LFInst_2_n17) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_2_U4 ( .A1(PermutationOutput[57]), 
        .A2(SubCellInst_LFInst_14_LFInst_2_n16), .ZN(
        SubCellInst_LFInst_14_LFInst_2_n18) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_2_U3 ( .A1(
        SubCellInst_LFInst_14_LFInst_2_n15), .A2(
        SubCellInst_LFInst_14_LFInst_2_n14), .ZN(
        SubCellInst_LFInst_14_LFInst_2_n16) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_2_U2 ( .A1(PermutationOutput[56]), 
        .A2(PermutationOutput[59]), .ZN(SubCellInst_LFInst_14_LFInst_2_n14) );
  INV_X1 SubCellInst_LFInst_14_LFInst_2_U1 ( .A(PermutationOutput[58]), .ZN(
        SubCellInst_LFInst_14_LFInst_2_n15) );
  OR2_X1 SubCellInst_LFInst_14_LFInst_3_U4 ( .A1(
        SubCellInst_LFInst_14_LFInst_3_n9), .A2(
        SubCellInst_LFInst_14_LFInst_3_n8), .ZN(SboxOut[59]) );
  NOR2_X1 SubCellInst_LFInst_14_LFInst_3_U3 ( .A1(PermutationOutput[57]), .A2(
        PermutationOutput[58]), .ZN(SubCellInst_LFInst_14_LFInst_3_n8) );
  NOR2_X1 SubCellInst_LFInst_14_LFInst_3_U2 ( .A1(PermutationOutput[59]), .A2(
        SubCellInst_LFInst_14_LFInst_3_n7), .ZN(
        SubCellInst_LFInst_14_LFInst_3_n9) );
  AND2_X1 SubCellInst_LFInst_14_LFInst_3_U1 ( .A1(PermutationOutput[57]), .A2(
        PermutationOutput[56]), .ZN(SubCellInst_LFInst_14_LFInst_3_n7) );
  NOR2_X1 SubCellInst_LFInst_15_LFInst_0_U6 ( .A1(
        SubCellInst_LFInst_15_LFInst_0_n15), .A2(
        SubCellInst_LFInst_15_LFInst_0_n14), .ZN(SboxOut[60]) );
  AND2_X1 SubCellInst_LFInst_15_LFInst_0_U5 ( .A1(PermutationOutput[63]), .A2(
        PermutationOutput[62]), .ZN(SubCellInst_LFInst_15_LFInst_0_n14) );
  NOR2_X1 SubCellInst_LFInst_15_LFInst_0_U4 ( .A1(PermutationOutput[61]), .A2(
        SubCellInst_LFInst_15_LFInst_0_n13), .ZN(
        SubCellInst_LFInst_15_LFInst_0_n15) );
  NOR2_X1 SubCellInst_LFInst_15_LFInst_0_U3 ( .A1(
        SubCellInst_LFInst_15_LFInst_0_n12), .A2(
        SubCellInst_LFInst_15_LFInst_0_n11), .ZN(
        SubCellInst_LFInst_15_LFInst_0_n13) );
  NOR2_X1 SubCellInst_LFInst_15_LFInst_0_U2 ( .A1(PermutationOutput[63]), .A2(
        PermutationOutput[62]), .ZN(SubCellInst_LFInst_15_LFInst_0_n11) );
  INV_X1 SubCellInst_LFInst_15_LFInst_0_U1 ( .A(PermutationOutput[60]), .ZN(
        SubCellInst_LFInst_15_LFInst_0_n12) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_1_U4 ( .A1(
        SubCellInst_LFInst_15_LFInst_1_n9), .A2(
        SubCellInst_LFInst_15_LFInst_1_n8), .ZN(SboxOut[61]) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_1_U3 ( .A1(PermutationOutput[60]), 
        .A2(PermutationOutput[62]), .ZN(SubCellInst_LFInst_15_LFInst_1_n8) );
  OR2_X1 SubCellInst_LFInst_15_LFInst_1_U2 ( .A1(PermutationOutput[63]), .A2(
        SubCellInst_LFInst_15_LFInst_1_n7), .ZN(
        SubCellInst_LFInst_15_LFInst_1_n9) );
  NOR2_X1 SubCellInst_LFInst_15_LFInst_1_U1 ( .A1(PermutationOutput[60]), .A2(
        PermutationOutput[62]), .ZN(SubCellInst_LFInst_15_LFInst_1_n7) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_2_U6 ( .A1(
        SubCellInst_LFInst_15_LFInst_2_n18), .A2(
        SubCellInst_LFInst_15_LFInst_2_n17), .ZN(SboxOut[62]) );
  OR2_X1 SubCellInst_LFInst_15_LFInst_2_U5 ( .A1(PermutationOutput[60]), .A2(
        PermutationOutput[63]), .ZN(SubCellInst_LFInst_15_LFInst_2_n17) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_2_U4 ( .A1(PermutationOutput[61]), 
        .A2(SubCellInst_LFInst_15_LFInst_2_n16), .ZN(
        SubCellInst_LFInst_15_LFInst_2_n18) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_2_U3 ( .A1(
        SubCellInst_LFInst_15_LFInst_2_n15), .A2(
        SubCellInst_LFInst_15_LFInst_2_n14), .ZN(
        SubCellInst_LFInst_15_LFInst_2_n16) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_2_U2 ( .A1(PermutationOutput[60]), 
        .A2(PermutationOutput[63]), .ZN(SubCellInst_LFInst_15_LFInst_2_n14) );
  INV_X1 SubCellInst_LFInst_15_LFInst_2_U1 ( .A(PermutationOutput[62]), .ZN(
        SubCellInst_LFInst_15_LFInst_2_n15) );
  OR2_X1 SubCellInst_LFInst_15_LFInst_3_U4 ( .A1(
        SubCellInst_LFInst_15_LFInst_3_n9), .A2(
        SubCellInst_LFInst_15_LFInst_3_n8), .ZN(SboxOut[63]) );
  NOR2_X1 SubCellInst_LFInst_15_LFInst_3_U3 ( .A1(PermutationOutput[61]), .A2(
        PermutationOutput[62]), .ZN(SubCellInst_LFInst_15_LFInst_3_n8) );
  NOR2_X1 SubCellInst_LFInst_15_LFInst_3_U2 ( .A1(PermutationOutput[63]), .A2(
        SubCellInst_LFInst_15_LFInst_3_n7), .ZN(
        SubCellInst_LFInst_15_LFInst_3_n9) );
  AND2_X1 SubCellInst_LFInst_15_LFInst_3_U1 ( .A1(PermutationOutput[61]), .A2(
        PermutationOutput[60]), .ZN(SubCellInst_LFInst_15_LFInst_3_n7) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_0_U2 ( .A(MCInst2_XOR_r0_Inst_0_n5), .B(
        MCOutput2[16]), .ZN(MCOutput2[48]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_0_U1 ( .A(MCOutput2[0]), .B(SboxOut[48]), .ZN(
        MCInst2_XOR_r0_Inst_0_n5) );
  XOR2_X1 MCInst2_XOR_r1_Inst_0_U1 ( .A(SboxOut[32]), .B(MCOutput2[0]), .Z(
        MCOutput2[32]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_1_U2 ( .A(MCInst2_XOR_r0_Inst_1_n5), .B(
        MCOutput2[17]), .ZN(MCOutput2[49]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_1_U1 ( .A(MCOutput2[1]), .B(SboxOut[49]), .ZN(
        MCInst2_XOR_r0_Inst_1_n5) );
  XOR2_X1 MCInst2_XOR_r1_Inst_1_U1 ( .A(SboxOut[33]), .B(MCOutput2[1]), .Z(
        MCOutput2[33]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_2_U2 ( .A(MCInst2_XOR_r0_Inst_2_n5), .B(
        MCOutput2[18]), .ZN(MCOutput2[50]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_2_U1 ( .A(MCOutput2[2]), .B(SboxOut[50]), .ZN(
        MCInst2_XOR_r0_Inst_2_n5) );
  XOR2_X1 MCInst2_XOR_r1_Inst_2_U1 ( .A(SboxOut[34]), .B(MCOutput2[2]), .Z(
        MCOutput2[34]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_3_U2 ( .A(MCInst2_XOR_r0_Inst_3_n5), .B(
        MCOutput2[19]), .ZN(MCOutput2[51]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_3_U1 ( .A(MCOutput2[3]), .B(SboxOut[51]), .ZN(
        MCInst2_XOR_r0_Inst_3_n5) );
  XOR2_X1 MCInst2_XOR_r1_Inst_3_U1 ( .A(SboxOut[35]), .B(MCOutput2[3]), .Z(
        MCOutput2[35]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_4_U2 ( .A(MCInst2_XOR_r0_Inst_4_n5), .B(
        MCOutput2[20]), .ZN(MCOutput2[52]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_4_U1 ( .A(MCOutput2[4]), .B(SboxOut[52]), .ZN(
        MCInst2_XOR_r0_Inst_4_n5) );
  XOR2_X1 MCInst2_XOR_r1_Inst_4_U1 ( .A(SboxOut[36]), .B(MCOutput2[4]), .Z(
        MCOutput2[36]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_5_U2 ( .A(MCInst2_XOR_r0_Inst_5_n5), .B(
        MCOutput2[21]), .ZN(MCOutput2[53]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_5_U1 ( .A(MCOutput2[5]), .B(SboxOut[53]), .ZN(
        MCInst2_XOR_r0_Inst_5_n5) );
  XOR2_X1 MCInst2_XOR_r1_Inst_5_U1 ( .A(SboxOut[37]), .B(MCOutput2[5]), .Z(
        MCOutput2[37]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_6_U2 ( .A(MCInst2_XOR_r0_Inst_6_n5), .B(
        MCOutput2[22]), .ZN(MCOutput2[54]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_6_U1 ( .A(MCOutput2[6]), .B(SboxOut[54]), .ZN(
        MCInst2_XOR_r0_Inst_6_n5) );
  XOR2_X1 MCInst2_XOR_r1_Inst_6_U1 ( .A(SboxOut[38]), .B(MCOutput2[6]), .Z(
        MCOutput2[38]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_7_U2 ( .A(MCInst2_XOR_r0_Inst_7_n5), .B(
        MCOutput2[23]), .ZN(MCOutput2[55]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_7_U1 ( .A(MCOutput2[7]), .B(SboxOut[55]), .ZN(
        MCInst2_XOR_r0_Inst_7_n5) );
  XOR2_X1 MCInst2_XOR_r1_Inst_7_U1 ( .A(SboxOut[39]), .B(MCOutput2[7]), .Z(
        MCOutput2[39]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_8_U2 ( .A(MCInst2_XOR_r0_Inst_8_n5), .B(
        MCOutput2[24]), .ZN(MCOutput2[56]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_8_U1 ( .A(MCOutput2[8]), .B(SboxOut[56]), .ZN(
        MCInst2_XOR_r0_Inst_8_n5) );
  XOR2_X1 MCInst2_XOR_r1_Inst_8_U1 ( .A(SboxOut[40]), .B(MCOutput2[8]), .Z(
        MCOutput2[40]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_9_U2 ( .A(MCInst2_XOR_r0_Inst_9_n5), .B(
        MCOutput2[25]), .ZN(MCOutput2[57]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_9_U1 ( .A(MCOutput2[9]), .B(SboxOut[57]), .ZN(
        MCInst2_XOR_r0_Inst_9_n5) );
  XOR2_X1 MCInst2_XOR_r1_Inst_9_U1 ( .A(SboxOut[41]), .B(MCOutput2[9]), .Z(
        MCOutput2[41]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_10_U2 ( .A(MCInst2_XOR_r0_Inst_10_n5), .B(
        MCOutput2[26]), .ZN(MCOutput2[58]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_10_U1 ( .A(MCOutput2[10]), .B(SboxOut[58]), 
        .ZN(MCInst2_XOR_r0_Inst_10_n5) );
  XOR2_X1 MCInst2_XOR_r1_Inst_10_U1 ( .A(SboxOut[42]), .B(MCOutput2[10]), .Z(
        MCOutput2[42]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_11_U2 ( .A(MCInst2_XOR_r0_Inst_11_n5), .B(
        MCOutput2[27]), .ZN(MCOutput2[59]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_11_U1 ( .A(MCOutput2[11]), .B(SboxOut[59]), 
        .ZN(MCInst2_XOR_r0_Inst_11_n5) );
  XOR2_X1 MCInst2_XOR_r1_Inst_11_U1 ( .A(SboxOut[43]), .B(MCOutput2[11]), .Z(
        MCOutput2[43]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_12_U2 ( .A(MCInst2_XOR_r0_Inst_12_n5), .B(
        MCOutput2[28]), .ZN(MCOutput2[60]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_12_U1 ( .A(MCOutput2[12]), .B(SboxOut[60]), 
        .ZN(MCInst2_XOR_r0_Inst_12_n5) );
  XOR2_X1 MCInst2_XOR_r1_Inst_12_U1 ( .A(SboxOut[44]), .B(MCOutput2[12]), .Z(
        MCOutput2[44]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_13_U2 ( .A(MCInst2_XOR_r0_Inst_13_n5), .B(
        MCOutput2[29]), .ZN(MCOutput2[61]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_13_U1 ( .A(MCOutput2[13]), .B(SboxOut[61]), 
        .ZN(MCInst2_XOR_r0_Inst_13_n5) );
  XOR2_X1 MCInst2_XOR_r1_Inst_13_U1 ( .A(SboxOut[45]), .B(MCOutput2[13]), .Z(
        MCOutput2[45]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_14_U2 ( .A(MCInst2_XOR_r0_Inst_14_n5), .B(
        MCOutput2[30]), .ZN(MCOutput2[62]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_14_U1 ( .A(MCOutput2[14]), .B(SboxOut[62]), 
        .ZN(MCInst2_XOR_r0_Inst_14_n5) );
  XOR2_X1 MCInst2_XOR_r1_Inst_14_U1 ( .A(SboxOut[46]), .B(MCOutput2[14]), .Z(
        MCOutput2[46]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_15_U2 ( .A(MCInst2_XOR_r0_Inst_15_n5), .B(
        MCOutput2[31]), .ZN(MCOutput2[63]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_15_U1 ( .A(MCOutput2[15]), .B(SboxOut[63]), 
        .ZN(MCInst2_XOR_r0_Inst_15_n5) );
  XOR2_X1 MCInst2_XOR_r1_Inst_15_U1 ( .A(SboxOut[47]), .B(MCOutput2[15]), .Z(
        MCOutput2[47]) );
  XOR2_X1 AddKeyXOR12_XORInst_0_0_U1 ( .A(MCOutput2[48]), .B(Key[48]), .Z(
        AddRoundKeyOutput2[48]) );
  XOR2_X1 AddKeyXOR12_XORInst_0_1_U1 ( .A(MCOutput2[49]), .B(Key[49]), .Z(
        AddRoundKeyOutput2[49]) );
  XOR2_X1 AddKeyXOR12_XORInst_0_2_U1 ( .A(MCOutput2[50]), .B(Key[50]), .Z(
        AddRoundKeyOutput2[50]) );
  XOR2_X1 AddKeyXOR12_XORInst_0_3_U1 ( .A(MCOutput2[51]), .B(Key[51]), .Z(
        AddRoundKeyOutput2[51]) );
  XOR2_X1 AddKeyXOR12_XORInst_1_0_U1 ( .A(MCOutput2[52]), .B(Key[52]), .Z(
        AddRoundKeyOutput2[52]) );
  XOR2_X1 AddKeyXOR12_XORInst_1_1_U1 ( .A(MCOutput2[53]), .B(Key[53]), .Z(
        AddRoundKeyOutput2[53]) );
  XOR2_X1 AddKeyXOR12_XORInst_1_2_U1 ( .A(MCOutput2[54]), .B(Key[54]), .Z(
        AddRoundKeyOutput2[54]) );
  XOR2_X1 AddKeyXOR12_XORInst_1_3_U1 ( .A(MCOutput2[55]), .B(Key[55]), .Z(
        AddRoundKeyOutput2[55]) );
  XOR2_X1 AddKeyXOR12_XORInst_2_0_U1 ( .A(MCOutput2[56]), .B(Key[56]), .Z(
        AddRoundKeyOutput2[56]) );
  XOR2_X1 AddKeyXOR12_XORInst_2_1_U1 ( .A(MCOutput2[57]), .B(Key[57]), .Z(
        AddRoundKeyOutput2[57]) );
  XOR2_X1 AddKeyXOR12_XORInst_2_2_U1 ( .A(MCOutput2[58]), .B(Key[58]), .Z(
        AddRoundKeyOutput2[58]) );
  XOR2_X1 AddKeyXOR12_XORInst_2_3_U1 ( .A(MCOutput2[59]), .B(Key[59]), .Z(
        AddRoundKeyOutput2[59]) );
  XOR2_X1 AddKeyXOR12_XORInst_3_0_U1 ( .A(MCOutput2[60]), .B(Key[60]), .Z(
        AddRoundKeyOutput2[60]) );
  XOR2_X1 AddKeyXOR12_XORInst_3_1_U1 ( .A(MCOutput2[61]), .B(Key[61]), .Z(
        AddRoundKeyOutput2[61]) );
  XOR2_X1 AddKeyXOR12_XORInst_3_2_U1 ( .A(MCOutput2[62]), .B(Key[62]), .Z(
        AddRoundKeyOutput2[62]) );
  XOR2_X1 AddKeyXOR12_XORInst_3_3_U1 ( .A(MCOutput2[63]), .B(Key[63]), .Z(
        AddRoundKeyOutput2[63]) );
  XOR2_X1 AddKeyConstXOR2_XORInst_0_0_U1 ( .A(MCOutput2[40]), .B(Key[40]), .Z(
        AddRoundKeyOutput2[40]) );
  XOR2_X1 AddKeyConstXOR2_XORInst_0_1_U1 ( .A(MCOutput2[41]), .B(Key[41]), .Z(
        AddRoundKeyOutput2[41]) );
  XOR2_X1 AddKeyConstXOR2_XORInst_0_2_U1 ( .A(MCOutput2[42]), .B(Key[42]), .Z(
        AddRoundKeyOutput2[42]) );
  XOR2_X1 AddKeyConstXOR2_XORInst_0_3_U1 ( .A(MCOutput2[43]), .B(Key[43]), .Z(
        AddRoundKeyOutput2[43]) );
  XOR2_X1 AddKeyConstXOR2_XORInst_1_0_U1 ( .A(MCOutput2[44]), .B(Key[44]), .Z(
        AddRoundKeyOutput2[44]) );
  XOR2_X1 AddKeyConstXOR2_XORInst_1_1_U1 ( .A(MCOutput2[45]), .B(Key[45]), .Z(
        AddRoundKeyOutput2[45]) );
  XOR2_X1 AddKeyConstXOR2_XORInst_1_2_U1 ( .A(MCOutput2[46]), .B(Key[46]), .Z(
        AddRoundKeyOutput2[46]) );
  XOR2_X1 AddKeyConstXOR2_XORInst_1_3_U1 ( .A(MCOutput2[47]), .B(Key[47]), .Z(
        AddRoundKeyOutput2[47]) );
  XOR2_X1 AddKeyXOR22_XORInst_0_0_U1 ( .A(MCOutput2[0]), .B(Key[0]), .Z(
        AddRoundKeyOutput2[0]) );
  XOR2_X1 AddKeyXOR22_XORInst_0_1_U1 ( .A(MCOutput2[1]), .B(Key[1]), .Z(
        AddRoundKeyOutput2[1]) );
  XOR2_X1 AddKeyXOR22_XORInst_0_2_U1 ( .A(MCOutput2[2]), .B(Key[2]), .Z(
        AddRoundKeyOutput2[2]) );
  XOR2_X1 AddKeyXOR22_XORInst_0_3_U1 ( .A(MCOutput2[3]), .B(Key[3]), .Z(
        AddRoundKeyOutput2[3]) );
  XOR2_X1 AddKeyXOR22_XORInst_1_0_U1 ( .A(MCOutput2[4]), .B(Key[4]), .Z(
        AddRoundKeyOutput2[4]) );
  XOR2_X1 AddKeyXOR22_XORInst_1_1_U1 ( .A(MCOutput2[5]), .B(Key[5]), .Z(
        AddRoundKeyOutput2[5]) );
  XOR2_X1 AddKeyXOR22_XORInst_1_2_U1 ( .A(MCOutput2[6]), .B(Key[6]), .Z(
        AddRoundKeyOutput2[6]) );
  XOR2_X1 AddKeyXOR22_XORInst_1_3_U1 ( .A(MCOutput2[7]), .B(Key[7]), .Z(
        AddRoundKeyOutput2[7]) );
  XOR2_X1 AddKeyXOR22_XORInst_2_0_U1 ( .A(MCOutput2[8]), .B(Key[8]), .Z(
        AddRoundKeyOutput2[8]) );
  XOR2_X1 AddKeyXOR22_XORInst_2_1_U1 ( .A(MCOutput2[9]), .B(Key[9]), .Z(
        AddRoundKeyOutput2[9]) );
  XOR2_X1 AddKeyXOR22_XORInst_2_2_U1 ( .A(MCOutput2[10]), .B(Key[10]), .Z(
        AddRoundKeyOutput2[10]) );
  XOR2_X1 AddKeyXOR22_XORInst_2_3_U1 ( .A(MCOutput2[11]), .B(Key[11]), .Z(
        AddRoundKeyOutput2[11]) );
  XOR2_X1 AddKeyXOR22_XORInst_3_0_U1 ( .A(MCOutput2[12]), .B(Key[12]), .Z(
        AddRoundKeyOutput2[12]) );
  XOR2_X1 AddKeyXOR22_XORInst_3_1_U1 ( .A(MCOutput2[13]), .B(Key[13]), .Z(
        AddRoundKeyOutput2[13]) );
  XOR2_X1 AddKeyXOR22_XORInst_3_2_U1 ( .A(MCOutput2[14]), .B(Key[14]), .Z(
        AddRoundKeyOutput2[14]) );
  XOR2_X1 AddKeyXOR22_XORInst_3_3_U1 ( .A(MCOutput2[15]), .B(Key[15]), .Z(
        AddRoundKeyOutput2[15]) );
  XOR2_X1 AddKeyXOR22_XORInst_4_0_U1 ( .A(MCOutput2[16]), .B(Key[16]), .Z(
        AddRoundKeyOutput2[16]) );
  XOR2_X1 AddKeyXOR22_XORInst_4_1_U1 ( .A(MCOutput2[17]), .B(Key[17]), .Z(
        AddRoundKeyOutput2[17]) );
  XOR2_X1 AddKeyXOR22_XORInst_4_2_U1 ( .A(MCOutput2[18]), .B(Key[18]), .Z(
        AddRoundKeyOutput2[18]) );
  XOR2_X1 AddKeyXOR22_XORInst_4_3_U1 ( .A(MCOutput2[19]), .B(Key[19]), .Z(
        AddRoundKeyOutput2[19]) );
  XOR2_X1 AddKeyXOR22_XORInst_5_0_U1 ( .A(MCOutput2[20]), .B(Key[20]), .Z(
        AddRoundKeyOutput2[20]) );
  XOR2_X1 AddKeyXOR22_XORInst_5_1_U1 ( .A(MCOutput2[21]), .B(Key[21]), .Z(
        AddRoundKeyOutput2[21]) );
  XOR2_X1 AddKeyXOR22_XORInst_5_2_U1 ( .A(MCOutput2[22]), .B(Key[22]), .Z(
        AddRoundKeyOutput2[22]) );
  XOR2_X1 AddKeyXOR22_XORInst_5_3_U1 ( .A(MCOutput2[23]), .B(Key[23]), .Z(
        AddRoundKeyOutput2[23]) );
  XOR2_X1 AddKeyXOR22_XORInst_6_0_U1 ( .A(MCOutput2[24]), .B(Key[24]), .Z(
        AddRoundKeyOutput2[24]) );
  XOR2_X1 AddKeyXOR22_XORInst_6_1_U1 ( .A(MCOutput2[25]), .B(Key[25]), .Z(
        AddRoundKeyOutput2[25]) );
  XOR2_X1 AddKeyXOR22_XORInst_6_2_U1 ( .A(MCOutput2[26]), .B(Key[26]), .Z(
        AddRoundKeyOutput2[26]) );
  XOR2_X1 AddKeyXOR22_XORInst_6_3_U1 ( .A(MCOutput2[27]), .B(Key[27]), .Z(
        AddRoundKeyOutput2[27]) );
  XOR2_X1 AddKeyXOR22_XORInst_7_0_U1 ( .A(MCOutput2[28]), .B(Key[28]), .Z(
        AddRoundKeyOutput2[28]) );
  XOR2_X1 AddKeyXOR22_XORInst_7_1_U1 ( .A(MCOutput2[29]), .B(Key[29]), .Z(
        AddRoundKeyOutput2[29]) );
  XOR2_X1 AddKeyXOR22_XORInst_7_2_U1 ( .A(MCOutput2[30]), .B(Key[30]), .Z(
        AddRoundKeyOutput2[30]) );
  XOR2_X1 AddKeyXOR22_XORInst_7_3_U1 ( .A(MCOutput2[31]), .B(Key[31]), .Z(
        AddRoundKeyOutput2[31]) );
  XOR2_X1 AddKeyXOR22_XORInst_8_0_U1 ( .A(MCOutput2[32]), .B(Key[32]), .Z(
        AddRoundKeyOutput2[32]) );
  XOR2_X1 AddKeyXOR22_XORInst_8_1_U1 ( .A(MCOutput2[33]), .B(Key[33]), .Z(
        AddRoundKeyOutput2[33]) );
  XOR2_X1 AddKeyXOR22_XORInst_8_2_U1 ( .A(MCOutput2[34]), .B(Key[34]), .Z(
        AddRoundKeyOutput2[34]) );
  XOR2_X1 AddKeyXOR22_XORInst_8_3_U1 ( .A(MCOutput2[35]), .B(Key[35]), .Z(
        AddRoundKeyOutput2[35]) );
  XOR2_X1 AddKeyXOR22_XORInst_9_0_U1 ( .A(MCOutput2[36]), .B(Key[36]), .Z(
        AddRoundKeyOutput2[36]) );
  XOR2_X1 AddKeyXOR22_XORInst_9_1_U1 ( .A(MCOutput2[37]), .B(Key[37]), .Z(
        AddRoundKeyOutput2[37]) );
  XOR2_X1 AddKeyXOR22_XORInst_9_2_U1 ( .A(MCOutput2[38]), .B(Key[38]), .Z(
        AddRoundKeyOutput2[38]) );
  XOR2_X1 AddKeyXOR22_XORInst_9_3_U1 ( .A(MCOutput2[39]), .B(Key[39]), .Z(
        AddRoundKeyOutput2[39]) );
  DFF_X1 StateReg2_s_current_state_reg_0_ ( .D(AddRoundKeyOutput2[0]), .CK(clk), .Q(PermutationOutput2[60]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_1_ ( .D(AddRoundKeyOutput2[1]), .CK(clk), .Q(PermutationOutput2[61]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_2_ ( .D(AddRoundKeyOutput2[2]), .CK(clk), .Q(PermutationOutput2[62]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_3_ ( .D(AddRoundKeyOutput2[3]), .CK(clk), .Q(PermutationOutput2[63]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_4_ ( .D(AddRoundKeyOutput2[4]), .CK(clk), .Q(PermutationOutput2[48]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_5_ ( .D(AddRoundKeyOutput2[5]), .CK(clk), .Q(PermutationOutput2[49]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_6_ ( .D(AddRoundKeyOutput2[6]), .CK(clk), .Q(PermutationOutput2[50]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_7_ ( .D(AddRoundKeyOutput2[7]), .CK(clk), .Q(PermutationOutput2[51]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_8_ ( .D(AddRoundKeyOutput2[8]), .CK(clk), .Q(PermutationOutput2[52]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_9_ ( .D(AddRoundKeyOutput2[9]), .CK(clk), .Q(PermutationOutput2[53]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_10_ ( .D(AddRoundKeyOutput2[10]), .CK(
        clk), .Q(PermutationOutput2[54]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_11_ ( .D(AddRoundKeyOutput2[11]), .CK(
        clk), .Q(PermutationOutput2[55]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_12_ ( .D(AddRoundKeyOutput2[12]), .CK(
        clk), .Q(PermutationOutput2[56]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_13_ ( .D(AddRoundKeyOutput2[13]), .CK(
        clk), .Q(PermutationOutput2[57]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_14_ ( .D(AddRoundKeyOutput2[14]), .CK(
        clk), .Q(PermutationOutput2[58]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_15_ ( .D(AddRoundKeyOutput2[15]), .CK(
        clk), .Q(PermutationOutput2[59]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_16_ ( .D(AddRoundKeyOutput2[16]), .CK(
        clk), .Q(PermutationOutput2[32]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_17_ ( .D(AddRoundKeyOutput2[17]), .CK(
        clk), .Q(PermutationOutput2[33]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_18_ ( .D(AddRoundKeyOutput2[18]), .CK(
        clk), .Q(PermutationOutput2[34]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_19_ ( .D(AddRoundKeyOutput2[19]), .CK(
        clk), .Q(PermutationOutput2[35]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_20_ ( .D(AddRoundKeyOutput2[20]), .CK(
        clk), .Q(PermutationOutput2[44]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_21_ ( .D(AddRoundKeyOutput2[21]), .CK(
        clk), .Q(PermutationOutput2[45]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_22_ ( .D(AddRoundKeyOutput2[22]), .CK(
        clk), .Q(PermutationOutput2[46]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_23_ ( .D(AddRoundKeyOutput2[23]), .CK(
        clk), .Q(PermutationOutput2[47]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_24_ ( .D(AddRoundKeyOutput2[24]), .CK(
        clk), .Q(PermutationOutput2[40]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_25_ ( .D(AddRoundKeyOutput2[25]), .CK(
        clk), .Q(PermutationOutput2[41]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_26_ ( .D(AddRoundKeyOutput2[26]), .CK(
        clk), .Q(PermutationOutput2[42]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_27_ ( .D(AddRoundKeyOutput2[27]), .CK(
        clk), .Q(PermutationOutput2[43]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_28_ ( .D(AddRoundKeyOutput2[28]), .CK(
        clk), .Q(PermutationOutput2[36]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_29_ ( .D(AddRoundKeyOutput2[29]), .CK(
        clk), .Q(PermutationOutput2[37]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_30_ ( .D(AddRoundKeyOutput2[30]), .CK(
        clk), .Q(PermutationOutput2[38]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_31_ ( .D(AddRoundKeyOutput2[31]), .CK(
        clk), .Q(PermutationOutput2[39]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_32_ ( .D(AddRoundKeyOutput2[32]), .CK(
        clk), .Q(PermutationOutput2[16]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_33_ ( .D(AddRoundKeyOutput2[33]), .CK(
        clk), .Q(PermutationOutput2[17]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_34_ ( .D(AddRoundKeyOutput2[34]), .CK(
        clk), .Q(PermutationOutput2[18]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_35_ ( .D(AddRoundKeyOutput2[35]), .CK(
        clk), .Q(PermutationOutput2[19]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_36_ ( .D(AddRoundKeyOutput2[36]), .CK(
        clk), .Q(PermutationOutput2[28]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_37_ ( .D(AddRoundKeyOutput2[37]), .CK(
        clk), .Q(PermutationOutput2[29]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_38_ ( .D(AddRoundKeyOutput2[38]), .CK(
        clk), .Q(PermutationOutput2[30]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_39_ ( .D(AddRoundKeyOutput2[39]), .CK(
        clk), .Q(PermutationOutput2[31]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_40_ ( .D(AddRoundKeyOutput2[40]), .CK(
        clk), .Q(PermutationOutput2[24]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_41_ ( .D(AddRoundKeyOutput2[41]), .CK(
        clk), .Q(PermutationOutput2[25]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_42_ ( .D(AddRoundKeyOutput2[42]), .CK(
        clk), .Q(PermutationOutput2[26]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_43_ ( .D(AddRoundKeyOutput2[43]), .CK(
        clk), .Q(PermutationOutput2[27]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_44_ ( .D(AddRoundKeyOutput2[44]), .CK(
        clk), .Q(PermutationOutput2[20]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_45_ ( .D(AddRoundKeyOutput2[45]), .CK(
        clk), .Q(PermutationOutput2[21]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_46_ ( .D(AddRoundKeyOutput2[46]), .CK(
        clk), .Q(PermutationOutput2[22]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_47_ ( .D(AddRoundKeyOutput2[47]), .CK(
        clk), .Q(PermutationOutput2[23]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_48_ ( .D(AddRoundKeyOutput2[48]), .CK(
        clk), .Q(PermutationOutput2[4]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_49_ ( .D(AddRoundKeyOutput2[49]), .CK(
        clk), .Q(PermutationOutput2[5]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_50_ ( .D(AddRoundKeyOutput2[50]), .CK(
        clk), .Q(PermutationOutput2[6]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_51_ ( .D(AddRoundKeyOutput2[51]), .CK(
        clk), .Q(PermutationOutput2[7]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_52_ ( .D(AddRoundKeyOutput2[52]), .CK(
        clk), .Q(PermutationOutput2[8]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_53_ ( .D(AddRoundKeyOutput2[53]), .CK(
        clk), .Q(PermutationOutput2[9]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_54_ ( .D(AddRoundKeyOutput2[54]), .CK(
        clk), .Q(PermutationOutput2[10]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_55_ ( .D(AddRoundKeyOutput2[55]), .CK(
        clk), .Q(PermutationOutput2[11]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_56_ ( .D(AddRoundKeyOutput2[56]), .CK(
        clk), .Q(PermutationOutput2[12]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_57_ ( .D(AddRoundKeyOutput2[57]), .CK(
        clk), .Q(PermutationOutput2[13]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_58_ ( .D(AddRoundKeyOutput2[58]), .CK(
        clk), .Q(PermutationOutput2[14]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_59_ ( .D(AddRoundKeyOutput2[59]), .CK(
        clk), .Q(PermutationOutput2[15]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_60_ ( .D(AddRoundKeyOutput2[60]), .CK(
        clk), .Q(PermutationOutput2[0]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_61_ ( .D(AddRoundKeyOutput2[61]), .CK(
        clk), .Q(PermutationOutput2[1]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_62_ ( .D(AddRoundKeyOutput2[62]), .CK(
        clk), .Q(PermutationOutput2[2]), .QN() );
  DFF_X1 StateReg2_s_current_state_reg_63_ ( .D(AddRoundKeyOutput2[63]), .CK(
        clk), .Q(PermutationOutput2[3]), .QN() );
  NOR2_X1 SubCellInst2_LFInst_0_LFInst_0_U6 ( .A1(
        SubCellInst2_LFInst_0_LFInst_0_n15), .A2(
        SubCellInst2_LFInst_0_LFInst_0_n14), .ZN(Output[0]) );
  AND2_X1 SubCellInst2_LFInst_0_LFInst_0_U5 ( .A1(PermutationOutput2[3]), .A2(
        PermutationOutput2[2]), .ZN(SubCellInst2_LFInst_0_LFInst_0_n14) );
  NOR2_X1 SubCellInst2_LFInst_0_LFInst_0_U4 ( .A1(PermutationOutput2[1]), .A2(
        SubCellInst2_LFInst_0_LFInst_0_n13), .ZN(
        SubCellInst2_LFInst_0_LFInst_0_n15) );
  NOR2_X1 SubCellInst2_LFInst_0_LFInst_0_U3 ( .A1(
        SubCellInst2_LFInst_0_LFInst_0_n12), .A2(
        SubCellInst2_LFInst_0_LFInst_0_n11), .ZN(
        SubCellInst2_LFInst_0_LFInst_0_n13) );
  NOR2_X1 SubCellInst2_LFInst_0_LFInst_0_U2 ( .A1(PermutationOutput2[3]), .A2(
        PermutationOutput2[2]), .ZN(SubCellInst2_LFInst_0_LFInst_0_n11) );
  INV_X1 SubCellInst2_LFInst_0_LFInst_0_U1 ( .A(PermutationOutput2[0]), .ZN(
        SubCellInst2_LFInst_0_LFInst_0_n12) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_1_U4 ( .A1(
        SubCellInst2_LFInst_0_LFInst_1_n9), .A2(
        SubCellInst2_LFInst_0_LFInst_1_n8), .ZN(Output[1]) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_1_U3 ( .A1(PermutationOutput2[0]), 
        .A2(PermutationOutput2[2]), .ZN(SubCellInst2_LFInst_0_LFInst_1_n8) );
  OR2_X1 SubCellInst2_LFInst_0_LFInst_1_U2 ( .A1(PermutationOutput2[3]), .A2(
        SubCellInst2_LFInst_0_LFInst_1_n7), .ZN(
        SubCellInst2_LFInst_0_LFInst_1_n9) );
  NOR2_X1 SubCellInst2_LFInst_0_LFInst_1_U1 ( .A1(PermutationOutput2[0]), .A2(
        PermutationOutput2[2]), .ZN(SubCellInst2_LFInst_0_LFInst_1_n7) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_2_U6 ( .A1(
        SubCellInst2_LFInst_0_LFInst_2_n18), .A2(
        SubCellInst2_LFInst_0_LFInst_2_n17), .ZN(Output[2]) );
  OR2_X1 SubCellInst2_LFInst_0_LFInst_2_U5 ( .A1(PermutationOutput2[0]), .A2(
        PermutationOutput2[3]), .ZN(SubCellInst2_LFInst_0_LFInst_2_n17) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_2_U4 ( .A1(PermutationOutput2[1]), 
        .A2(SubCellInst2_LFInst_0_LFInst_2_n16), .ZN(
        SubCellInst2_LFInst_0_LFInst_2_n18) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_2_U3 ( .A1(
        SubCellInst2_LFInst_0_LFInst_2_n15), .A2(
        SubCellInst2_LFInst_0_LFInst_2_n14), .ZN(
        SubCellInst2_LFInst_0_LFInst_2_n16) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_2_U2 ( .A1(PermutationOutput2[0]), 
        .A2(PermutationOutput2[3]), .ZN(SubCellInst2_LFInst_0_LFInst_2_n14) );
  INV_X1 SubCellInst2_LFInst_0_LFInst_2_U1 ( .A(PermutationOutput2[2]), .ZN(
        SubCellInst2_LFInst_0_LFInst_2_n15) );
  OR2_X1 SubCellInst2_LFInst_0_LFInst_3_U4 ( .A1(
        SubCellInst2_LFInst_0_LFInst_3_n9), .A2(
        SubCellInst2_LFInst_0_LFInst_3_n8), .ZN(Output[3]) );
  NOR2_X1 SubCellInst2_LFInst_0_LFInst_3_U3 ( .A1(PermutationOutput2[1]), .A2(
        PermutationOutput2[2]), .ZN(SubCellInst2_LFInst_0_LFInst_3_n8) );
  NOR2_X1 SubCellInst2_LFInst_0_LFInst_3_U2 ( .A1(PermutationOutput2[3]), .A2(
        SubCellInst2_LFInst_0_LFInst_3_n7), .ZN(
        SubCellInst2_LFInst_0_LFInst_3_n9) );
  AND2_X1 SubCellInst2_LFInst_0_LFInst_3_U1 ( .A1(PermutationOutput2[1]), .A2(
        PermutationOutput2[0]), .ZN(SubCellInst2_LFInst_0_LFInst_3_n7) );
  NOR2_X1 SubCellInst2_LFInst_1_LFInst_0_U6 ( .A1(
        SubCellInst2_LFInst_1_LFInst_0_n15), .A2(
        SubCellInst2_LFInst_1_LFInst_0_n14), .ZN(Output[4]) );
  AND2_X1 SubCellInst2_LFInst_1_LFInst_0_U5 ( .A1(PermutationOutput2[7]), .A2(
        PermutationOutput2[6]), .ZN(SubCellInst2_LFInst_1_LFInst_0_n14) );
  NOR2_X1 SubCellInst2_LFInst_1_LFInst_0_U4 ( .A1(PermutationOutput2[5]), .A2(
        SubCellInst2_LFInst_1_LFInst_0_n13), .ZN(
        SubCellInst2_LFInst_1_LFInst_0_n15) );
  NOR2_X1 SubCellInst2_LFInst_1_LFInst_0_U3 ( .A1(
        SubCellInst2_LFInst_1_LFInst_0_n12), .A2(
        SubCellInst2_LFInst_1_LFInst_0_n11), .ZN(
        SubCellInst2_LFInst_1_LFInst_0_n13) );
  NOR2_X1 SubCellInst2_LFInst_1_LFInst_0_U2 ( .A1(PermutationOutput2[7]), .A2(
        PermutationOutput2[6]), .ZN(SubCellInst2_LFInst_1_LFInst_0_n11) );
  INV_X1 SubCellInst2_LFInst_1_LFInst_0_U1 ( .A(PermutationOutput2[4]), .ZN(
        SubCellInst2_LFInst_1_LFInst_0_n12) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_1_U4 ( .A1(
        SubCellInst2_LFInst_1_LFInst_1_n9), .A2(
        SubCellInst2_LFInst_1_LFInst_1_n8), .ZN(Output[5]) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_1_U3 ( .A1(PermutationOutput2[4]), 
        .A2(PermutationOutput2[6]), .ZN(SubCellInst2_LFInst_1_LFInst_1_n8) );
  OR2_X1 SubCellInst2_LFInst_1_LFInst_1_U2 ( .A1(PermutationOutput2[7]), .A2(
        SubCellInst2_LFInst_1_LFInst_1_n7), .ZN(
        SubCellInst2_LFInst_1_LFInst_1_n9) );
  NOR2_X1 SubCellInst2_LFInst_1_LFInst_1_U1 ( .A1(PermutationOutput2[4]), .A2(
        PermutationOutput2[6]), .ZN(SubCellInst2_LFInst_1_LFInst_1_n7) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_2_U6 ( .A1(
        SubCellInst2_LFInst_1_LFInst_2_n18), .A2(
        SubCellInst2_LFInst_1_LFInst_2_n17), .ZN(Output[6]) );
  OR2_X1 SubCellInst2_LFInst_1_LFInst_2_U5 ( .A1(PermutationOutput2[4]), .A2(
        PermutationOutput2[7]), .ZN(SubCellInst2_LFInst_1_LFInst_2_n17) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_2_U4 ( .A1(PermutationOutput2[5]), 
        .A2(SubCellInst2_LFInst_1_LFInst_2_n16), .ZN(
        SubCellInst2_LFInst_1_LFInst_2_n18) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_2_U3 ( .A1(
        SubCellInst2_LFInst_1_LFInst_2_n15), .A2(
        SubCellInst2_LFInst_1_LFInst_2_n14), .ZN(
        SubCellInst2_LFInst_1_LFInst_2_n16) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_2_U2 ( .A1(PermutationOutput2[4]), 
        .A2(PermutationOutput2[7]), .ZN(SubCellInst2_LFInst_1_LFInst_2_n14) );
  INV_X1 SubCellInst2_LFInst_1_LFInst_2_U1 ( .A(PermutationOutput2[6]), .ZN(
        SubCellInst2_LFInst_1_LFInst_2_n15) );
  OR2_X1 SubCellInst2_LFInst_1_LFInst_3_U4 ( .A1(
        SubCellInst2_LFInst_1_LFInst_3_n9), .A2(
        SubCellInst2_LFInst_1_LFInst_3_n8), .ZN(Output[7]) );
  NOR2_X1 SubCellInst2_LFInst_1_LFInst_3_U3 ( .A1(PermutationOutput2[5]), .A2(
        PermutationOutput2[6]), .ZN(SubCellInst2_LFInst_1_LFInst_3_n8) );
  NOR2_X1 SubCellInst2_LFInst_1_LFInst_3_U2 ( .A1(PermutationOutput2[7]), .A2(
        SubCellInst2_LFInst_1_LFInst_3_n7), .ZN(
        SubCellInst2_LFInst_1_LFInst_3_n9) );
  AND2_X1 SubCellInst2_LFInst_1_LFInst_3_U1 ( .A1(PermutationOutput2[5]), .A2(
        PermutationOutput2[4]), .ZN(SubCellInst2_LFInst_1_LFInst_3_n7) );
  NOR2_X1 SubCellInst2_LFInst_2_LFInst_0_U6 ( .A1(
        SubCellInst2_LFInst_2_LFInst_0_n15), .A2(
        SubCellInst2_LFInst_2_LFInst_0_n14), .ZN(Output[8]) );
  AND2_X1 SubCellInst2_LFInst_2_LFInst_0_U5 ( .A1(PermutationOutput2[11]), 
        .A2(PermutationOutput2[10]), .ZN(SubCellInst2_LFInst_2_LFInst_0_n14)
         );
  NOR2_X1 SubCellInst2_LFInst_2_LFInst_0_U4 ( .A1(PermutationOutput2[9]), .A2(
        SubCellInst2_LFInst_2_LFInst_0_n13), .ZN(
        SubCellInst2_LFInst_2_LFInst_0_n15) );
  NOR2_X1 SubCellInst2_LFInst_2_LFInst_0_U3 ( .A1(
        SubCellInst2_LFInst_2_LFInst_0_n12), .A2(
        SubCellInst2_LFInst_2_LFInst_0_n11), .ZN(
        SubCellInst2_LFInst_2_LFInst_0_n13) );
  NOR2_X1 SubCellInst2_LFInst_2_LFInst_0_U2 ( .A1(PermutationOutput2[11]), 
        .A2(PermutationOutput2[10]), .ZN(SubCellInst2_LFInst_2_LFInst_0_n11)
         );
  INV_X1 SubCellInst2_LFInst_2_LFInst_0_U1 ( .A(PermutationOutput2[8]), .ZN(
        SubCellInst2_LFInst_2_LFInst_0_n12) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_1_U4 ( .A1(
        SubCellInst2_LFInst_2_LFInst_1_n9), .A2(
        SubCellInst2_LFInst_2_LFInst_1_n8), .ZN(Output[9]) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_1_U3 ( .A1(PermutationOutput2[8]), 
        .A2(PermutationOutput2[10]), .ZN(SubCellInst2_LFInst_2_LFInst_1_n8) );
  OR2_X1 SubCellInst2_LFInst_2_LFInst_1_U2 ( .A1(PermutationOutput2[11]), .A2(
        SubCellInst2_LFInst_2_LFInst_1_n7), .ZN(
        SubCellInst2_LFInst_2_LFInst_1_n9) );
  NOR2_X1 SubCellInst2_LFInst_2_LFInst_1_U1 ( .A1(PermutationOutput2[8]), .A2(
        PermutationOutput2[10]), .ZN(SubCellInst2_LFInst_2_LFInst_1_n7) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_2_U6 ( .A1(
        SubCellInst2_LFInst_2_LFInst_2_n18), .A2(
        SubCellInst2_LFInst_2_LFInst_2_n17), .ZN(Output[10]) );
  OR2_X1 SubCellInst2_LFInst_2_LFInst_2_U5 ( .A1(PermutationOutput2[8]), .A2(
        PermutationOutput2[11]), .ZN(SubCellInst2_LFInst_2_LFInst_2_n17) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_2_U4 ( .A1(PermutationOutput2[9]), 
        .A2(SubCellInst2_LFInst_2_LFInst_2_n16), .ZN(
        SubCellInst2_LFInst_2_LFInst_2_n18) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_2_U3 ( .A1(
        SubCellInst2_LFInst_2_LFInst_2_n15), .A2(
        SubCellInst2_LFInst_2_LFInst_2_n14), .ZN(
        SubCellInst2_LFInst_2_LFInst_2_n16) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_2_U2 ( .A1(PermutationOutput2[8]), 
        .A2(PermutationOutput2[11]), .ZN(SubCellInst2_LFInst_2_LFInst_2_n14)
         );
  INV_X1 SubCellInst2_LFInst_2_LFInst_2_U1 ( .A(PermutationOutput2[10]), .ZN(
        SubCellInst2_LFInst_2_LFInst_2_n15) );
  OR2_X1 SubCellInst2_LFInst_2_LFInst_3_U4 ( .A1(
        SubCellInst2_LFInst_2_LFInst_3_n9), .A2(
        SubCellInst2_LFInst_2_LFInst_3_n8), .ZN(Output[11]) );
  NOR2_X1 SubCellInst2_LFInst_2_LFInst_3_U3 ( .A1(PermutationOutput2[9]), .A2(
        PermutationOutput2[10]), .ZN(SubCellInst2_LFInst_2_LFInst_3_n8) );
  NOR2_X1 SubCellInst2_LFInst_2_LFInst_3_U2 ( .A1(PermutationOutput2[11]), 
        .A2(SubCellInst2_LFInst_2_LFInst_3_n7), .ZN(
        SubCellInst2_LFInst_2_LFInst_3_n9) );
  AND2_X1 SubCellInst2_LFInst_2_LFInst_3_U1 ( .A1(PermutationOutput2[9]), .A2(
        PermutationOutput2[8]), .ZN(SubCellInst2_LFInst_2_LFInst_3_n7) );
  NOR2_X1 SubCellInst2_LFInst_3_LFInst_0_U6 ( .A1(
        SubCellInst2_LFInst_3_LFInst_0_n15), .A2(
        SubCellInst2_LFInst_3_LFInst_0_n14), .ZN(Output[12]) );
  AND2_X1 SubCellInst2_LFInst_3_LFInst_0_U5 ( .A1(PermutationOutput2[15]), 
        .A2(PermutationOutput2[14]), .ZN(SubCellInst2_LFInst_3_LFInst_0_n14)
         );
  NOR2_X1 SubCellInst2_LFInst_3_LFInst_0_U4 ( .A1(PermutationOutput2[13]), 
        .A2(SubCellInst2_LFInst_3_LFInst_0_n13), .ZN(
        SubCellInst2_LFInst_3_LFInst_0_n15) );
  NOR2_X1 SubCellInst2_LFInst_3_LFInst_0_U3 ( .A1(
        SubCellInst2_LFInst_3_LFInst_0_n12), .A2(
        SubCellInst2_LFInst_3_LFInst_0_n11), .ZN(
        SubCellInst2_LFInst_3_LFInst_0_n13) );
  NOR2_X1 SubCellInst2_LFInst_3_LFInst_0_U2 ( .A1(PermutationOutput2[15]), 
        .A2(PermutationOutput2[14]), .ZN(SubCellInst2_LFInst_3_LFInst_0_n11)
         );
  INV_X1 SubCellInst2_LFInst_3_LFInst_0_U1 ( .A(PermutationOutput2[12]), .ZN(
        SubCellInst2_LFInst_3_LFInst_0_n12) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_1_U4 ( .A1(
        SubCellInst2_LFInst_3_LFInst_1_n9), .A2(
        SubCellInst2_LFInst_3_LFInst_1_n8), .ZN(Output[13]) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_1_U3 ( .A1(PermutationOutput2[12]), 
        .A2(PermutationOutput2[14]), .ZN(SubCellInst2_LFInst_3_LFInst_1_n8) );
  OR2_X1 SubCellInst2_LFInst_3_LFInst_1_U2 ( .A1(PermutationOutput2[15]), .A2(
        SubCellInst2_LFInst_3_LFInst_1_n7), .ZN(
        SubCellInst2_LFInst_3_LFInst_1_n9) );
  NOR2_X1 SubCellInst2_LFInst_3_LFInst_1_U1 ( .A1(PermutationOutput2[12]), 
        .A2(PermutationOutput2[14]), .ZN(SubCellInst2_LFInst_3_LFInst_1_n7) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_2_U6 ( .A1(
        SubCellInst2_LFInst_3_LFInst_2_n18), .A2(
        SubCellInst2_LFInst_3_LFInst_2_n17), .ZN(Output[14]) );
  OR2_X1 SubCellInst2_LFInst_3_LFInst_2_U5 ( .A1(PermutationOutput2[12]), .A2(
        PermutationOutput2[15]), .ZN(SubCellInst2_LFInst_3_LFInst_2_n17) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_2_U4 ( .A1(PermutationOutput2[13]), 
        .A2(SubCellInst2_LFInst_3_LFInst_2_n16), .ZN(
        SubCellInst2_LFInst_3_LFInst_2_n18) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_2_U3 ( .A1(
        SubCellInst2_LFInst_3_LFInst_2_n15), .A2(
        SubCellInst2_LFInst_3_LFInst_2_n14), .ZN(
        SubCellInst2_LFInst_3_LFInst_2_n16) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_2_U2 ( .A1(PermutationOutput2[12]), 
        .A2(PermutationOutput2[15]), .ZN(SubCellInst2_LFInst_3_LFInst_2_n14)
         );
  INV_X1 SubCellInst2_LFInst_3_LFInst_2_U1 ( .A(PermutationOutput2[14]), .ZN(
        SubCellInst2_LFInst_3_LFInst_2_n15) );
  OR2_X1 SubCellInst2_LFInst_3_LFInst_3_U4 ( .A1(
        SubCellInst2_LFInst_3_LFInst_3_n9), .A2(
        SubCellInst2_LFInst_3_LFInst_3_n8), .ZN(Output[15]) );
  NOR2_X1 SubCellInst2_LFInst_3_LFInst_3_U3 ( .A1(PermutationOutput2[13]), 
        .A2(PermutationOutput2[14]), .ZN(SubCellInst2_LFInst_3_LFInst_3_n8) );
  NOR2_X1 SubCellInst2_LFInst_3_LFInst_3_U2 ( .A1(PermutationOutput2[15]), 
        .A2(SubCellInst2_LFInst_3_LFInst_3_n7), .ZN(
        SubCellInst2_LFInst_3_LFInst_3_n9) );
  AND2_X1 SubCellInst2_LFInst_3_LFInst_3_U1 ( .A1(PermutationOutput2[13]), 
        .A2(PermutationOutput2[12]), .ZN(SubCellInst2_LFInst_3_LFInst_3_n7) );
  NOR2_X1 SubCellInst2_LFInst_4_LFInst_0_U6 ( .A1(
        SubCellInst2_LFInst_4_LFInst_0_n15), .A2(
        SubCellInst2_LFInst_4_LFInst_0_n14), .ZN(Output[16]) );
  AND2_X1 SubCellInst2_LFInst_4_LFInst_0_U5 ( .A1(PermutationOutput2[19]), 
        .A2(PermutationOutput2[18]), .ZN(SubCellInst2_LFInst_4_LFInst_0_n14)
         );
  NOR2_X1 SubCellInst2_LFInst_4_LFInst_0_U4 ( .A1(PermutationOutput2[17]), 
        .A2(SubCellInst2_LFInst_4_LFInst_0_n13), .ZN(
        SubCellInst2_LFInst_4_LFInst_0_n15) );
  NOR2_X1 SubCellInst2_LFInst_4_LFInst_0_U3 ( .A1(
        SubCellInst2_LFInst_4_LFInst_0_n12), .A2(
        SubCellInst2_LFInst_4_LFInst_0_n11), .ZN(
        SubCellInst2_LFInst_4_LFInst_0_n13) );
  NOR2_X1 SubCellInst2_LFInst_4_LFInst_0_U2 ( .A1(PermutationOutput2[19]), 
        .A2(PermutationOutput2[18]), .ZN(SubCellInst2_LFInst_4_LFInst_0_n11)
         );
  INV_X1 SubCellInst2_LFInst_4_LFInst_0_U1 ( .A(PermutationOutput2[16]), .ZN(
        SubCellInst2_LFInst_4_LFInst_0_n12) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_1_U4 ( .A1(
        SubCellInst2_LFInst_4_LFInst_1_n9), .A2(
        SubCellInst2_LFInst_4_LFInst_1_n8), .ZN(Output[17]) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_1_U3 ( .A1(PermutationOutput2[16]), 
        .A2(PermutationOutput2[18]), .ZN(SubCellInst2_LFInst_4_LFInst_1_n8) );
  OR2_X1 SubCellInst2_LFInst_4_LFInst_1_U2 ( .A1(PermutationOutput2[19]), .A2(
        SubCellInst2_LFInst_4_LFInst_1_n7), .ZN(
        SubCellInst2_LFInst_4_LFInst_1_n9) );
  NOR2_X1 SubCellInst2_LFInst_4_LFInst_1_U1 ( .A1(PermutationOutput2[16]), 
        .A2(PermutationOutput2[18]), .ZN(SubCellInst2_LFInst_4_LFInst_1_n7) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_2_U6 ( .A1(
        SubCellInst2_LFInst_4_LFInst_2_n18), .A2(
        SubCellInst2_LFInst_4_LFInst_2_n17), .ZN(Output[18]) );
  OR2_X1 SubCellInst2_LFInst_4_LFInst_2_U5 ( .A1(PermutationOutput2[16]), .A2(
        PermutationOutput2[19]), .ZN(SubCellInst2_LFInst_4_LFInst_2_n17) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_2_U4 ( .A1(PermutationOutput2[17]), 
        .A2(SubCellInst2_LFInst_4_LFInst_2_n16), .ZN(
        SubCellInst2_LFInst_4_LFInst_2_n18) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_2_U3 ( .A1(
        SubCellInst2_LFInst_4_LFInst_2_n15), .A2(
        SubCellInst2_LFInst_4_LFInst_2_n14), .ZN(
        SubCellInst2_LFInst_4_LFInst_2_n16) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_2_U2 ( .A1(PermutationOutput2[16]), 
        .A2(PermutationOutput2[19]), .ZN(SubCellInst2_LFInst_4_LFInst_2_n14)
         );
  INV_X1 SubCellInst2_LFInst_4_LFInst_2_U1 ( .A(PermutationOutput2[18]), .ZN(
        SubCellInst2_LFInst_4_LFInst_2_n15) );
  OR2_X1 SubCellInst2_LFInst_4_LFInst_3_U4 ( .A1(
        SubCellInst2_LFInst_4_LFInst_3_n9), .A2(
        SubCellInst2_LFInst_4_LFInst_3_n8), .ZN(Output[19]) );
  NOR2_X1 SubCellInst2_LFInst_4_LFInst_3_U3 ( .A1(PermutationOutput2[17]), 
        .A2(PermutationOutput2[18]), .ZN(SubCellInst2_LFInst_4_LFInst_3_n8) );
  NOR2_X1 SubCellInst2_LFInst_4_LFInst_3_U2 ( .A1(PermutationOutput2[19]), 
        .A2(SubCellInst2_LFInst_4_LFInst_3_n7), .ZN(
        SubCellInst2_LFInst_4_LFInst_3_n9) );
  AND2_X1 SubCellInst2_LFInst_4_LFInst_3_U1 ( .A1(PermutationOutput2[17]), 
        .A2(PermutationOutput2[16]), .ZN(SubCellInst2_LFInst_4_LFInst_3_n7) );
  NOR2_X1 SubCellInst2_LFInst_5_LFInst_0_U6 ( .A1(
        SubCellInst2_LFInst_5_LFInst_0_n15), .A2(
        SubCellInst2_LFInst_5_LFInst_0_n14), .ZN(Output[20]) );
  AND2_X1 SubCellInst2_LFInst_5_LFInst_0_U5 ( .A1(PermutationOutput2[23]), 
        .A2(PermutationOutput2[22]), .ZN(SubCellInst2_LFInst_5_LFInst_0_n14)
         );
  NOR2_X1 SubCellInst2_LFInst_5_LFInst_0_U4 ( .A1(PermutationOutput2[21]), 
        .A2(SubCellInst2_LFInst_5_LFInst_0_n13), .ZN(
        SubCellInst2_LFInst_5_LFInst_0_n15) );
  NOR2_X1 SubCellInst2_LFInst_5_LFInst_0_U3 ( .A1(
        SubCellInst2_LFInst_5_LFInst_0_n12), .A2(
        SubCellInst2_LFInst_5_LFInst_0_n11), .ZN(
        SubCellInst2_LFInst_5_LFInst_0_n13) );
  NOR2_X1 SubCellInst2_LFInst_5_LFInst_0_U2 ( .A1(PermutationOutput2[23]), 
        .A2(PermutationOutput2[22]), .ZN(SubCellInst2_LFInst_5_LFInst_0_n11)
         );
  INV_X1 SubCellInst2_LFInst_5_LFInst_0_U1 ( .A(PermutationOutput2[20]), .ZN(
        SubCellInst2_LFInst_5_LFInst_0_n12) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_1_U4 ( .A1(
        SubCellInst2_LFInst_5_LFInst_1_n9), .A2(
        SubCellInst2_LFInst_5_LFInst_1_n8), .ZN(Output[21]) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_1_U3 ( .A1(PermutationOutput2[20]), 
        .A2(PermutationOutput2[22]), .ZN(SubCellInst2_LFInst_5_LFInst_1_n8) );
  OR2_X1 SubCellInst2_LFInst_5_LFInst_1_U2 ( .A1(PermutationOutput2[23]), .A2(
        SubCellInst2_LFInst_5_LFInst_1_n7), .ZN(
        SubCellInst2_LFInst_5_LFInst_1_n9) );
  NOR2_X1 SubCellInst2_LFInst_5_LFInst_1_U1 ( .A1(PermutationOutput2[20]), 
        .A2(PermutationOutput2[22]), .ZN(SubCellInst2_LFInst_5_LFInst_1_n7) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_2_U6 ( .A1(
        SubCellInst2_LFInst_5_LFInst_2_n18), .A2(
        SubCellInst2_LFInst_5_LFInst_2_n17), .ZN(Output[22]) );
  OR2_X1 SubCellInst2_LFInst_5_LFInst_2_U5 ( .A1(PermutationOutput2[20]), .A2(
        PermutationOutput2[23]), .ZN(SubCellInst2_LFInst_5_LFInst_2_n17) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_2_U4 ( .A1(PermutationOutput2[21]), 
        .A2(SubCellInst2_LFInst_5_LFInst_2_n16), .ZN(
        SubCellInst2_LFInst_5_LFInst_2_n18) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_2_U3 ( .A1(
        SubCellInst2_LFInst_5_LFInst_2_n15), .A2(
        SubCellInst2_LFInst_5_LFInst_2_n14), .ZN(
        SubCellInst2_LFInst_5_LFInst_2_n16) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_2_U2 ( .A1(PermutationOutput2[20]), 
        .A2(PermutationOutput2[23]), .ZN(SubCellInst2_LFInst_5_LFInst_2_n14)
         );
  INV_X1 SubCellInst2_LFInst_5_LFInst_2_U1 ( .A(PermutationOutput2[22]), .ZN(
        SubCellInst2_LFInst_5_LFInst_2_n15) );
  OR2_X1 SubCellInst2_LFInst_5_LFInst_3_U4 ( .A1(
        SubCellInst2_LFInst_5_LFInst_3_n9), .A2(
        SubCellInst2_LFInst_5_LFInst_3_n8), .ZN(Output[23]) );
  NOR2_X1 SubCellInst2_LFInst_5_LFInst_3_U3 ( .A1(PermutationOutput2[21]), 
        .A2(PermutationOutput2[22]), .ZN(SubCellInst2_LFInst_5_LFInst_3_n8) );
  NOR2_X1 SubCellInst2_LFInst_5_LFInst_3_U2 ( .A1(PermutationOutput2[23]), 
        .A2(SubCellInst2_LFInst_5_LFInst_3_n7), .ZN(
        SubCellInst2_LFInst_5_LFInst_3_n9) );
  AND2_X1 SubCellInst2_LFInst_5_LFInst_3_U1 ( .A1(PermutationOutput2[21]), 
        .A2(PermutationOutput2[20]), .ZN(SubCellInst2_LFInst_5_LFInst_3_n7) );
  NOR2_X1 SubCellInst2_LFInst_6_LFInst_0_U6 ( .A1(
        SubCellInst2_LFInst_6_LFInst_0_n15), .A2(
        SubCellInst2_LFInst_6_LFInst_0_n14), .ZN(Output[24]) );
  AND2_X1 SubCellInst2_LFInst_6_LFInst_0_U5 ( .A1(PermutationOutput2[27]), 
        .A2(PermutationOutput2[26]), .ZN(SubCellInst2_LFInst_6_LFInst_0_n14)
         );
  NOR2_X1 SubCellInst2_LFInst_6_LFInst_0_U4 ( .A1(PermutationOutput2[25]), 
        .A2(SubCellInst2_LFInst_6_LFInst_0_n13), .ZN(
        SubCellInst2_LFInst_6_LFInst_0_n15) );
  NOR2_X1 SubCellInst2_LFInst_6_LFInst_0_U3 ( .A1(
        SubCellInst2_LFInst_6_LFInst_0_n12), .A2(
        SubCellInst2_LFInst_6_LFInst_0_n11), .ZN(
        SubCellInst2_LFInst_6_LFInst_0_n13) );
  NOR2_X1 SubCellInst2_LFInst_6_LFInst_0_U2 ( .A1(PermutationOutput2[27]), 
        .A2(PermutationOutput2[26]), .ZN(SubCellInst2_LFInst_6_LFInst_0_n11)
         );
  INV_X1 SubCellInst2_LFInst_6_LFInst_0_U1 ( .A(PermutationOutput2[24]), .ZN(
        SubCellInst2_LFInst_6_LFInst_0_n12) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_1_U4 ( .A1(
        SubCellInst2_LFInst_6_LFInst_1_n9), .A2(
        SubCellInst2_LFInst_6_LFInst_1_n8), .ZN(Output[25]) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_1_U3 ( .A1(PermutationOutput2[24]), 
        .A2(PermutationOutput2[26]), .ZN(SubCellInst2_LFInst_6_LFInst_1_n8) );
  OR2_X1 SubCellInst2_LFInst_6_LFInst_1_U2 ( .A1(PermutationOutput2[27]), .A2(
        SubCellInst2_LFInst_6_LFInst_1_n7), .ZN(
        SubCellInst2_LFInst_6_LFInst_1_n9) );
  NOR2_X1 SubCellInst2_LFInst_6_LFInst_1_U1 ( .A1(PermutationOutput2[24]), 
        .A2(PermutationOutput2[26]), .ZN(SubCellInst2_LFInst_6_LFInst_1_n7) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_2_U6 ( .A1(
        SubCellInst2_LFInst_6_LFInst_2_n18), .A2(
        SubCellInst2_LFInst_6_LFInst_2_n17), .ZN(Output[26]) );
  OR2_X1 SubCellInst2_LFInst_6_LFInst_2_U5 ( .A1(PermutationOutput2[24]), .A2(
        PermutationOutput2[27]), .ZN(SubCellInst2_LFInst_6_LFInst_2_n17) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_2_U4 ( .A1(PermutationOutput2[25]), 
        .A2(SubCellInst2_LFInst_6_LFInst_2_n16), .ZN(
        SubCellInst2_LFInst_6_LFInst_2_n18) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_2_U3 ( .A1(
        SubCellInst2_LFInst_6_LFInst_2_n15), .A2(
        SubCellInst2_LFInst_6_LFInst_2_n14), .ZN(
        SubCellInst2_LFInst_6_LFInst_2_n16) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_2_U2 ( .A1(PermutationOutput2[24]), 
        .A2(PermutationOutput2[27]), .ZN(SubCellInst2_LFInst_6_LFInst_2_n14)
         );
  INV_X1 SubCellInst2_LFInst_6_LFInst_2_U1 ( .A(PermutationOutput2[26]), .ZN(
        SubCellInst2_LFInst_6_LFInst_2_n15) );
  OR2_X1 SubCellInst2_LFInst_6_LFInst_3_U4 ( .A1(
        SubCellInst2_LFInst_6_LFInst_3_n9), .A2(
        SubCellInst2_LFInst_6_LFInst_3_n8), .ZN(Output[27]) );
  NOR2_X1 SubCellInst2_LFInst_6_LFInst_3_U3 ( .A1(PermutationOutput2[25]), 
        .A2(PermutationOutput2[26]), .ZN(SubCellInst2_LFInst_6_LFInst_3_n8) );
  NOR2_X1 SubCellInst2_LFInst_6_LFInst_3_U2 ( .A1(PermutationOutput2[27]), 
        .A2(SubCellInst2_LFInst_6_LFInst_3_n7), .ZN(
        SubCellInst2_LFInst_6_LFInst_3_n9) );
  AND2_X1 SubCellInst2_LFInst_6_LFInst_3_U1 ( .A1(PermutationOutput2[25]), 
        .A2(PermutationOutput2[24]), .ZN(SubCellInst2_LFInst_6_LFInst_3_n7) );
  NOR2_X1 SubCellInst2_LFInst_7_LFInst_0_U6 ( .A1(
        SubCellInst2_LFInst_7_LFInst_0_n15), .A2(
        SubCellInst2_LFInst_7_LFInst_0_n14), .ZN(Output[28]) );
  AND2_X1 SubCellInst2_LFInst_7_LFInst_0_U5 ( .A1(PermutationOutput2[31]), 
        .A2(PermutationOutput2[30]), .ZN(SubCellInst2_LFInst_7_LFInst_0_n14)
         );
  NOR2_X1 SubCellInst2_LFInst_7_LFInst_0_U4 ( .A1(PermutationOutput2[29]), 
        .A2(SubCellInst2_LFInst_7_LFInst_0_n13), .ZN(
        SubCellInst2_LFInst_7_LFInst_0_n15) );
  NOR2_X1 SubCellInst2_LFInst_7_LFInst_0_U3 ( .A1(
        SubCellInst2_LFInst_7_LFInst_0_n12), .A2(
        SubCellInst2_LFInst_7_LFInst_0_n11), .ZN(
        SubCellInst2_LFInst_7_LFInst_0_n13) );
  NOR2_X1 SubCellInst2_LFInst_7_LFInst_0_U2 ( .A1(PermutationOutput2[31]), 
        .A2(PermutationOutput2[30]), .ZN(SubCellInst2_LFInst_7_LFInst_0_n11)
         );
  INV_X1 SubCellInst2_LFInst_7_LFInst_0_U1 ( .A(PermutationOutput2[28]), .ZN(
        SubCellInst2_LFInst_7_LFInst_0_n12) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_1_U4 ( .A1(
        SubCellInst2_LFInst_7_LFInst_1_n9), .A2(
        SubCellInst2_LFInst_7_LFInst_1_n8), .ZN(Output[29]) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_1_U3 ( .A1(PermutationOutput2[28]), 
        .A2(PermutationOutput2[30]), .ZN(SubCellInst2_LFInst_7_LFInst_1_n8) );
  OR2_X1 SubCellInst2_LFInst_7_LFInst_1_U2 ( .A1(PermutationOutput2[31]), .A2(
        SubCellInst2_LFInst_7_LFInst_1_n7), .ZN(
        SubCellInst2_LFInst_7_LFInst_1_n9) );
  NOR2_X1 SubCellInst2_LFInst_7_LFInst_1_U1 ( .A1(PermutationOutput2[28]), 
        .A2(PermutationOutput2[30]), .ZN(SubCellInst2_LFInst_7_LFInst_1_n7) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_2_U6 ( .A1(
        SubCellInst2_LFInst_7_LFInst_2_n18), .A2(
        SubCellInst2_LFInst_7_LFInst_2_n17), .ZN(Output[30]) );
  OR2_X1 SubCellInst2_LFInst_7_LFInst_2_U5 ( .A1(PermutationOutput2[28]), .A2(
        PermutationOutput2[31]), .ZN(SubCellInst2_LFInst_7_LFInst_2_n17) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_2_U4 ( .A1(PermutationOutput2[29]), 
        .A2(SubCellInst2_LFInst_7_LFInst_2_n16), .ZN(
        SubCellInst2_LFInst_7_LFInst_2_n18) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_2_U3 ( .A1(
        SubCellInst2_LFInst_7_LFInst_2_n15), .A2(
        SubCellInst2_LFInst_7_LFInst_2_n14), .ZN(
        SubCellInst2_LFInst_7_LFInst_2_n16) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_2_U2 ( .A1(PermutationOutput2[28]), 
        .A2(PermutationOutput2[31]), .ZN(SubCellInst2_LFInst_7_LFInst_2_n14)
         );
  INV_X1 SubCellInst2_LFInst_7_LFInst_2_U1 ( .A(PermutationOutput2[30]), .ZN(
        SubCellInst2_LFInst_7_LFInst_2_n15) );
  OR2_X1 SubCellInst2_LFInst_7_LFInst_3_U4 ( .A1(
        SubCellInst2_LFInst_7_LFInst_3_n9), .A2(
        SubCellInst2_LFInst_7_LFInst_3_n8), .ZN(Output[31]) );
  NOR2_X1 SubCellInst2_LFInst_7_LFInst_3_U3 ( .A1(PermutationOutput2[29]), 
        .A2(PermutationOutput2[30]), .ZN(SubCellInst2_LFInst_7_LFInst_3_n8) );
  NOR2_X1 SubCellInst2_LFInst_7_LFInst_3_U2 ( .A1(PermutationOutput2[31]), 
        .A2(SubCellInst2_LFInst_7_LFInst_3_n7), .ZN(
        SubCellInst2_LFInst_7_LFInst_3_n9) );
  AND2_X1 SubCellInst2_LFInst_7_LFInst_3_U1 ( .A1(PermutationOutput2[29]), 
        .A2(PermutationOutput2[28]), .ZN(SubCellInst2_LFInst_7_LFInst_3_n7) );
  NOR2_X1 SubCellInst2_LFInst_8_LFInst_0_U6 ( .A1(
        SubCellInst2_LFInst_8_LFInst_0_n15), .A2(
        SubCellInst2_LFInst_8_LFInst_0_n14), .ZN(Output[32]) );
  AND2_X1 SubCellInst2_LFInst_8_LFInst_0_U5 ( .A1(PermutationOutput2[35]), 
        .A2(PermutationOutput2[34]), .ZN(SubCellInst2_LFInst_8_LFInst_0_n14)
         );
  NOR2_X1 SubCellInst2_LFInst_8_LFInst_0_U4 ( .A1(PermutationOutput2[33]), 
        .A2(SubCellInst2_LFInst_8_LFInst_0_n13), .ZN(
        SubCellInst2_LFInst_8_LFInst_0_n15) );
  NOR2_X1 SubCellInst2_LFInst_8_LFInst_0_U3 ( .A1(
        SubCellInst2_LFInst_8_LFInst_0_n12), .A2(
        SubCellInst2_LFInst_8_LFInst_0_n11), .ZN(
        SubCellInst2_LFInst_8_LFInst_0_n13) );
  NOR2_X1 SubCellInst2_LFInst_8_LFInst_0_U2 ( .A1(PermutationOutput2[35]), 
        .A2(PermutationOutput2[34]), .ZN(SubCellInst2_LFInst_8_LFInst_0_n11)
         );
  INV_X1 SubCellInst2_LFInst_8_LFInst_0_U1 ( .A(PermutationOutput2[32]), .ZN(
        SubCellInst2_LFInst_8_LFInst_0_n12) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_1_U4 ( .A1(
        SubCellInst2_LFInst_8_LFInst_1_n9), .A2(
        SubCellInst2_LFInst_8_LFInst_1_n8), .ZN(Output[33]) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_1_U3 ( .A1(PermutationOutput2[32]), 
        .A2(PermutationOutput2[34]), .ZN(SubCellInst2_LFInst_8_LFInst_1_n8) );
  OR2_X1 SubCellInst2_LFInst_8_LFInst_1_U2 ( .A1(PermutationOutput2[35]), .A2(
        SubCellInst2_LFInst_8_LFInst_1_n7), .ZN(
        SubCellInst2_LFInst_8_LFInst_1_n9) );
  NOR2_X1 SubCellInst2_LFInst_8_LFInst_1_U1 ( .A1(PermutationOutput2[32]), 
        .A2(PermutationOutput2[34]), .ZN(SubCellInst2_LFInst_8_LFInst_1_n7) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_2_U6 ( .A1(
        SubCellInst2_LFInst_8_LFInst_2_n18), .A2(
        SubCellInst2_LFInst_8_LFInst_2_n17), .ZN(Output[34]) );
  OR2_X1 SubCellInst2_LFInst_8_LFInst_2_U5 ( .A1(PermutationOutput2[32]), .A2(
        PermutationOutput2[35]), .ZN(SubCellInst2_LFInst_8_LFInst_2_n17) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_2_U4 ( .A1(PermutationOutput2[33]), 
        .A2(SubCellInst2_LFInst_8_LFInst_2_n16), .ZN(
        SubCellInst2_LFInst_8_LFInst_2_n18) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_2_U3 ( .A1(
        SubCellInst2_LFInst_8_LFInst_2_n15), .A2(
        SubCellInst2_LFInst_8_LFInst_2_n14), .ZN(
        SubCellInst2_LFInst_8_LFInst_2_n16) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_2_U2 ( .A1(PermutationOutput2[32]), 
        .A2(PermutationOutput2[35]), .ZN(SubCellInst2_LFInst_8_LFInst_2_n14)
         );
  INV_X1 SubCellInst2_LFInst_8_LFInst_2_U1 ( .A(PermutationOutput2[34]), .ZN(
        SubCellInst2_LFInst_8_LFInst_2_n15) );
  OR2_X1 SubCellInst2_LFInst_8_LFInst_3_U4 ( .A1(
        SubCellInst2_LFInst_8_LFInst_3_n9), .A2(
        SubCellInst2_LFInst_8_LFInst_3_n8), .ZN(Output[35]) );
  NOR2_X1 SubCellInst2_LFInst_8_LFInst_3_U3 ( .A1(PermutationOutput2[33]), 
        .A2(PermutationOutput2[34]), .ZN(SubCellInst2_LFInst_8_LFInst_3_n8) );
  NOR2_X1 SubCellInst2_LFInst_8_LFInst_3_U2 ( .A1(PermutationOutput2[35]), 
        .A2(SubCellInst2_LFInst_8_LFInst_3_n7), .ZN(
        SubCellInst2_LFInst_8_LFInst_3_n9) );
  AND2_X1 SubCellInst2_LFInst_8_LFInst_3_U1 ( .A1(PermutationOutput2[33]), 
        .A2(PermutationOutput2[32]), .ZN(SubCellInst2_LFInst_8_LFInst_3_n7) );
  NOR2_X1 SubCellInst2_LFInst_9_LFInst_0_U6 ( .A1(
        SubCellInst2_LFInst_9_LFInst_0_n15), .A2(
        SubCellInst2_LFInst_9_LFInst_0_n14), .ZN(Output[36]) );
  AND2_X1 SubCellInst2_LFInst_9_LFInst_0_U5 ( .A1(PermutationOutput2[39]), 
        .A2(PermutationOutput2[38]), .ZN(SubCellInst2_LFInst_9_LFInst_0_n14)
         );
  NOR2_X1 SubCellInst2_LFInst_9_LFInst_0_U4 ( .A1(PermutationOutput2[37]), 
        .A2(SubCellInst2_LFInst_9_LFInst_0_n13), .ZN(
        SubCellInst2_LFInst_9_LFInst_0_n15) );
  NOR2_X1 SubCellInst2_LFInst_9_LFInst_0_U3 ( .A1(
        SubCellInst2_LFInst_9_LFInst_0_n12), .A2(
        SubCellInst2_LFInst_9_LFInst_0_n11), .ZN(
        SubCellInst2_LFInst_9_LFInst_0_n13) );
  NOR2_X1 SubCellInst2_LFInst_9_LFInst_0_U2 ( .A1(PermutationOutput2[39]), 
        .A2(PermutationOutput2[38]), .ZN(SubCellInst2_LFInst_9_LFInst_0_n11)
         );
  INV_X1 SubCellInst2_LFInst_9_LFInst_0_U1 ( .A(PermutationOutput2[36]), .ZN(
        SubCellInst2_LFInst_9_LFInst_0_n12) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_1_U4 ( .A1(
        SubCellInst2_LFInst_9_LFInst_1_n9), .A2(
        SubCellInst2_LFInst_9_LFInst_1_n8), .ZN(Output[37]) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_1_U3 ( .A1(PermutationOutput2[36]), 
        .A2(PermutationOutput2[38]), .ZN(SubCellInst2_LFInst_9_LFInst_1_n8) );
  OR2_X1 SubCellInst2_LFInst_9_LFInst_1_U2 ( .A1(PermutationOutput2[39]), .A2(
        SubCellInst2_LFInst_9_LFInst_1_n7), .ZN(
        SubCellInst2_LFInst_9_LFInst_1_n9) );
  NOR2_X1 SubCellInst2_LFInst_9_LFInst_1_U1 ( .A1(PermutationOutput2[36]), 
        .A2(PermutationOutput2[38]), .ZN(SubCellInst2_LFInst_9_LFInst_1_n7) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_2_U6 ( .A1(
        SubCellInst2_LFInst_9_LFInst_2_n18), .A2(
        SubCellInst2_LFInst_9_LFInst_2_n17), .ZN(Output[38]) );
  OR2_X1 SubCellInst2_LFInst_9_LFInst_2_U5 ( .A1(PermutationOutput2[36]), .A2(
        PermutationOutput2[39]), .ZN(SubCellInst2_LFInst_9_LFInst_2_n17) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_2_U4 ( .A1(PermutationOutput2[37]), 
        .A2(SubCellInst2_LFInst_9_LFInst_2_n16), .ZN(
        SubCellInst2_LFInst_9_LFInst_2_n18) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_2_U3 ( .A1(
        SubCellInst2_LFInst_9_LFInst_2_n15), .A2(
        SubCellInst2_LFInst_9_LFInst_2_n14), .ZN(
        SubCellInst2_LFInst_9_LFInst_2_n16) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_2_U2 ( .A1(PermutationOutput2[36]), 
        .A2(PermutationOutput2[39]), .ZN(SubCellInst2_LFInst_9_LFInst_2_n14)
         );
  INV_X1 SubCellInst2_LFInst_9_LFInst_2_U1 ( .A(PermutationOutput2[38]), .ZN(
        SubCellInst2_LFInst_9_LFInst_2_n15) );
  OR2_X1 SubCellInst2_LFInst_9_LFInst_3_U4 ( .A1(
        SubCellInst2_LFInst_9_LFInst_3_n9), .A2(
        SubCellInst2_LFInst_9_LFInst_3_n8), .ZN(Output[39]) );
  NOR2_X1 SubCellInst2_LFInst_9_LFInst_3_U3 ( .A1(PermutationOutput2[37]), 
        .A2(PermutationOutput2[38]), .ZN(SubCellInst2_LFInst_9_LFInst_3_n8) );
  NOR2_X1 SubCellInst2_LFInst_9_LFInst_3_U2 ( .A1(PermutationOutput2[39]), 
        .A2(SubCellInst2_LFInst_9_LFInst_3_n7), .ZN(
        SubCellInst2_LFInst_9_LFInst_3_n9) );
  AND2_X1 SubCellInst2_LFInst_9_LFInst_3_U1 ( .A1(PermutationOutput2[37]), 
        .A2(PermutationOutput2[36]), .ZN(SubCellInst2_LFInst_9_LFInst_3_n7) );
  NOR2_X1 SubCellInst2_LFInst_10_LFInst_0_U6 ( .A1(
        SubCellInst2_LFInst_10_LFInst_0_n15), .A2(
        SubCellInst2_LFInst_10_LFInst_0_n14), .ZN(Output[40]) );
  AND2_X1 SubCellInst2_LFInst_10_LFInst_0_U5 ( .A1(PermutationOutput2[43]), 
        .A2(PermutationOutput2[42]), .ZN(SubCellInst2_LFInst_10_LFInst_0_n14)
         );
  NOR2_X1 SubCellInst2_LFInst_10_LFInst_0_U4 ( .A1(PermutationOutput2[41]), 
        .A2(SubCellInst2_LFInst_10_LFInst_0_n13), .ZN(
        SubCellInst2_LFInst_10_LFInst_0_n15) );
  NOR2_X1 SubCellInst2_LFInst_10_LFInst_0_U3 ( .A1(
        SubCellInst2_LFInst_10_LFInst_0_n12), .A2(
        SubCellInst2_LFInst_10_LFInst_0_n11), .ZN(
        SubCellInst2_LFInst_10_LFInst_0_n13) );
  NOR2_X1 SubCellInst2_LFInst_10_LFInst_0_U2 ( .A1(PermutationOutput2[43]), 
        .A2(PermutationOutput2[42]), .ZN(SubCellInst2_LFInst_10_LFInst_0_n11)
         );
  INV_X1 SubCellInst2_LFInst_10_LFInst_0_U1 ( .A(PermutationOutput2[40]), .ZN(
        SubCellInst2_LFInst_10_LFInst_0_n12) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_1_U4 ( .A1(
        SubCellInst2_LFInst_10_LFInst_1_n9), .A2(
        SubCellInst2_LFInst_10_LFInst_1_n8), .ZN(Output[41]) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_1_U3 ( .A1(PermutationOutput2[40]), 
        .A2(PermutationOutput2[42]), .ZN(SubCellInst2_LFInst_10_LFInst_1_n8)
         );
  OR2_X1 SubCellInst2_LFInst_10_LFInst_1_U2 ( .A1(PermutationOutput2[43]), 
        .A2(SubCellInst2_LFInst_10_LFInst_1_n7), .ZN(
        SubCellInst2_LFInst_10_LFInst_1_n9) );
  NOR2_X1 SubCellInst2_LFInst_10_LFInst_1_U1 ( .A1(PermutationOutput2[40]), 
        .A2(PermutationOutput2[42]), .ZN(SubCellInst2_LFInst_10_LFInst_1_n7)
         );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_2_U6 ( .A1(
        SubCellInst2_LFInst_10_LFInst_2_n18), .A2(
        SubCellInst2_LFInst_10_LFInst_2_n17), .ZN(Output[42]) );
  OR2_X1 SubCellInst2_LFInst_10_LFInst_2_U5 ( .A1(PermutationOutput2[40]), 
        .A2(PermutationOutput2[43]), .ZN(SubCellInst2_LFInst_10_LFInst_2_n17)
         );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_2_U4 ( .A1(PermutationOutput2[41]), 
        .A2(SubCellInst2_LFInst_10_LFInst_2_n16), .ZN(
        SubCellInst2_LFInst_10_LFInst_2_n18) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_2_U3 ( .A1(
        SubCellInst2_LFInst_10_LFInst_2_n15), .A2(
        SubCellInst2_LFInst_10_LFInst_2_n14), .ZN(
        SubCellInst2_LFInst_10_LFInst_2_n16) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_2_U2 ( .A1(PermutationOutput2[40]), 
        .A2(PermutationOutput2[43]), .ZN(SubCellInst2_LFInst_10_LFInst_2_n14)
         );
  INV_X1 SubCellInst2_LFInst_10_LFInst_2_U1 ( .A(PermutationOutput2[42]), .ZN(
        SubCellInst2_LFInst_10_LFInst_2_n15) );
  OR2_X1 SubCellInst2_LFInst_10_LFInst_3_U4 ( .A1(
        SubCellInst2_LFInst_10_LFInst_3_n9), .A2(
        SubCellInst2_LFInst_10_LFInst_3_n8), .ZN(Output[43]) );
  NOR2_X1 SubCellInst2_LFInst_10_LFInst_3_U3 ( .A1(PermutationOutput2[41]), 
        .A2(PermutationOutput2[42]), .ZN(SubCellInst2_LFInst_10_LFInst_3_n8)
         );
  NOR2_X1 SubCellInst2_LFInst_10_LFInst_3_U2 ( .A1(PermutationOutput2[43]), 
        .A2(SubCellInst2_LFInst_10_LFInst_3_n7), .ZN(
        SubCellInst2_LFInst_10_LFInst_3_n9) );
  AND2_X1 SubCellInst2_LFInst_10_LFInst_3_U1 ( .A1(PermutationOutput2[41]), 
        .A2(PermutationOutput2[40]), .ZN(SubCellInst2_LFInst_10_LFInst_3_n7)
         );
  NOR2_X1 SubCellInst2_LFInst_11_LFInst_0_U6 ( .A1(
        SubCellInst2_LFInst_11_LFInst_0_n15), .A2(
        SubCellInst2_LFInst_11_LFInst_0_n14), .ZN(Output[44]) );
  AND2_X1 SubCellInst2_LFInst_11_LFInst_0_U5 ( .A1(PermutationOutput2[47]), 
        .A2(PermutationOutput2[46]), .ZN(SubCellInst2_LFInst_11_LFInst_0_n14)
         );
  NOR2_X1 SubCellInst2_LFInst_11_LFInst_0_U4 ( .A1(PermutationOutput2[45]), 
        .A2(SubCellInst2_LFInst_11_LFInst_0_n13), .ZN(
        SubCellInst2_LFInst_11_LFInst_0_n15) );
  NOR2_X1 SubCellInst2_LFInst_11_LFInst_0_U3 ( .A1(
        SubCellInst2_LFInst_11_LFInst_0_n12), .A2(
        SubCellInst2_LFInst_11_LFInst_0_n11), .ZN(
        SubCellInst2_LFInst_11_LFInst_0_n13) );
  NOR2_X1 SubCellInst2_LFInst_11_LFInst_0_U2 ( .A1(PermutationOutput2[47]), 
        .A2(PermutationOutput2[46]), .ZN(SubCellInst2_LFInst_11_LFInst_0_n11)
         );
  INV_X1 SubCellInst2_LFInst_11_LFInst_0_U1 ( .A(PermutationOutput2[44]), .ZN(
        SubCellInst2_LFInst_11_LFInst_0_n12) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_1_U4 ( .A1(
        SubCellInst2_LFInst_11_LFInst_1_n9), .A2(
        SubCellInst2_LFInst_11_LFInst_1_n8), .ZN(Output[45]) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_1_U3 ( .A1(PermutationOutput2[44]), 
        .A2(PermutationOutput2[46]), .ZN(SubCellInst2_LFInst_11_LFInst_1_n8)
         );
  OR2_X1 SubCellInst2_LFInst_11_LFInst_1_U2 ( .A1(PermutationOutput2[47]), 
        .A2(SubCellInst2_LFInst_11_LFInst_1_n7), .ZN(
        SubCellInst2_LFInst_11_LFInst_1_n9) );
  NOR2_X1 SubCellInst2_LFInst_11_LFInst_1_U1 ( .A1(PermutationOutput2[44]), 
        .A2(PermutationOutput2[46]), .ZN(SubCellInst2_LFInst_11_LFInst_1_n7)
         );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_2_U6 ( .A1(
        SubCellInst2_LFInst_11_LFInst_2_n18), .A2(
        SubCellInst2_LFInst_11_LFInst_2_n17), .ZN(Output[46]) );
  OR2_X1 SubCellInst2_LFInst_11_LFInst_2_U5 ( .A1(PermutationOutput2[44]), 
        .A2(PermutationOutput2[47]), .ZN(SubCellInst2_LFInst_11_LFInst_2_n17)
         );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_2_U4 ( .A1(PermutationOutput2[45]), 
        .A2(SubCellInst2_LFInst_11_LFInst_2_n16), .ZN(
        SubCellInst2_LFInst_11_LFInst_2_n18) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_2_U3 ( .A1(
        SubCellInst2_LFInst_11_LFInst_2_n15), .A2(
        SubCellInst2_LFInst_11_LFInst_2_n14), .ZN(
        SubCellInst2_LFInst_11_LFInst_2_n16) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_2_U2 ( .A1(PermutationOutput2[44]), 
        .A2(PermutationOutput2[47]), .ZN(SubCellInst2_LFInst_11_LFInst_2_n14)
         );
  INV_X1 SubCellInst2_LFInst_11_LFInst_2_U1 ( .A(PermutationOutput2[46]), .ZN(
        SubCellInst2_LFInst_11_LFInst_2_n15) );
  OR2_X1 SubCellInst2_LFInst_11_LFInst_3_U4 ( .A1(
        SubCellInst2_LFInst_11_LFInst_3_n9), .A2(
        SubCellInst2_LFInst_11_LFInst_3_n8), .ZN(Output[47]) );
  NOR2_X1 SubCellInst2_LFInst_11_LFInst_3_U3 ( .A1(PermutationOutput2[45]), 
        .A2(PermutationOutput2[46]), .ZN(SubCellInst2_LFInst_11_LFInst_3_n8)
         );
  NOR2_X1 SubCellInst2_LFInst_11_LFInst_3_U2 ( .A1(PermutationOutput2[47]), 
        .A2(SubCellInst2_LFInst_11_LFInst_3_n7), .ZN(
        SubCellInst2_LFInst_11_LFInst_3_n9) );
  AND2_X1 SubCellInst2_LFInst_11_LFInst_3_U1 ( .A1(PermutationOutput2[45]), 
        .A2(PermutationOutput2[44]), .ZN(SubCellInst2_LFInst_11_LFInst_3_n7)
         );
  NOR2_X1 SubCellInst2_LFInst_12_LFInst_0_U6 ( .A1(
        SubCellInst2_LFInst_12_LFInst_0_n15), .A2(
        SubCellInst2_LFInst_12_LFInst_0_n14), .ZN(Output[48]) );
  AND2_X1 SubCellInst2_LFInst_12_LFInst_0_U5 ( .A1(PermutationOutput2[51]), 
        .A2(PermutationOutput2[50]), .ZN(SubCellInst2_LFInst_12_LFInst_0_n14)
         );
  NOR2_X1 SubCellInst2_LFInst_12_LFInst_0_U4 ( .A1(PermutationOutput2[49]), 
        .A2(SubCellInst2_LFInst_12_LFInst_0_n13), .ZN(
        SubCellInst2_LFInst_12_LFInst_0_n15) );
  NOR2_X1 SubCellInst2_LFInst_12_LFInst_0_U3 ( .A1(
        SubCellInst2_LFInst_12_LFInst_0_n12), .A2(
        SubCellInst2_LFInst_12_LFInst_0_n11), .ZN(
        SubCellInst2_LFInst_12_LFInst_0_n13) );
  NOR2_X1 SubCellInst2_LFInst_12_LFInst_0_U2 ( .A1(PermutationOutput2[51]), 
        .A2(PermutationOutput2[50]), .ZN(SubCellInst2_LFInst_12_LFInst_0_n11)
         );
  INV_X1 SubCellInst2_LFInst_12_LFInst_0_U1 ( .A(PermutationOutput2[48]), .ZN(
        SubCellInst2_LFInst_12_LFInst_0_n12) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_1_U4 ( .A1(
        SubCellInst2_LFInst_12_LFInst_1_n9), .A2(
        SubCellInst2_LFInst_12_LFInst_1_n8), .ZN(Output[49]) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_1_U3 ( .A1(PermutationOutput2[48]), 
        .A2(PermutationOutput2[50]), .ZN(SubCellInst2_LFInst_12_LFInst_1_n8)
         );
  OR2_X1 SubCellInst2_LFInst_12_LFInst_1_U2 ( .A1(PermutationOutput2[51]), 
        .A2(SubCellInst2_LFInst_12_LFInst_1_n7), .ZN(
        SubCellInst2_LFInst_12_LFInst_1_n9) );
  NOR2_X1 SubCellInst2_LFInst_12_LFInst_1_U1 ( .A1(PermutationOutput2[48]), 
        .A2(PermutationOutput2[50]), .ZN(SubCellInst2_LFInst_12_LFInst_1_n7)
         );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_2_U6 ( .A1(
        SubCellInst2_LFInst_12_LFInst_2_n18), .A2(
        SubCellInst2_LFInst_12_LFInst_2_n17), .ZN(Output[50]) );
  OR2_X1 SubCellInst2_LFInst_12_LFInst_2_U5 ( .A1(PermutationOutput2[48]), 
        .A2(PermutationOutput2[51]), .ZN(SubCellInst2_LFInst_12_LFInst_2_n17)
         );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_2_U4 ( .A1(PermutationOutput2[49]), 
        .A2(SubCellInst2_LFInst_12_LFInst_2_n16), .ZN(
        SubCellInst2_LFInst_12_LFInst_2_n18) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_2_U3 ( .A1(
        SubCellInst2_LFInst_12_LFInst_2_n15), .A2(
        SubCellInst2_LFInst_12_LFInst_2_n14), .ZN(
        SubCellInst2_LFInst_12_LFInst_2_n16) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_2_U2 ( .A1(PermutationOutput2[48]), 
        .A2(PermutationOutput2[51]), .ZN(SubCellInst2_LFInst_12_LFInst_2_n14)
         );
  INV_X1 SubCellInst2_LFInst_12_LFInst_2_U1 ( .A(PermutationOutput2[50]), .ZN(
        SubCellInst2_LFInst_12_LFInst_2_n15) );
  OR2_X1 SubCellInst2_LFInst_12_LFInst_3_U4 ( .A1(
        SubCellInst2_LFInst_12_LFInst_3_n9), .A2(
        SubCellInst2_LFInst_12_LFInst_3_n8), .ZN(Output[51]) );
  NOR2_X1 SubCellInst2_LFInst_12_LFInst_3_U3 ( .A1(PermutationOutput2[49]), 
        .A2(PermutationOutput2[50]), .ZN(SubCellInst2_LFInst_12_LFInst_3_n8)
         );
  NOR2_X1 SubCellInst2_LFInst_12_LFInst_3_U2 ( .A1(PermutationOutput2[51]), 
        .A2(SubCellInst2_LFInst_12_LFInst_3_n7), .ZN(
        SubCellInst2_LFInst_12_LFInst_3_n9) );
  AND2_X1 SubCellInst2_LFInst_12_LFInst_3_U1 ( .A1(PermutationOutput2[49]), 
        .A2(PermutationOutput2[48]), .ZN(SubCellInst2_LFInst_12_LFInst_3_n7)
         );
  NOR2_X1 SubCellInst2_LFInst_13_LFInst_0_U6 ( .A1(
        SubCellInst2_LFInst_13_LFInst_0_n15), .A2(
        SubCellInst2_LFInst_13_LFInst_0_n14), .ZN(Output[52]) );
  AND2_X1 SubCellInst2_LFInst_13_LFInst_0_U5 ( .A1(PermutationOutput2[55]), 
        .A2(PermutationOutput2[54]), .ZN(SubCellInst2_LFInst_13_LFInst_0_n14)
         );
  NOR2_X1 SubCellInst2_LFInst_13_LFInst_0_U4 ( .A1(PermutationOutput2[53]), 
        .A2(SubCellInst2_LFInst_13_LFInst_0_n13), .ZN(
        SubCellInst2_LFInst_13_LFInst_0_n15) );
  NOR2_X1 SubCellInst2_LFInst_13_LFInst_0_U3 ( .A1(
        SubCellInst2_LFInst_13_LFInst_0_n12), .A2(
        SubCellInst2_LFInst_13_LFInst_0_n11), .ZN(
        SubCellInst2_LFInst_13_LFInst_0_n13) );
  NOR2_X1 SubCellInst2_LFInst_13_LFInst_0_U2 ( .A1(PermutationOutput2[55]), 
        .A2(PermutationOutput2[54]), .ZN(SubCellInst2_LFInst_13_LFInst_0_n11)
         );
  INV_X1 SubCellInst2_LFInst_13_LFInst_0_U1 ( .A(PermutationOutput2[52]), .ZN(
        SubCellInst2_LFInst_13_LFInst_0_n12) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_1_U4 ( .A1(
        SubCellInst2_LFInst_13_LFInst_1_n9), .A2(
        SubCellInst2_LFInst_13_LFInst_1_n8), .ZN(Output[53]) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_1_U3 ( .A1(PermutationOutput2[52]), 
        .A2(PermutationOutput2[54]), .ZN(SubCellInst2_LFInst_13_LFInst_1_n8)
         );
  OR2_X1 SubCellInst2_LFInst_13_LFInst_1_U2 ( .A1(PermutationOutput2[55]), 
        .A2(SubCellInst2_LFInst_13_LFInst_1_n7), .ZN(
        SubCellInst2_LFInst_13_LFInst_1_n9) );
  NOR2_X1 SubCellInst2_LFInst_13_LFInst_1_U1 ( .A1(PermutationOutput2[52]), 
        .A2(PermutationOutput2[54]), .ZN(SubCellInst2_LFInst_13_LFInst_1_n7)
         );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_2_U6 ( .A1(
        SubCellInst2_LFInst_13_LFInst_2_n18), .A2(
        SubCellInst2_LFInst_13_LFInst_2_n17), .ZN(Output[54]) );
  OR2_X1 SubCellInst2_LFInst_13_LFInst_2_U5 ( .A1(PermutationOutput2[52]), 
        .A2(PermutationOutput2[55]), .ZN(SubCellInst2_LFInst_13_LFInst_2_n17)
         );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_2_U4 ( .A1(PermutationOutput2[53]), 
        .A2(SubCellInst2_LFInst_13_LFInst_2_n16), .ZN(
        SubCellInst2_LFInst_13_LFInst_2_n18) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_2_U3 ( .A1(
        SubCellInst2_LFInst_13_LFInst_2_n15), .A2(
        SubCellInst2_LFInst_13_LFInst_2_n14), .ZN(
        SubCellInst2_LFInst_13_LFInst_2_n16) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_2_U2 ( .A1(PermutationOutput2[52]), 
        .A2(PermutationOutput2[55]), .ZN(SubCellInst2_LFInst_13_LFInst_2_n14)
         );
  INV_X1 SubCellInst2_LFInst_13_LFInst_2_U1 ( .A(PermutationOutput2[54]), .ZN(
        SubCellInst2_LFInst_13_LFInst_2_n15) );
  OR2_X1 SubCellInst2_LFInst_13_LFInst_3_U4 ( .A1(
        SubCellInst2_LFInst_13_LFInst_3_n9), .A2(
        SubCellInst2_LFInst_13_LFInst_3_n8), .ZN(Output[55]) );
  NOR2_X1 SubCellInst2_LFInst_13_LFInst_3_U3 ( .A1(PermutationOutput2[53]), 
        .A2(PermutationOutput2[54]), .ZN(SubCellInst2_LFInst_13_LFInst_3_n8)
         );
  NOR2_X1 SubCellInst2_LFInst_13_LFInst_3_U2 ( .A1(PermutationOutput2[55]), 
        .A2(SubCellInst2_LFInst_13_LFInst_3_n7), .ZN(
        SubCellInst2_LFInst_13_LFInst_3_n9) );
  AND2_X1 SubCellInst2_LFInst_13_LFInst_3_U1 ( .A1(PermutationOutput2[53]), 
        .A2(PermutationOutput2[52]), .ZN(SubCellInst2_LFInst_13_LFInst_3_n7)
         );
  NOR2_X1 SubCellInst2_LFInst_14_LFInst_0_U6 ( .A1(
        SubCellInst2_LFInst_14_LFInst_0_n15), .A2(
        SubCellInst2_LFInst_14_LFInst_0_n14), .ZN(Output[56]) );
  AND2_X1 SubCellInst2_LFInst_14_LFInst_0_U5 ( .A1(PermutationOutput2[59]), 
        .A2(PermutationOutput2[58]), .ZN(SubCellInst2_LFInst_14_LFInst_0_n14)
         );
  NOR2_X1 SubCellInst2_LFInst_14_LFInst_0_U4 ( .A1(PermutationOutput2[57]), 
        .A2(SubCellInst2_LFInst_14_LFInst_0_n13), .ZN(
        SubCellInst2_LFInst_14_LFInst_0_n15) );
  NOR2_X1 SubCellInst2_LFInst_14_LFInst_0_U3 ( .A1(
        SubCellInst2_LFInst_14_LFInst_0_n12), .A2(
        SubCellInst2_LFInst_14_LFInst_0_n11), .ZN(
        SubCellInst2_LFInst_14_LFInst_0_n13) );
  NOR2_X1 SubCellInst2_LFInst_14_LFInst_0_U2 ( .A1(PermutationOutput2[59]), 
        .A2(PermutationOutput2[58]), .ZN(SubCellInst2_LFInst_14_LFInst_0_n11)
         );
  INV_X1 SubCellInst2_LFInst_14_LFInst_0_U1 ( .A(PermutationOutput2[56]), .ZN(
        SubCellInst2_LFInst_14_LFInst_0_n12) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_1_U4 ( .A1(
        SubCellInst2_LFInst_14_LFInst_1_n9), .A2(
        SubCellInst2_LFInst_14_LFInst_1_n8), .ZN(Output[57]) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_1_U3 ( .A1(PermutationOutput2[56]), 
        .A2(PermutationOutput2[58]), .ZN(SubCellInst2_LFInst_14_LFInst_1_n8)
         );
  OR2_X1 SubCellInst2_LFInst_14_LFInst_1_U2 ( .A1(PermutationOutput2[59]), 
        .A2(SubCellInst2_LFInst_14_LFInst_1_n7), .ZN(
        SubCellInst2_LFInst_14_LFInst_1_n9) );
  NOR2_X1 SubCellInst2_LFInst_14_LFInst_1_U1 ( .A1(PermutationOutput2[56]), 
        .A2(PermutationOutput2[58]), .ZN(SubCellInst2_LFInst_14_LFInst_1_n7)
         );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_2_U6 ( .A1(
        SubCellInst2_LFInst_14_LFInst_2_n18), .A2(
        SubCellInst2_LFInst_14_LFInst_2_n17), .ZN(Output[58]) );
  OR2_X1 SubCellInst2_LFInst_14_LFInst_2_U5 ( .A1(PermutationOutput2[56]), 
        .A2(PermutationOutput2[59]), .ZN(SubCellInst2_LFInst_14_LFInst_2_n17)
         );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_2_U4 ( .A1(PermutationOutput2[57]), 
        .A2(SubCellInst2_LFInst_14_LFInst_2_n16), .ZN(
        SubCellInst2_LFInst_14_LFInst_2_n18) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_2_U3 ( .A1(
        SubCellInst2_LFInst_14_LFInst_2_n15), .A2(
        SubCellInst2_LFInst_14_LFInst_2_n14), .ZN(
        SubCellInst2_LFInst_14_LFInst_2_n16) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_2_U2 ( .A1(PermutationOutput2[56]), 
        .A2(PermutationOutput2[59]), .ZN(SubCellInst2_LFInst_14_LFInst_2_n14)
         );
  INV_X1 SubCellInst2_LFInst_14_LFInst_2_U1 ( .A(PermutationOutput2[58]), .ZN(
        SubCellInst2_LFInst_14_LFInst_2_n15) );
  OR2_X1 SubCellInst2_LFInst_14_LFInst_3_U4 ( .A1(
        SubCellInst2_LFInst_14_LFInst_3_n9), .A2(
        SubCellInst2_LFInst_14_LFInst_3_n8), .ZN(Output[59]) );
  NOR2_X1 SubCellInst2_LFInst_14_LFInst_3_U3 ( .A1(PermutationOutput2[57]), 
        .A2(PermutationOutput2[58]), .ZN(SubCellInst2_LFInst_14_LFInst_3_n8)
         );
  NOR2_X1 SubCellInst2_LFInst_14_LFInst_3_U2 ( .A1(PermutationOutput2[59]), 
        .A2(SubCellInst2_LFInst_14_LFInst_3_n7), .ZN(
        SubCellInst2_LFInst_14_LFInst_3_n9) );
  AND2_X1 SubCellInst2_LFInst_14_LFInst_3_U1 ( .A1(PermutationOutput2[57]), 
        .A2(PermutationOutput2[56]), .ZN(SubCellInst2_LFInst_14_LFInst_3_n7)
         );
  NOR2_X1 SubCellInst2_LFInst_15_LFInst_0_U6 ( .A1(
        SubCellInst2_LFInst_15_LFInst_0_n15), .A2(
        SubCellInst2_LFInst_15_LFInst_0_n14), .ZN(Output[60]) );
  AND2_X1 SubCellInst2_LFInst_15_LFInst_0_U5 ( .A1(PermutationOutput2[63]), 
        .A2(PermutationOutput2[62]), .ZN(SubCellInst2_LFInst_15_LFInst_0_n14)
         );
  NOR2_X1 SubCellInst2_LFInst_15_LFInst_0_U4 ( .A1(PermutationOutput2[61]), 
        .A2(SubCellInst2_LFInst_15_LFInst_0_n13), .ZN(
        SubCellInst2_LFInst_15_LFInst_0_n15) );
  NOR2_X1 SubCellInst2_LFInst_15_LFInst_0_U3 ( .A1(
        SubCellInst2_LFInst_15_LFInst_0_n12), .A2(
        SubCellInst2_LFInst_15_LFInst_0_n11), .ZN(
        SubCellInst2_LFInst_15_LFInst_0_n13) );
  NOR2_X1 SubCellInst2_LFInst_15_LFInst_0_U2 ( .A1(PermutationOutput2[63]), 
        .A2(PermutationOutput2[62]), .ZN(SubCellInst2_LFInst_15_LFInst_0_n11)
         );
  INV_X1 SubCellInst2_LFInst_15_LFInst_0_U1 ( .A(PermutationOutput2[60]), .ZN(
        SubCellInst2_LFInst_15_LFInst_0_n12) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_1_U4 ( .A1(
        SubCellInst2_LFInst_15_LFInst_1_n9), .A2(
        SubCellInst2_LFInst_15_LFInst_1_n8), .ZN(Output[61]) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_1_U3 ( .A1(PermutationOutput2[60]), 
        .A2(PermutationOutput2[62]), .ZN(SubCellInst2_LFInst_15_LFInst_1_n8)
         );
  OR2_X1 SubCellInst2_LFInst_15_LFInst_1_U2 ( .A1(PermutationOutput2[63]), 
        .A2(SubCellInst2_LFInst_15_LFInst_1_n7), .ZN(
        SubCellInst2_LFInst_15_LFInst_1_n9) );
  NOR2_X1 SubCellInst2_LFInst_15_LFInst_1_U1 ( .A1(PermutationOutput2[60]), 
        .A2(PermutationOutput2[62]), .ZN(SubCellInst2_LFInst_15_LFInst_1_n7)
         );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_2_U6 ( .A1(
        SubCellInst2_LFInst_15_LFInst_2_n18), .A2(
        SubCellInst2_LFInst_15_LFInst_2_n17), .ZN(Output[62]) );
  OR2_X1 SubCellInst2_LFInst_15_LFInst_2_U5 ( .A1(PermutationOutput2[60]), 
        .A2(PermutationOutput2[63]), .ZN(SubCellInst2_LFInst_15_LFInst_2_n17)
         );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_2_U4 ( .A1(PermutationOutput2[61]), 
        .A2(SubCellInst2_LFInst_15_LFInst_2_n16), .ZN(
        SubCellInst2_LFInst_15_LFInst_2_n18) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_2_U3 ( .A1(
        SubCellInst2_LFInst_15_LFInst_2_n15), .A2(
        SubCellInst2_LFInst_15_LFInst_2_n14), .ZN(
        SubCellInst2_LFInst_15_LFInst_2_n16) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_2_U2 ( .A1(PermutationOutput2[60]), 
        .A2(PermutationOutput2[63]), .ZN(SubCellInst2_LFInst_15_LFInst_2_n14)
         );
  INV_X1 SubCellInst2_LFInst_15_LFInst_2_U1 ( .A(PermutationOutput2[62]), .ZN(
        SubCellInst2_LFInst_15_LFInst_2_n15) );
  OR2_X1 SubCellInst2_LFInst_15_LFInst_3_U4 ( .A1(
        SubCellInst2_LFInst_15_LFInst_3_n9), .A2(
        SubCellInst2_LFInst_15_LFInst_3_n8), .ZN(Output[63]) );
  NOR2_X1 SubCellInst2_LFInst_15_LFInst_3_U3 ( .A1(PermutationOutput2[61]), 
        .A2(PermutationOutput2[62]), .ZN(SubCellInst2_LFInst_15_LFInst_3_n8)
         );
  NOR2_X1 SubCellInst2_LFInst_15_LFInst_3_U2 ( .A1(PermutationOutput2[63]), 
        .A2(SubCellInst2_LFInst_15_LFInst_3_n7), .ZN(
        SubCellInst2_LFInst_15_LFInst_3_n9) );
  AND2_X1 SubCellInst2_LFInst_15_LFInst_3_U1 ( .A1(PermutationOutput2[61]), 
        .A2(PermutationOutput2[60]), .ZN(SubCellInst2_LFInst_15_LFInst_3_n7)
         );
  XNOR2_X1 Red_PlaintextInst_LFInst_0_LFInst_0_U3 ( .A(
        Red_PlaintextInst_LFInst_0_LFInst_0_n6), .B(
        Red_PlaintextInst_LFInst_0_LFInst_0_n5), .ZN(Red_MCOutput[0]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_0_LFInst_0_U2 ( .A(Input[2]), .B(Input[3]), 
        .ZN(Red_PlaintextInst_LFInst_0_LFInst_0_n5) );
  XOR2_X1 Red_PlaintextInst_LFInst_0_LFInst_0_U1 ( .A(Input[0]), .B(Input[1]), 
        .Z(Red_PlaintextInst_LFInst_0_LFInst_0_n6) );
  XNOR2_X1 Red_PlaintextInst_LFInst_1_LFInst_0_U3 ( .A(
        Red_PlaintextInst_LFInst_1_LFInst_0_n6), .B(
        Red_PlaintextInst_LFInst_1_LFInst_0_n5), .ZN(Red_MCOutput[1]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_1_LFInst_0_U2 ( .A(Input[6]), .B(Input[7]), 
        .ZN(Red_PlaintextInst_LFInst_1_LFInst_0_n5) );
  XOR2_X1 Red_PlaintextInst_LFInst_1_LFInst_0_U1 ( .A(Input[4]), .B(Input[5]), 
        .Z(Red_PlaintextInst_LFInst_1_LFInst_0_n6) );
  XNOR2_X1 Red_PlaintextInst_LFInst_2_LFInst_0_U3 ( .A(
        Red_PlaintextInst_LFInst_2_LFInst_0_n6), .B(
        Red_PlaintextInst_LFInst_2_LFInst_0_n5), .ZN(Red_MCOutput[2]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_2_LFInst_0_U2 ( .A(Input[10]), .B(
        Input[11]), .ZN(Red_PlaintextInst_LFInst_2_LFInst_0_n5) );
  XOR2_X1 Red_PlaintextInst_LFInst_2_LFInst_0_U1 ( .A(Input[8]), .B(Input[9]), 
        .Z(Red_PlaintextInst_LFInst_2_LFInst_0_n6) );
  XNOR2_X1 Red_PlaintextInst_LFInst_3_LFInst_0_U3 ( .A(
        Red_PlaintextInst_LFInst_3_LFInst_0_n6), .B(
        Red_PlaintextInst_LFInst_3_LFInst_0_n5), .ZN(Red_MCOutput[3]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_3_LFInst_0_U2 ( .A(Input[14]), .B(
        Input[15]), .ZN(Red_PlaintextInst_LFInst_3_LFInst_0_n5) );
  XOR2_X1 Red_PlaintextInst_LFInst_3_LFInst_0_U1 ( .A(Input[12]), .B(Input[13]), .Z(Red_PlaintextInst_LFInst_3_LFInst_0_n6) );
  XNOR2_X1 Red_PlaintextInst_LFInst_4_LFInst_0_U3 ( .A(
        Red_PlaintextInst_LFInst_4_LFInst_0_n6), .B(
        Red_PlaintextInst_LFInst_4_LFInst_0_n5), .ZN(Red_MCOutput[4]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_4_LFInst_0_U2 ( .A(Input[18]), .B(
        Input[19]), .ZN(Red_PlaintextInst_LFInst_4_LFInst_0_n5) );
  XOR2_X1 Red_PlaintextInst_LFInst_4_LFInst_0_U1 ( .A(Input[16]), .B(Input[17]), .Z(Red_PlaintextInst_LFInst_4_LFInst_0_n6) );
  XNOR2_X1 Red_PlaintextInst_LFInst_5_LFInst_0_U3 ( .A(
        Red_PlaintextInst_LFInst_5_LFInst_0_n6), .B(
        Red_PlaintextInst_LFInst_5_LFInst_0_n5), .ZN(Red_MCOutput[5]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_5_LFInst_0_U2 ( .A(Input[22]), .B(
        Input[23]), .ZN(Red_PlaintextInst_LFInst_5_LFInst_0_n5) );
  XOR2_X1 Red_PlaintextInst_LFInst_5_LFInst_0_U1 ( .A(Input[20]), .B(Input[21]), .Z(Red_PlaintextInst_LFInst_5_LFInst_0_n6) );
  XNOR2_X1 Red_PlaintextInst_LFInst_6_LFInst_0_U3 ( .A(
        Red_PlaintextInst_LFInst_6_LFInst_0_n6), .B(
        Red_PlaintextInst_LFInst_6_LFInst_0_n5), .ZN(Red_MCOutput[6]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_6_LFInst_0_U2 ( .A(Input[26]), .B(
        Input[27]), .ZN(Red_PlaintextInst_LFInst_6_LFInst_0_n5) );
  XOR2_X1 Red_PlaintextInst_LFInst_6_LFInst_0_U1 ( .A(Input[24]), .B(Input[25]), .Z(Red_PlaintextInst_LFInst_6_LFInst_0_n6) );
  XNOR2_X1 Red_PlaintextInst_LFInst_7_LFInst_0_U3 ( .A(
        Red_PlaintextInst_LFInst_7_LFInst_0_n6), .B(
        Red_PlaintextInst_LFInst_7_LFInst_0_n5), .ZN(Red_MCOutput[7]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_7_LFInst_0_U2 ( .A(Input[30]), .B(
        Input[31]), .ZN(Red_PlaintextInst_LFInst_7_LFInst_0_n5) );
  XOR2_X1 Red_PlaintextInst_LFInst_7_LFInst_0_U1 ( .A(Input[28]), .B(Input[29]), .Z(Red_PlaintextInst_LFInst_7_LFInst_0_n6) );
  XNOR2_X1 Red_PlaintextInst_LFInst_8_LFInst_0_U3 ( .A(
        Red_PlaintextInst_LFInst_8_LFInst_0_n6), .B(
        Red_PlaintextInst_LFInst_8_LFInst_0_n5), .ZN(Red_Input[8]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_8_LFInst_0_U2 ( .A(Input[34]), .B(
        Input[35]), .ZN(Red_PlaintextInst_LFInst_8_LFInst_0_n5) );
  XOR2_X1 Red_PlaintextInst_LFInst_8_LFInst_0_U1 ( .A(Input[32]), .B(Input[33]), .Z(Red_PlaintextInst_LFInst_8_LFInst_0_n6) );
  XNOR2_X1 Red_PlaintextInst_LFInst_9_LFInst_0_U3 ( .A(
        Red_PlaintextInst_LFInst_9_LFInst_0_n6), .B(
        Red_PlaintextInst_LFInst_9_LFInst_0_n5), .ZN(Red_Input[9]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_9_LFInst_0_U2 ( .A(Input[38]), .B(
        Input[39]), .ZN(Red_PlaintextInst_LFInst_9_LFInst_0_n5) );
  XOR2_X1 Red_PlaintextInst_LFInst_9_LFInst_0_U1 ( .A(Input[36]), .B(Input[37]), .Z(Red_PlaintextInst_LFInst_9_LFInst_0_n6) );
  XNOR2_X1 Red_PlaintextInst_LFInst_10_LFInst_0_U3 ( .A(
        Red_PlaintextInst_LFInst_10_LFInst_0_n6), .B(
        Red_PlaintextInst_LFInst_10_LFInst_0_n5), .ZN(Red_Input[10]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_10_LFInst_0_U2 ( .A(Input[42]), .B(
        Input[43]), .ZN(Red_PlaintextInst_LFInst_10_LFInst_0_n5) );
  XOR2_X1 Red_PlaintextInst_LFInst_10_LFInst_0_U1 ( .A(Input[40]), .B(
        Input[41]), .Z(Red_PlaintextInst_LFInst_10_LFInst_0_n6) );
  XNOR2_X1 Red_PlaintextInst_LFInst_11_LFInst_0_U3 ( .A(
        Red_PlaintextInst_LFInst_11_LFInst_0_n6), .B(
        Red_PlaintextInst_LFInst_11_LFInst_0_n5), .ZN(Red_Input[11]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_11_LFInst_0_U2 ( .A(Input[46]), .B(
        Input[47]), .ZN(Red_PlaintextInst_LFInst_11_LFInst_0_n5) );
  XOR2_X1 Red_PlaintextInst_LFInst_11_LFInst_0_U1 ( .A(Input[44]), .B(
        Input[45]), .Z(Red_PlaintextInst_LFInst_11_LFInst_0_n6) );
  XNOR2_X1 Red_PlaintextInst_LFInst_12_LFInst_0_U3 ( .A(
        Red_PlaintextInst_LFInst_12_LFInst_0_n6), .B(
        Red_PlaintextInst_LFInst_12_LFInst_0_n5), .ZN(Red_Input[12]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_12_LFInst_0_U2 ( .A(Input[50]), .B(
        Input[51]), .ZN(Red_PlaintextInst_LFInst_12_LFInst_0_n5) );
  XOR2_X1 Red_PlaintextInst_LFInst_12_LFInst_0_U1 ( .A(Input[48]), .B(
        Input[49]), .Z(Red_PlaintextInst_LFInst_12_LFInst_0_n6) );
  XNOR2_X1 Red_PlaintextInst_LFInst_13_LFInst_0_U3 ( .A(
        Red_PlaintextInst_LFInst_13_LFInst_0_n6), .B(
        Red_PlaintextInst_LFInst_13_LFInst_0_n5), .ZN(Red_Input[13]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_13_LFInst_0_U2 ( .A(Input[54]), .B(
        Input[55]), .ZN(Red_PlaintextInst_LFInst_13_LFInst_0_n5) );
  XOR2_X1 Red_PlaintextInst_LFInst_13_LFInst_0_U1 ( .A(Input[52]), .B(
        Input[53]), .Z(Red_PlaintextInst_LFInst_13_LFInst_0_n6) );
  XNOR2_X1 Red_PlaintextInst_LFInst_14_LFInst_0_U3 ( .A(
        Red_PlaintextInst_LFInst_14_LFInst_0_n6), .B(
        Red_PlaintextInst_LFInst_14_LFInst_0_n5), .ZN(Red_Input[14]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_14_LFInst_0_U2 ( .A(Input[58]), .B(
        Input[59]), .ZN(Red_PlaintextInst_LFInst_14_LFInst_0_n5) );
  XOR2_X1 Red_PlaintextInst_LFInst_14_LFInst_0_U1 ( .A(Input[56]), .B(
        Input[57]), .Z(Red_PlaintextInst_LFInst_14_LFInst_0_n6) );
  XNOR2_X1 Red_PlaintextInst_LFInst_15_LFInst_0_U3 ( .A(
        Red_PlaintextInst_LFInst_15_LFInst_0_n6), .B(
        Red_PlaintextInst_LFInst_15_LFInst_0_n5), .ZN(Red_Input[15]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_15_LFInst_0_U2 ( .A(Input[62]), .B(
        Input[63]), .ZN(Red_PlaintextInst_LFInst_15_LFInst_0_n5) );
  XOR2_X1 Red_PlaintextInst_LFInst_15_LFInst_0_U1 ( .A(Input[60]), .B(
        Input[61]), .Z(Red_PlaintextInst_LFInst_15_LFInst_0_n6) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_0_U2 ( .A(Red_MCInst_XOR_r0_Inst_0_n5), .B(
        Red_MCOutput[4]), .ZN(Red_MCOutput[12]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_0_U1 ( .A(Red_MCOutput[0]), .B(Red_Input[12]), .ZN(Red_MCInst_XOR_r0_Inst_0_n5) );
  XOR2_X1 Red_MCInst_XOR_r1_Inst_0_U1 ( .A(Red_Input[8]), .B(Red_MCOutput[0]), 
        .Z(Red_MCOutput[8]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_1_U2 ( .A(Red_MCInst_XOR_r0_Inst_1_n5), .B(
        Red_MCOutput[5]), .ZN(Red_MCOutput[13]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_1_U1 ( .A(Red_MCOutput[1]), .B(Red_Input[13]), .ZN(Red_MCInst_XOR_r0_Inst_1_n5) );
  XOR2_X1 Red_MCInst_XOR_r1_Inst_1_U1 ( .A(Red_Input[9]), .B(Red_MCOutput[1]), 
        .Z(Red_MCOutput[9]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_2_U2 ( .A(Red_MCInst_XOR_r0_Inst_2_n5), .B(
        Red_MCOutput[6]), .ZN(Red_MCOutput[14]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_2_U1 ( .A(Red_MCOutput[2]), .B(Red_Input[14]), .ZN(Red_MCInst_XOR_r0_Inst_2_n5) );
  XOR2_X1 Red_MCInst_XOR_r1_Inst_2_U1 ( .A(Red_Input[10]), .B(Red_MCOutput[2]), 
        .Z(Red_MCOutput[10]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_3_U2 ( .A(Red_MCInst_XOR_r0_Inst_3_n5), .B(
        Red_MCOutput[7]), .ZN(Red_MCOutput[15]) );
  XNOR2_X1 Red_MCInst_XOR_r0_Inst_3_U1 ( .A(Red_MCOutput[3]), .B(Red_Input[15]), .ZN(Red_MCInst_XOR_r0_Inst_3_n5) );
  XOR2_X1 Red_MCInst_XOR_r1_Inst_3_U1 ( .A(Red_Input[11]), .B(Red_MCOutput[3]), 
        .Z(Red_MCOutput[11]) );
  XOR2_X1 Red_AddKeyXOR1_XORInst_0_0_U1 ( .A(Red_MCOutput[12]), .B(Red_K0[12]), 
        .Z(Red_final[28]) );
  XOR2_X1 Red_AddKeyXOR1_XORInst_1_0_U1 ( .A(Red_MCOutput[13]), .B(Red_K0[13]), 
        .Z(Red_final[29]) );
  XOR2_X1 Red_AddKeyXOR1_XORInst_2_0_U1 ( .A(Red_MCOutput[14]), .B(Red_K0[14]), 
        .Z(Red_final[30]) );
  XOR2_X1 Red_AddKeyXOR1_XORInst_3_0_U1 ( .A(Red_MCOutput[15]), .B(Red_K0[15]), 
        .Z(Red_final[31]) );
  XOR2_X1 Red_AddKeyConstXOR_XORInst_0_0_U1 ( .A(Red_MCOutput[10]), .B(
        Red_K0[10]), .Z(Red_final[26]) );
  XOR2_X1 Red_AddKeyConstXOR_XORInst_1_0_U1 ( .A(Red_MCOutput[11]), .B(
        Red_K0[11]), .Z(Red_final[27]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_0_0_U1 ( .A(Red_MCOutput[0]), .B(Red_K0[0]), 
        .Z(Red_final[16]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_1_0_U1 ( .A(Red_MCOutput[1]), .B(Red_K0[1]), 
        .Z(Red_final[17]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_2_0_U1 ( .A(Red_MCOutput[2]), .B(Red_K0[2]), 
        .Z(Red_final[18]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_3_0_U1 ( .A(Red_MCOutput[3]), .B(Red_K0[3]), 
        .Z(Red_final[19]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_4_0_U1 ( .A(Red_MCOutput[4]), .B(Red_K0[4]), 
        .Z(Red_final[20]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_5_0_U1 ( .A(Red_MCOutput[5]), .B(Red_K0[5]), 
        .Z(Red_final[21]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_6_0_U1 ( .A(Red_MCOutput[6]), .B(Red_K0[6]), 
        .Z(Red_final[22]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_7_0_U1 ( .A(Red_MCOutput[7]), .B(Red_K0[7]), 
        .Z(Red_final[23]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_8_0_U1 ( .A(Red_MCOutput[8]), .B(Red_K0[8]), 
        .Z(Red_final[24]) );
  XOR2_X1 Red_AddKeyXOR2_XORInst_9_0_U1 ( .A(Red_MCOutput[9]), .B(Red_K0[9]), 
        .Z(Red_final[25]) );
  DFF_X1 Red_StateReg_s_current_state_reg_0_ ( .D(Red_final[16]), .CK(clk), 
        .Q(Red_StateRegOutput[0]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_1_ ( .D(Red_final[17]), .CK(clk), 
        .Q(Red_StateRegOutput[1]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_2_ ( .D(Red_final[18]), .CK(clk), 
        .Q(Red_StateRegOutput[2]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_3_ ( .D(Red_final[19]), .CK(clk), 
        .Q(Red_StateRegOutput[3]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_4_ ( .D(Red_final[20]), .CK(clk), 
        .Q(Red_StateRegOutput[4]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_5_ ( .D(Red_final[21]), .CK(clk), 
        .Q(Red_StateRegOutput[5]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_6_ ( .D(Red_final[22]), .CK(clk), 
        .Q(Red_StateRegOutput[6]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_7_ ( .D(Red_final[23]), .CK(clk), 
        .Q(Red_StateRegOutput[7]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_8_ ( .D(Red_final[24]), .CK(clk), 
        .Q(Red_StateRegOutput[8]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_9_ ( .D(Red_final[25]), .CK(clk), 
        .Q(Red_StateRegOutput[9]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_10_ ( .D(Red_final[26]), .CK(clk), 
        .Q(Red_StateRegOutput[10]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_11_ ( .D(Red_final[27]), .CK(clk), 
        .Q(Red_StateRegOutput[11]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_12_ ( .D(Red_final[28]), .CK(clk), 
        .Q(Red_StateRegOutput[12]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_13_ ( .D(Red_final[29]), .CK(clk), 
        .Q(Red_StateRegOutput[13]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_14_ ( .D(Red_final[30]), .CK(clk), 
        .Q(Red_StateRegOutput[14]), .QN() );
  DFF_X1 Red_StateReg_s_current_state_reg_15_ ( .D(Red_final[31]), .CK(clk), 
        .Q(Red_StateRegOutput[15]), .QN() );
  NAND2_X1 Red_SubCellInst_LFInst_0_LFInst_0_U10 ( .A1(
        Red_SubCellInst_LFInst_0_LFInst_0_n20), .A2(
        Red_SubCellInst_LFInst_0_LFInst_0_n19), .ZN(
        Red_SubCellInst_LFInst_0_LFInst_0_n21) );
  INV_X1 Red_SubCellInst_LFInst_0_LFInst_0_U9 ( .A(PermutationOutput[2]), .ZN(
        Red_SubCellInst_LFInst_0_LFInst_0_n19) );
  NAND2_X1 Red_SubCellInst_LFInst_0_LFInst_0_U8 ( .A1(
        Red_SubCellInst_LFInst_0_LFInst_0_n18), .A2(PermutationOutput[2]), 
        .ZN(Red_SubCellInst_LFInst_0_LFInst_0_n22) );
  XNOR2_X1 Red_SubCellInst_LFInst_0_LFInst_0_U7 ( .A(
        Red_SubCellInst_LFInst_0_LFInst_0_n17), .B(
        Red_SubCellInst_LFInst_0_LFInst_0_n20), .ZN(
        Red_SubCellInst_LFInst_0_LFInst_0_n18) );
  NOR2_X1 Red_SubCellInst_LFInst_0_LFInst_0_U6 ( .A1(
        Red_SubCellInst_LFInst_0_LFInst_0_n16), .A2(
        Red_SubCellInst_LFInst_0_LFInst_0_n15), .ZN(
        Red_SubCellInst_LFInst_0_LFInst_0_n17) );
  INV_X1 Red_SubCellInst_LFInst_0_LFInst_0_U5 ( .A(PermutationOutput[1]), .ZN(
        Red_SubCellInst_LFInst_0_LFInst_0_n15) );
  INV_X1 Red_SubCellInst_LFInst_0_LFInst_0_U4 ( .A(PermutationOutput[3]), .ZN(
        Red_SubCellInst_LFInst_0_LFInst_0_n16) );
  AND2_X1 Red_SubCellInst_LFInst_0_LFInst_0_U3 ( .A1(
        Red_SubCellInst_LFInst_0_LFInst_0_n22), .A2(
        Red_SubCellInst_LFInst_0_LFInst_0_n21), .ZN(Red_MCOutput2[0]) );
  OR2_X1 Red_SubCellInst_LFInst_0_LFInst_0_U2 ( .A1(
        Red_SubCellInst_LFInst_0_LFInst_0_n14), .A2(PermutationOutput[0]), 
        .ZN(Red_SubCellInst_LFInst_0_LFInst_0_n20) );
  AND2_X1 Red_SubCellInst_LFInst_0_LFInst_0_U1 ( .A1(
        Red_SubCellInst_LFInst_0_LFInst_0_n15), .A2(
        Red_SubCellInst_LFInst_0_LFInst_0_n16), .ZN(
        Red_SubCellInst_LFInst_0_LFInst_0_n14) );
  NAND2_X1 Red_SubCellInst_LFInst_1_LFInst_0_U10 ( .A1(
        Red_SubCellInst_LFInst_1_LFInst_0_n20), .A2(
        Red_SubCellInst_LFInst_1_LFInst_0_n19), .ZN(
        Red_SubCellInst_LFInst_1_LFInst_0_n21) );
  INV_X1 Red_SubCellInst_LFInst_1_LFInst_0_U9 ( .A(PermutationOutput[6]), .ZN(
        Red_SubCellInst_LFInst_1_LFInst_0_n19) );
  NAND2_X1 Red_SubCellInst_LFInst_1_LFInst_0_U8 ( .A1(
        Red_SubCellInst_LFInst_1_LFInst_0_n18), .A2(PermutationOutput[6]), 
        .ZN(Red_SubCellInst_LFInst_1_LFInst_0_n22) );
  XNOR2_X1 Red_SubCellInst_LFInst_1_LFInst_0_U7 ( .A(
        Red_SubCellInst_LFInst_1_LFInst_0_n17), .B(
        Red_SubCellInst_LFInst_1_LFInst_0_n20), .ZN(
        Red_SubCellInst_LFInst_1_LFInst_0_n18) );
  NOR2_X1 Red_SubCellInst_LFInst_1_LFInst_0_U6 ( .A1(
        Red_SubCellInst_LFInst_1_LFInst_0_n16), .A2(
        Red_SubCellInst_LFInst_1_LFInst_0_n15), .ZN(
        Red_SubCellInst_LFInst_1_LFInst_0_n17) );
  INV_X1 Red_SubCellInst_LFInst_1_LFInst_0_U5 ( .A(PermutationOutput[5]), .ZN(
        Red_SubCellInst_LFInst_1_LFInst_0_n15) );
  INV_X1 Red_SubCellInst_LFInst_1_LFInst_0_U4 ( .A(PermutationOutput[7]), .ZN(
        Red_SubCellInst_LFInst_1_LFInst_0_n16) );
  AND2_X1 Red_SubCellInst_LFInst_1_LFInst_0_U3 ( .A1(
        Red_SubCellInst_LFInst_1_LFInst_0_n22), .A2(
        Red_SubCellInst_LFInst_1_LFInst_0_n21), .ZN(Red_MCOutput2[1]) );
  OR2_X1 Red_SubCellInst_LFInst_1_LFInst_0_U2 ( .A1(
        Red_SubCellInst_LFInst_1_LFInst_0_n14), .A2(PermutationOutput[4]), 
        .ZN(Red_SubCellInst_LFInst_1_LFInst_0_n20) );
  AND2_X1 Red_SubCellInst_LFInst_1_LFInst_0_U1 ( .A1(
        Red_SubCellInst_LFInst_1_LFInst_0_n15), .A2(
        Red_SubCellInst_LFInst_1_LFInst_0_n16), .ZN(
        Red_SubCellInst_LFInst_1_LFInst_0_n14) );
  NAND2_X1 Red_SubCellInst_LFInst_2_LFInst_0_U10 ( .A1(
        Red_SubCellInst_LFInst_2_LFInst_0_n20), .A2(
        Red_SubCellInst_LFInst_2_LFInst_0_n19), .ZN(
        Red_SubCellInst_LFInst_2_LFInst_0_n21) );
  INV_X1 Red_SubCellInst_LFInst_2_LFInst_0_U9 ( .A(PermutationOutput[10]), 
        .ZN(Red_SubCellInst_LFInst_2_LFInst_0_n19) );
  NAND2_X1 Red_SubCellInst_LFInst_2_LFInst_0_U8 ( .A1(
        Red_SubCellInst_LFInst_2_LFInst_0_n18), .A2(PermutationOutput[10]), 
        .ZN(Red_SubCellInst_LFInst_2_LFInst_0_n22) );
  XNOR2_X1 Red_SubCellInst_LFInst_2_LFInst_0_U7 ( .A(
        Red_SubCellInst_LFInst_2_LFInst_0_n17), .B(
        Red_SubCellInst_LFInst_2_LFInst_0_n20), .ZN(
        Red_SubCellInst_LFInst_2_LFInst_0_n18) );
  NOR2_X1 Red_SubCellInst_LFInst_2_LFInst_0_U6 ( .A1(
        Red_SubCellInst_LFInst_2_LFInst_0_n16), .A2(
        Red_SubCellInst_LFInst_2_LFInst_0_n15), .ZN(
        Red_SubCellInst_LFInst_2_LFInst_0_n17) );
  INV_X1 Red_SubCellInst_LFInst_2_LFInst_0_U5 ( .A(PermutationOutput[9]), .ZN(
        Red_SubCellInst_LFInst_2_LFInst_0_n15) );
  INV_X1 Red_SubCellInst_LFInst_2_LFInst_0_U4 ( .A(PermutationOutput[11]), 
        .ZN(Red_SubCellInst_LFInst_2_LFInst_0_n16) );
  AND2_X1 Red_SubCellInst_LFInst_2_LFInst_0_U3 ( .A1(
        Red_SubCellInst_LFInst_2_LFInst_0_n22), .A2(
        Red_SubCellInst_LFInst_2_LFInst_0_n21), .ZN(Red_MCOutput2[2]) );
  OR2_X1 Red_SubCellInst_LFInst_2_LFInst_0_U2 ( .A1(
        Red_SubCellInst_LFInst_2_LFInst_0_n14), .A2(PermutationOutput[8]), 
        .ZN(Red_SubCellInst_LFInst_2_LFInst_0_n20) );
  AND2_X1 Red_SubCellInst_LFInst_2_LFInst_0_U1 ( .A1(
        Red_SubCellInst_LFInst_2_LFInst_0_n15), .A2(
        Red_SubCellInst_LFInst_2_LFInst_0_n16), .ZN(
        Red_SubCellInst_LFInst_2_LFInst_0_n14) );
  NAND2_X1 Red_SubCellInst_LFInst_3_LFInst_0_U10 ( .A1(
        Red_SubCellInst_LFInst_3_LFInst_0_n20), .A2(
        Red_SubCellInst_LFInst_3_LFInst_0_n19), .ZN(
        Red_SubCellInst_LFInst_3_LFInst_0_n21) );
  INV_X1 Red_SubCellInst_LFInst_3_LFInst_0_U9 ( .A(PermutationOutput[14]), 
        .ZN(Red_SubCellInst_LFInst_3_LFInst_0_n19) );
  NAND2_X1 Red_SubCellInst_LFInst_3_LFInst_0_U8 ( .A1(
        Red_SubCellInst_LFInst_3_LFInst_0_n18), .A2(PermutationOutput[14]), 
        .ZN(Red_SubCellInst_LFInst_3_LFInst_0_n22) );
  XNOR2_X1 Red_SubCellInst_LFInst_3_LFInst_0_U7 ( .A(
        Red_SubCellInst_LFInst_3_LFInst_0_n17), .B(
        Red_SubCellInst_LFInst_3_LFInst_0_n20), .ZN(
        Red_SubCellInst_LFInst_3_LFInst_0_n18) );
  NOR2_X1 Red_SubCellInst_LFInst_3_LFInst_0_U6 ( .A1(
        Red_SubCellInst_LFInst_3_LFInst_0_n16), .A2(
        Red_SubCellInst_LFInst_3_LFInst_0_n15), .ZN(
        Red_SubCellInst_LFInst_3_LFInst_0_n17) );
  INV_X1 Red_SubCellInst_LFInst_3_LFInst_0_U5 ( .A(PermutationOutput[13]), 
        .ZN(Red_SubCellInst_LFInst_3_LFInst_0_n15) );
  INV_X1 Red_SubCellInst_LFInst_3_LFInst_0_U4 ( .A(PermutationOutput[15]), 
        .ZN(Red_SubCellInst_LFInst_3_LFInst_0_n16) );
  AND2_X1 Red_SubCellInst_LFInst_3_LFInst_0_U3 ( .A1(
        Red_SubCellInst_LFInst_3_LFInst_0_n22), .A2(
        Red_SubCellInst_LFInst_3_LFInst_0_n21), .ZN(Red_MCOutput2[3]) );
  OR2_X1 Red_SubCellInst_LFInst_3_LFInst_0_U2 ( .A1(
        Red_SubCellInst_LFInst_3_LFInst_0_n14), .A2(PermutationOutput[12]), 
        .ZN(Red_SubCellInst_LFInst_3_LFInst_0_n20) );
  AND2_X1 Red_SubCellInst_LFInst_3_LFInst_0_U1 ( .A1(
        Red_SubCellInst_LFInst_3_LFInst_0_n15), .A2(
        Red_SubCellInst_LFInst_3_LFInst_0_n16), .ZN(
        Red_SubCellInst_LFInst_3_LFInst_0_n14) );
  INV_X1 Red_SubCellInst_LFInst_4_LFInst_0_U7 ( .A(PermutationOutput[17]), 
        .ZN(Red_SubCellInst_LFInst_4_LFInst_0_n18) );
  INV_X1 Red_SubCellInst_LFInst_4_LFInst_0_U6 ( .A(PermutationOutput[19]), 
        .ZN(Red_SubCellInst_LFInst_4_LFInst_0_n19) );
  XNOR2_X1 Red_SubCellInst_LFInst_4_LFInst_0_U5 ( .A(
        Red_SubCellInst_LFInst_4_LFInst_0_n15), .B(
        Red_SubCellInst_LFInst_4_LFInst_0_n17), .ZN(Red_MCOutput2[4]) );
  NOR2_X1 Red_SubCellInst_LFInst_4_LFInst_0_U4 ( .A1(
        Red_SubCellInst_LFInst_4_LFInst_0_n16), .A2(PermutationOutput[16]), 
        .ZN(Red_SubCellInst_LFInst_4_LFInst_0_n17) );
  AND2_X1 Red_SubCellInst_LFInst_4_LFInst_0_U3 ( .A1(
        Red_SubCellInst_LFInst_4_LFInst_0_n19), .A2(
        Red_SubCellInst_LFInst_4_LFInst_0_n18), .ZN(
        Red_SubCellInst_LFInst_4_LFInst_0_n16) );
  NAND2_X1 Red_SubCellInst_LFInst_4_LFInst_0_U2 ( .A1(
        Red_SubCellInst_LFInst_4_LFInst_0_n14), .A2(PermutationOutput[18]), 
        .ZN(Red_SubCellInst_LFInst_4_LFInst_0_n15) );
  OR2_X1 Red_SubCellInst_LFInst_4_LFInst_0_U1 ( .A1(
        Red_SubCellInst_LFInst_4_LFInst_0_n19), .A2(
        Red_SubCellInst_LFInst_4_LFInst_0_n18), .ZN(
        Red_SubCellInst_LFInst_4_LFInst_0_n14) );
  INV_X1 Red_SubCellInst_LFInst_5_LFInst_0_U7 ( .A(PermutationOutput[21]), 
        .ZN(Red_SubCellInst_LFInst_5_LFInst_0_n18) );
  INV_X1 Red_SubCellInst_LFInst_5_LFInst_0_U6 ( .A(PermutationOutput[23]), 
        .ZN(Red_SubCellInst_LFInst_5_LFInst_0_n19) );
  XNOR2_X1 Red_SubCellInst_LFInst_5_LFInst_0_U5 ( .A(
        Red_SubCellInst_LFInst_5_LFInst_0_n15), .B(
        Red_SubCellInst_LFInst_5_LFInst_0_n17), .ZN(Red_MCOutput2[5]) );
  NOR2_X1 Red_SubCellInst_LFInst_5_LFInst_0_U4 ( .A1(
        Red_SubCellInst_LFInst_5_LFInst_0_n16), .A2(PermutationOutput[20]), 
        .ZN(Red_SubCellInst_LFInst_5_LFInst_0_n17) );
  AND2_X1 Red_SubCellInst_LFInst_5_LFInst_0_U3 ( .A1(
        Red_SubCellInst_LFInst_5_LFInst_0_n19), .A2(
        Red_SubCellInst_LFInst_5_LFInst_0_n18), .ZN(
        Red_SubCellInst_LFInst_5_LFInst_0_n16) );
  NAND2_X1 Red_SubCellInst_LFInst_5_LFInst_0_U2 ( .A1(
        Red_SubCellInst_LFInst_5_LFInst_0_n14), .A2(PermutationOutput[22]), 
        .ZN(Red_SubCellInst_LFInst_5_LFInst_0_n15) );
  OR2_X1 Red_SubCellInst_LFInst_5_LFInst_0_U1 ( .A1(
        Red_SubCellInst_LFInst_5_LFInst_0_n19), .A2(
        Red_SubCellInst_LFInst_5_LFInst_0_n18), .ZN(
        Red_SubCellInst_LFInst_5_LFInst_0_n14) );
  INV_X1 Red_SubCellInst_LFInst_6_LFInst_0_U7 ( .A(PermutationOutput[25]), 
        .ZN(Red_SubCellInst_LFInst_6_LFInst_0_n18) );
  INV_X1 Red_SubCellInst_LFInst_6_LFInst_0_U6 ( .A(PermutationOutput[27]), 
        .ZN(Red_SubCellInst_LFInst_6_LFInst_0_n19) );
  XNOR2_X1 Red_SubCellInst_LFInst_6_LFInst_0_U5 ( .A(
        Red_SubCellInst_LFInst_6_LFInst_0_n15), .B(
        Red_SubCellInst_LFInst_6_LFInst_0_n17), .ZN(Red_MCOutput2[6]) );
  NOR2_X1 Red_SubCellInst_LFInst_6_LFInst_0_U4 ( .A1(
        Red_SubCellInst_LFInst_6_LFInst_0_n16), .A2(PermutationOutput[24]), 
        .ZN(Red_SubCellInst_LFInst_6_LFInst_0_n17) );
  AND2_X1 Red_SubCellInst_LFInst_6_LFInst_0_U3 ( .A1(
        Red_SubCellInst_LFInst_6_LFInst_0_n19), .A2(
        Red_SubCellInst_LFInst_6_LFInst_0_n18), .ZN(
        Red_SubCellInst_LFInst_6_LFInst_0_n16) );
  NAND2_X1 Red_SubCellInst_LFInst_6_LFInst_0_U2 ( .A1(
        Red_SubCellInst_LFInst_6_LFInst_0_n14), .A2(PermutationOutput[26]), 
        .ZN(Red_SubCellInst_LFInst_6_LFInst_0_n15) );
  OR2_X1 Red_SubCellInst_LFInst_6_LFInst_0_U1 ( .A1(
        Red_SubCellInst_LFInst_6_LFInst_0_n19), .A2(
        Red_SubCellInst_LFInst_6_LFInst_0_n18), .ZN(
        Red_SubCellInst_LFInst_6_LFInst_0_n14) );
  INV_X1 Red_SubCellInst_LFInst_7_LFInst_0_U7 ( .A(PermutationOutput[29]), 
        .ZN(Red_SubCellInst_LFInst_7_LFInst_0_n18) );
  INV_X1 Red_SubCellInst_LFInst_7_LFInst_0_U6 ( .A(PermutationOutput[31]), 
        .ZN(Red_SubCellInst_LFInst_7_LFInst_0_n19) );
  XNOR2_X1 Red_SubCellInst_LFInst_7_LFInst_0_U5 ( .A(
        Red_SubCellInst_LFInst_7_LFInst_0_n17), .B(
        Red_SubCellInst_LFInst_7_LFInst_0_n16), .ZN(Red_MCOutput2[7]) );
  NAND2_X1 Red_SubCellInst_LFInst_7_LFInst_0_U4 ( .A1(
        Red_SubCellInst_LFInst_7_LFInst_0_n14), .A2(PermutationOutput[30]), 
        .ZN(Red_SubCellInst_LFInst_7_LFInst_0_n17) );
  NOR2_X1 Red_SubCellInst_LFInst_7_LFInst_0_U3 ( .A1(
        Red_SubCellInst_LFInst_7_LFInst_0_n15), .A2(PermutationOutput[28]), 
        .ZN(Red_SubCellInst_LFInst_7_LFInst_0_n16) );
  AND2_X1 Red_SubCellInst_LFInst_7_LFInst_0_U2 ( .A1(
        Red_SubCellInst_LFInst_7_LFInst_0_n19), .A2(
        Red_SubCellInst_LFInst_7_LFInst_0_n18), .ZN(
        Red_SubCellInst_LFInst_7_LFInst_0_n15) );
  OR2_X1 Red_SubCellInst_LFInst_7_LFInst_0_U1 ( .A1(
        Red_SubCellInst_LFInst_7_LFInst_0_n19), .A2(
        Red_SubCellInst_LFInst_7_LFInst_0_n18), .ZN(
        Red_SubCellInst_LFInst_7_LFInst_0_n14) );
  AND2_X1 Red_SubCellInst_LFInst_8_LFInst_0_U10 ( .A1(
        Red_SubCellInst_LFInst_8_LFInst_0_n22), .A2(
        Red_SubCellInst_LFInst_8_LFInst_0_n21), .ZN(Red_SboxOut[8]) );
  NAND2_X1 Red_SubCellInst_LFInst_8_LFInst_0_U9 ( .A1(
        Red_SubCellInst_LFInst_8_LFInst_0_n20), .A2(
        Red_SubCellInst_LFInst_8_LFInst_0_n19), .ZN(
        Red_SubCellInst_LFInst_8_LFInst_0_n21) );
  INV_X1 Red_SubCellInst_LFInst_8_LFInst_0_U8 ( .A(PermutationOutput[34]), 
        .ZN(Red_SubCellInst_LFInst_8_LFInst_0_n19) );
  NAND2_X1 Red_SubCellInst_LFInst_8_LFInst_0_U7 ( .A1(
        Red_SubCellInst_LFInst_8_LFInst_0_n18), .A2(PermutationOutput[34]), 
        .ZN(Red_SubCellInst_LFInst_8_LFInst_0_n22) );
  XNOR2_X1 Red_SubCellInst_LFInst_8_LFInst_0_U6 ( .A(
        Red_SubCellInst_LFInst_8_LFInst_0_n17), .B(
        Red_SubCellInst_LFInst_8_LFInst_0_n20), .ZN(
        Red_SubCellInst_LFInst_8_LFInst_0_n18) );
  NOR2_X1 Red_SubCellInst_LFInst_8_LFInst_0_U5 ( .A1(
        Red_SubCellInst_LFInst_8_LFInst_0_n16), .A2(
        Red_SubCellInst_LFInst_8_LFInst_0_n15), .ZN(
        Red_SubCellInst_LFInst_8_LFInst_0_n17) );
  INV_X1 Red_SubCellInst_LFInst_8_LFInst_0_U4 ( .A(PermutationOutput[33]), 
        .ZN(Red_SubCellInst_LFInst_8_LFInst_0_n15) );
  INV_X1 Red_SubCellInst_LFInst_8_LFInst_0_U3 ( .A(PermutationOutput[35]), 
        .ZN(Red_SubCellInst_LFInst_8_LFInst_0_n16) );
  OR2_X1 Red_SubCellInst_LFInst_8_LFInst_0_U2 ( .A1(
        Red_SubCellInst_LFInst_8_LFInst_0_n14), .A2(PermutationOutput[32]), 
        .ZN(Red_SubCellInst_LFInst_8_LFInst_0_n20) );
  AND2_X1 Red_SubCellInst_LFInst_8_LFInst_0_U1 ( .A1(
        Red_SubCellInst_LFInst_8_LFInst_0_n15), .A2(
        Red_SubCellInst_LFInst_8_LFInst_0_n16), .ZN(
        Red_SubCellInst_LFInst_8_LFInst_0_n14) );
  AND2_X1 Red_SubCellInst_LFInst_9_LFInst_0_U10 ( .A1(
        Red_SubCellInst_LFInst_9_LFInst_0_n22), .A2(
        Red_SubCellInst_LFInst_9_LFInst_0_n21), .ZN(Red_SboxOut[9]) );
  NAND2_X1 Red_SubCellInst_LFInst_9_LFInst_0_U9 ( .A1(
        Red_SubCellInst_LFInst_9_LFInst_0_n20), .A2(
        Red_SubCellInst_LFInst_9_LFInst_0_n19), .ZN(
        Red_SubCellInst_LFInst_9_LFInst_0_n21) );
  INV_X1 Red_SubCellInst_LFInst_9_LFInst_0_U8 ( .A(PermutationOutput[38]), 
        .ZN(Red_SubCellInst_LFInst_9_LFInst_0_n19) );
  NAND2_X1 Red_SubCellInst_LFInst_9_LFInst_0_U7 ( .A1(
        Red_SubCellInst_LFInst_9_LFInst_0_n18), .A2(PermutationOutput[38]), 
        .ZN(Red_SubCellInst_LFInst_9_LFInst_0_n22) );
  XNOR2_X1 Red_SubCellInst_LFInst_9_LFInst_0_U6 ( .A(
        Red_SubCellInst_LFInst_9_LFInst_0_n17), .B(
        Red_SubCellInst_LFInst_9_LFInst_0_n20), .ZN(
        Red_SubCellInst_LFInst_9_LFInst_0_n18) );
  NOR2_X1 Red_SubCellInst_LFInst_9_LFInst_0_U5 ( .A1(
        Red_SubCellInst_LFInst_9_LFInst_0_n16), .A2(
        Red_SubCellInst_LFInst_9_LFInst_0_n15), .ZN(
        Red_SubCellInst_LFInst_9_LFInst_0_n17) );
  INV_X1 Red_SubCellInst_LFInst_9_LFInst_0_U4 ( .A(PermutationOutput[37]), 
        .ZN(Red_SubCellInst_LFInst_9_LFInst_0_n15) );
  INV_X1 Red_SubCellInst_LFInst_9_LFInst_0_U3 ( .A(PermutationOutput[39]), 
        .ZN(Red_SubCellInst_LFInst_9_LFInst_0_n16) );
  OR2_X1 Red_SubCellInst_LFInst_9_LFInst_0_U2 ( .A1(
        Red_SubCellInst_LFInst_9_LFInst_0_n14), .A2(PermutationOutput[36]), 
        .ZN(Red_SubCellInst_LFInst_9_LFInst_0_n20) );
  AND2_X1 Red_SubCellInst_LFInst_9_LFInst_0_U1 ( .A1(
        Red_SubCellInst_LFInst_9_LFInst_0_n15), .A2(
        Red_SubCellInst_LFInst_9_LFInst_0_n16), .ZN(
        Red_SubCellInst_LFInst_9_LFInst_0_n14) );
  AND2_X1 Red_SubCellInst_LFInst_10_LFInst_0_U10 ( .A1(
        Red_SubCellInst_LFInst_10_LFInst_0_n22), .A2(
        Red_SubCellInst_LFInst_10_LFInst_0_n21), .ZN(Red_SboxOut[10]) );
  NAND2_X1 Red_SubCellInst_LFInst_10_LFInst_0_U9 ( .A1(
        Red_SubCellInst_LFInst_10_LFInst_0_n20), .A2(
        Red_SubCellInst_LFInst_10_LFInst_0_n19), .ZN(
        Red_SubCellInst_LFInst_10_LFInst_0_n21) );
  INV_X1 Red_SubCellInst_LFInst_10_LFInst_0_U8 ( .A(PermutationOutput[42]), 
        .ZN(Red_SubCellInst_LFInst_10_LFInst_0_n19) );
  NAND2_X1 Red_SubCellInst_LFInst_10_LFInst_0_U7 ( .A1(
        Red_SubCellInst_LFInst_10_LFInst_0_n18), .A2(PermutationOutput[42]), 
        .ZN(Red_SubCellInst_LFInst_10_LFInst_0_n22) );
  XNOR2_X1 Red_SubCellInst_LFInst_10_LFInst_0_U6 ( .A(
        Red_SubCellInst_LFInst_10_LFInst_0_n17), .B(
        Red_SubCellInst_LFInst_10_LFInst_0_n20), .ZN(
        Red_SubCellInst_LFInst_10_LFInst_0_n18) );
  NOR2_X1 Red_SubCellInst_LFInst_10_LFInst_0_U5 ( .A1(
        Red_SubCellInst_LFInst_10_LFInst_0_n16), .A2(
        Red_SubCellInst_LFInst_10_LFInst_0_n15), .ZN(
        Red_SubCellInst_LFInst_10_LFInst_0_n17) );
  INV_X1 Red_SubCellInst_LFInst_10_LFInst_0_U4 ( .A(PermutationOutput[41]), 
        .ZN(Red_SubCellInst_LFInst_10_LFInst_0_n15) );
  INV_X1 Red_SubCellInst_LFInst_10_LFInst_0_U3 ( .A(PermutationOutput[43]), 
        .ZN(Red_SubCellInst_LFInst_10_LFInst_0_n16) );
  OR2_X1 Red_SubCellInst_LFInst_10_LFInst_0_U2 ( .A1(
        Red_SubCellInst_LFInst_10_LFInst_0_n14), .A2(PermutationOutput[40]), 
        .ZN(Red_SubCellInst_LFInst_10_LFInst_0_n20) );
  AND2_X1 Red_SubCellInst_LFInst_10_LFInst_0_U1 ( .A1(
        Red_SubCellInst_LFInst_10_LFInst_0_n15), .A2(
        Red_SubCellInst_LFInst_10_LFInst_0_n16), .ZN(
        Red_SubCellInst_LFInst_10_LFInst_0_n14) );
  AND2_X1 Red_SubCellInst_LFInst_11_LFInst_0_U10 ( .A1(
        Red_SubCellInst_LFInst_11_LFInst_0_n22), .A2(
        Red_SubCellInst_LFInst_11_LFInst_0_n21), .ZN(Red_SboxOut[11]) );
  NAND2_X1 Red_SubCellInst_LFInst_11_LFInst_0_U9 ( .A1(
        Red_SubCellInst_LFInst_11_LFInst_0_n20), .A2(
        Red_SubCellInst_LFInst_11_LFInst_0_n19), .ZN(
        Red_SubCellInst_LFInst_11_LFInst_0_n21) );
  INV_X1 Red_SubCellInst_LFInst_11_LFInst_0_U8 ( .A(PermutationOutput[46]), 
        .ZN(Red_SubCellInst_LFInst_11_LFInst_0_n19) );
  NAND2_X1 Red_SubCellInst_LFInst_11_LFInst_0_U7 ( .A1(
        Red_SubCellInst_LFInst_11_LFInst_0_n18), .A2(PermutationOutput[46]), 
        .ZN(Red_SubCellInst_LFInst_11_LFInst_0_n22) );
  XNOR2_X1 Red_SubCellInst_LFInst_11_LFInst_0_U6 ( .A(
        Red_SubCellInst_LFInst_11_LFInst_0_n17), .B(
        Red_SubCellInst_LFInst_11_LFInst_0_n20), .ZN(
        Red_SubCellInst_LFInst_11_LFInst_0_n18) );
  NOR2_X1 Red_SubCellInst_LFInst_11_LFInst_0_U5 ( .A1(
        Red_SubCellInst_LFInst_11_LFInst_0_n16), .A2(
        Red_SubCellInst_LFInst_11_LFInst_0_n15), .ZN(
        Red_SubCellInst_LFInst_11_LFInst_0_n17) );
  INV_X1 Red_SubCellInst_LFInst_11_LFInst_0_U4 ( .A(PermutationOutput[45]), 
        .ZN(Red_SubCellInst_LFInst_11_LFInst_0_n15) );
  INV_X1 Red_SubCellInst_LFInst_11_LFInst_0_U3 ( .A(PermutationOutput[47]), 
        .ZN(Red_SubCellInst_LFInst_11_LFInst_0_n16) );
  OR2_X1 Red_SubCellInst_LFInst_11_LFInst_0_U2 ( .A1(
        Red_SubCellInst_LFInst_11_LFInst_0_n14), .A2(PermutationOutput[44]), 
        .ZN(Red_SubCellInst_LFInst_11_LFInst_0_n20) );
  AND2_X1 Red_SubCellInst_LFInst_11_LFInst_0_U1 ( .A1(
        Red_SubCellInst_LFInst_11_LFInst_0_n15), .A2(
        Red_SubCellInst_LFInst_11_LFInst_0_n16), .ZN(
        Red_SubCellInst_LFInst_11_LFInst_0_n14) );
  AND2_X1 Red_SubCellInst_LFInst_12_LFInst_0_U10 ( .A1(
        Red_SubCellInst_LFInst_12_LFInst_0_n22), .A2(
        Red_SubCellInst_LFInst_12_LFInst_0_n21), .ZN(Red_SboxOut[12]) );
  NAND2_X1 Red_SubCellInst_LFInst_12_LFInst_0_U9 ( .A1(
        Red_SubCellInst_LFInst_12_LFInst_0_n20), .A2(
        Red_SubCellInst_LFInst_12_LFInst_0_n19), .ZN(
        Red_SubCellInst_LFInst_12_LFInst_0_n21) );
  INV_X1 Red_SubCellInst_LFInst_12_LFInst_0_U8 ( .A(PermutationOutput[50]), 
        .ZN(Red_SubCellInst_LFInst_12_LFInst_0_n19) );
  NAND2_X1 Red_SubCellInst_LFInst_12_LFInst_0_U7 ( .A1(
        Red_SubCellInst_LFInst_12_LFInst_0_n18), .A2(PermutationOutput[50]), 
        .ZN(Red_SubCellInst_LFInst_12_LFInst_0_n22) );
  XNOR2_X1 Red_SubCellInst_LFInst_12_LFInst_0_U6 ( .A(
        Red_SubCellInst_LFInst_12_LFInst_0_n17), .B(
        Red_SubCellInst_LFInst_12_LFInst_0_n20), .ZN(
        Red_SubCellInst_LFInst_12_LFInst_0_n18) );
  NOR2_X1 Red_SubCellInst_LFInst_12_LFInst_0_U5 ( .A1(
        Red_SubCellInst_LFInst_12_LFInst_0_n16), .A2(
        Red_SubCellInst_LFInst_12_LFInst_0_n15), .ZN(
        Red_SubCellInst_LFInst_12_LFInst_0_n17) );
  INV_X1 Red_SubCellInst_LFInst_12_LFInst_0_U4 ( .A(PermutationOutput[49]), 
        .ZN(Red_SubCellInst_LFInst_12_LFInst_0_n15) );
  INV_X1 Red_SubCellInst_LFInst_12_LFInst_0_U3 ( .A(PermutationOutput[51]), 
        .ZN(Red_SubCellInst_LFInst_12_LFInst_0_n16) );
  OR2_X1 Red_SubCellInst_LFInst_12_LFInst_0_U2 ( .A1(
        Red_SubCellInst_LFInst_12_LFInst_0_n14), .A2(PermutationOutput[48]), 
        .ZN(Red_SubCellInst_LFInst_12_LFInst_0_n20) );
  AND2_X1 Red_SubCellInst_LFInst_12_LFInst_0_U1 ( .A1(
        Red_SubCellInst_LFInst_12_LFInst_0_n15), .A2(
        Red_SubCellInst_LFInst_12_LFInst_0_n16), .ZN(
        Red_SubCellInst_LFInst_12_LFInst_0_n14) );
  AND2_X1 Red_SubCellInst_LFInst_13_LFInst_0_U10 ( .A1(
        Red_SubCellInst_LFInst_13_LFInst_0_n22), .A2(
        Red_SubCellInst_LFInst_13_LFInst_0_n21), .ZN(Red_SboxOut[13]) );
  NAND2_X1 Red_SubCellInst_LFInst_13_LFInst_0_U9 ( .A1(
        Red_SubCellInst_LFInst_13_LFInst_0_n20), .A2(
        Red_SubCellInst_LFInst_13_LFInst_0_n19), .ZN(
        Red_SubCellInst_LFInst_13_LFInst_0_n21) );
  INV_X1 Red_SubCellInst_LFInst_13_LFInst_0_U8 ( .A(PermutationOutput[54]), 
        .ZN(Red_SubCellInst_LFInst_13_LFInst_0_n19) );
  NAND2_X1 Red_SubCellInst_LFInst_13_LFInst_0_U7 ( .A1(
        Red_SubCellInst_LFInst_13_LFInst_0_n18), .A2(PermutationOutput[54]), 
        .ZN(Red_SubCellInst_LFInst_13_LFInst_0_n22) );
  XNOR2_X1 Red_SubCellInst_LFInst_13_LFInst_0_U6 ( .A(
        Red_SubCellInst_LFInst_13_LFInst_0_n17), .B(
        Red_SubCellInst_LFInst_13_LFInst_0_n20), .ZN(
        Red_SubCellInst_LFInst_13_LFInst_0_n18) );
  NOR2_X1 Red_SubCellInst_LFInst_13_LFInst_0_U5 ( .A1(
        Red_SubCellInst_LFInst_13_LFInst_0_n16), .A2(
        Red_SubCellInst_LFInst_13_LFInst_0_n15), .ZN(
        Red_SubCellInst_LFInst_13_LFInst_0_n17) );
  INV_X1 Red_SubCellInst_LFInst_13_LFInst_0_U4 ( .A(PermutationOutput[53]), 
        .ZN(Red_SubCellInst_LFInst_13_LFInst_0_n15) );
  INV_X1 Red_SubCellInst_LFInst_13_LFInst_0_U3 ( .A(PermutationOutput[55]), 
        .ZN(Red_SubCellInst_LFInst_13_LFInst_0_n16) );
  OR2_X1 Red_SubCellInst_LFInst_13_LFInst_0_U2 ( .A1(
        Red_SubCellInst_LFInst_13_LFInst_0_n14), .A2(PermutationOutput[52]), 
        .ZN(Red_SubCellInst_LFInst_13_LFInst_0_n20) );
  AND2_X1 Red_SubCellInst_LFInst_13_LFInst_0_U1 ( .A1(
        Red_SubCellInst_LFInst_13_LFInst_0_n15), .A2(
        Red_SubCellInst_LFInst_13_LFInst_0_n16), .ZN(
        Red_SubCellInst_LFInst_13_LFInst_0_n14) );
  AND2_X1 Red_SubCellInst_LFInst_14_LFInst_0_U10 ( .A1(
        Red_SubCellInst_LFInst_14_LFInst_0_n22), .A2(
        Red_SubCellInst_LFInst_14_LFInst_0_n21), .ZN(Red_SboxOut[14]) );
  NAND2_X1 Red_SubCellInst_LFInst_14_LFInst_0_U9 ( .A1(
        Red_SubCellInst_LFInst_14_LFInst_0_n20), .A2(
        Red_SubCellInst_LFInst_14_LFInst_0_n19), .ZN(
        Red_SubCellInst_LFInst_14_LFInst_0_n21) );
  INV_X1 Red_SubCellInst_LFInst_14_LFInst_0_U8 ( .A(PermutationOutput[58]), 
        .ZN(Red_SubCellInst_LFInst_14_LFInst_0_n19) );
  NAND2_X1 Red_SubCellInst_LFInst_14_LFInst_0_U7 ( .A1(
        Red_SubCellInst_LFInst_14_LFInst_0_n18), .A2(PermutationOutput[58]), 
        .ZN(Red_SubCellInst_LFInst_14_LFInst_0_n22) );
  XNOR2_X1 Red_SubCellInst_LFInst_14_LFInst_0_U6 ( .A(
        Red_SubCellInst_LFInst_14_LFInst_0_n17), .B(
        Red_SubCellInst_LFInst_14_LFInst_0_n20), .ZN(
        Red_SubCellInst_LFInst_14_LFInst_0_n18) );
  NOR2_X1 Red_SubCellInst_LFInst_14_LFInst_0_U5 ( .A1(
        Red_SubCellInst_LFInst_14_LFInst_0_n16), .A2(
        Red_SubCellInst_LFInst_14_LFInst_0_n15), .ZN(
        Red_SubCellInst_LFInst_14_LFInst_0_n17) );
  INV_X1 Red_SubCellInst_LFInst_14_LFInst_0_U4 ( .A(PermutationOutput[57]), 
        .ZN(Red_SubCellInst_LFInst_14_LFInst_0_n15) );
  INV_X1 Red_SubCellInst_LFInst_14_LFInst_0_U3 ( .A(PermutationOutput[59]), 
        .ZN(Red_SubCellInst_LFInst_14_LFInst_0_n16) );
  OR2_X1 Red_SubCellInst_LFInst_14_LFInst_0_U2 ( .A1(
        Red_SubCellInst_LFInst_14_LFInst_0_n14), .A2(PermutationOutput[56]), 
        .ZN(Red_SubCellInst_LFInst_14_LFInst_0_n20) );
  AND2_X1 Red_SubCellInst_LFInst_14_LFInst_0_U1 ( .A1(
        Red_SubCellInst_LFInst_14_LFInst_0_n15), .A2(
        Red_SubCellInst_LFInst_14_LFInst_0_n16), .ZN(
        Red_SubCellInst_LFInst_14_LFInst_0_n14) );
  AND2_X1 Red_SubCellInst_LFInst_15_LFInst_0_U10 ( .A1(
        Red_SubCellInst_LFInst_15_LFInst_0_n22), .A2(
        Red_SubCellInst_LFInst_15_LFInst_0_n21), .ZN(Red_SboxOut[15]) );
  NAND2_X1 Red_SubCellInst_LFInst_15_LFInst_0_U9 ( .A1(
        Red_SubCellInst_LFInst_15_LFInst_0_n20), .A2(
        Red_SubCellInst_LFInst_15_LFInst_0_n19), .ZN(
        Red_SubCellInst_LFInst_15_LFInst_0_n21) );
  INV_X1 Red_SubCellInst_LFInst_15_LFInst_0_U8 ( .A(PermutationOutput[62]), 
        .ZN(Red_SubCellInst_LFInst_15_LFInst_0_n19) );
  NAND2_X1 Red_SubCellInst_LFInst_15_LFInst_0_U7 ( .A1(
        Red_SubCellInst_LFInst_15_LFInst_0_n18), .A2(PermutationOutput[62]), 
        .ZN(Red_SubCellInst_LFInst_15_LFInst_0_n22) );
  XNOR2_X1 Red_SubCellInst_LFInst_15_LFInst_0_U6 ( .A(
        Red_SubCellInst_LFInst_15_LFInst_0_n17), .B(
        Red_SubCellInst_LFInst_15_LFInst_0_n20), .ZN(
        Red_SubCellInst_LFInst_15_LFInst_0_n18) );
  NOR2_X1 Red_SubCellInst_LFInst_15_LFInst_0_U5 ( .A1(
        Red_SubCellInst_LFInst_15_LFInst_0_n16), .A2(
        Red_SubCellInst_LFInst_15_LFInst_0_n15), .ZN(
        Red_SubCellInst_LFInst_15_LFInst_0_n17) );
  INV_X1 Red_SubCellInst_LFInst_15_LFInst_0_U4 ( .A(PermutationOutput[61]), 
        .ZN(Red_SubCellInst_LFInst_15_LFInst_0_n15) );
  INV_X1 Red_SubCellInst_LFInst_15_LFInst_0_U3 ( .A(PermutationOutput[63]), 
        .ZN(Red_SubCellInst_LFInst_15_LFInst_0_n16) );
  OR2_X1 Red_SubCellInst_LFInst_15_LFInst_0_U2 ( .A1(
        Red_SubCellInst_LFInst_15_LFInst_0_n14), .A2(PermutationOutput[60]), 
        .ZN(Red_SubCellInst_LFInst_15_LFInst_0_n20) );
  AND2_X1 Red_SubCellInst_LFInst_15_LFInst_0_U1 ( .A1(
        Red_SubCellInst_LFInst_15_LFInst_0_n15), .A2(
        Red_SubCellInst_LFInst_15_LFInst_0_n16), .ZN(
        Red_SubCellInst_LFInst_15_LFInst_0_n14) );
  XNOR2_X1 Red_MCInst2_XOR_r0_Inst_0_U2 ( .A(Red_MCInst2_XOR_r0_Inst_0_n5), 
        .B(Red_MCOutput2[4]), .ZN(Red_MCOutput2[12]) );
  XNOR2_X1 Red_MCInst2_XOR_r0_Inst_0_U1 ( .A(Red_MCOutput2[0]), .B(
        Red_SboxOut[12]), .ZN(Red_MCInst2_XOR_r0_Inst_0_n5) );
  XOR2_X1 Red_MCInst2_XOR_r1_Inst_0_U1 ( .A(Red_SboxOut[8]), .B(
        Red_MCOutput2[0]), .Z(Red_MCOutput2[8]) );
  XNOR2_X1 Red_MCInst2_XOR_r0_Inst_1_U2 ( .A(Red_MCInst2_XOR_r0_Inst_1_n5), 
        .B(Red_MCOutput2[5]), .ZN(Red_MCOutput2[13]) );
  XNOR2_X1 Red_MCInst2_XOR_r0_Inst_1_U1 ( .A(Red_MCOutput2[1]), .B(
        Red_SboxOut[13]), .ZN(Red_MCInst2_XOR_r0_Inst_1_n5) );
  XOR2_X1 Red_MCInst2_XOR_r1_Inst_1_U1 ( .A(Red_SboxOut[9]), .B(
        Red_MCOutput2[1]), .Z(Red_MCOutput2[9]) );
  XNOR2_X1 Red_MCInst2_XOR_r0_Inst_2_U2 ( .A(Red_MCInst2_XOR_r0_Inst_2_n5), 
        .B(Red_MCOutput2[6]), .ZN(Red_MCOutput2[14]) );
  XNOR2_X1 Red_MCInst2_XOR_r0_Inst_2_U1 ( .A(Red_MCOutput2[2]), .B(
        Red_SboxOut[14]), .ZN(Red_MCInst2_XOR_r0_Inst_2_n5) );
  XOR2_X1 Red_MCInst2_XOR_r1_Inst_2_U1 ( .A(Red_SboxOut[10]), .B(
        Red_MCOutput2[2]), .Z(Red_MCOutput2[10]) );
  XNOR2_X1 Red_MCInst2_XOR_r0_Inst_3_U2 ( .A(Red_MCInst2_XOR_r0_Inst_3_n5), 
        .B(Red_MCOutput2[7]), .ZN(Red_MCOutput2[15]) );
  XNOR2_X1 Red_MCInst2_XOR_r0_Inst_3_U1 ( .A(Red_MCOutput2[3]), .B(
        Red_SboxOut[15]), .ZN(Red_MCInst2_XOR_r0_Inst_3_n5) );
  XOR2_X1 Red_MCInst2_XOR_r1_Inst_3_U1 ( .A(Red_SboxOut[11]), .B(
        Red_MCOutput2[3]), .Z(Red_MCOutput2[11]) );
  XOR2_X1 Red_AddKeyXOR12_XORInst_0_0_U1 ( .A(Red_MCOutput2[12]), .B(
        Red_K1[12]), .Z(Red_final[12]) );
  XOR2_X1 Red_AddKeyXOR12_XORInst_1_0_U1 ( .A(Red_MCOutput2[13]), .B(
        Red_K1[13]), .Z(Red_final[13]) );
  XOR2_X1 Red_AddKeyXOR12_XORInst_2_0_U1 ( .A(Red_MCOutput2[14]), .B(
        Red_K1[14]), .Z(Red_final[14]) );
  XOR2_X1 Red_AddKeyXOR12_XORInst_3_0_U1 ( .A(Red_MCOutput2[15]), .B(
        Red_K1[15]), .Z(Red_final[15]) );
  XOR2_X1 Red_AddKeyConstXOR2_XORInst_0_0_U1 ( .A(Red_MCOutput2[10]), .B(
        Red_K1[10]), .Z(Red_final[10]) );
  XOR2_X1 Red_AddKeyConstXOR2_XORInst_1_0_U1 ( .A(Red_MCOutput2[11]), .B(
        Red_K1[11]), .Z(Red_final[11]) );
  XOR2_X1 Red_AddKeyXOR22_XORInst_0_0_U1 ( .A(Red_MCOutput2[0]), .B(Red_K1[0]), 
        .Z(Red_final[0]) );
  XOR2_X1 Red_AddKeyXOR22_XORInst_1_0_U1 ( .A(Red_MCOutput2[1]), .B(Red_K1[1]), 
        .Z(Red_final[1]) );
  XOR2_X1 Red_AddKeyXOR22_XORInst_2_0_U1 ( .A(Red_MCOutput2[2]), .B(Red_K1[2]), 
        .Z(Red_final[2]) );
  XOR2_X1 Red_AddKeyXOR22_XORInst_3_0_U1 ( .A(Red_MCOutput2[3]), .B(Red_K1[3]), 
        .Z(Red_final[3]) );
  XOR2_X1 Red_AddKeyXOR22_XORInst_4_0_U1 ( .A(Red_MCOutput2[4]), .B(Red_K1[4]), 
        .Z(Red_final[4]) );
  XOR2_X1 Red_AddKeyXOR22_XORInst_5_0_U1 ( .A(Red_MCOutput2[5]), .B(Red_K1[5]), 
        .Z(Red_final[5]) );
  XOR2_X1 Red_AddKeyXOR22_XORInst_6_0_U1 ( .A(Red_MCOutput2[6]), .B(Red_K1[6]), 
        .Z(Red_final[6]) );
  XOR2_X1 Red_AddKeyXOR22_XORInst_7_0_U1 ( .A(Red_MCOutput2[7]), .B(Red_K1[7]), 
        .Z(Red_final[7]) );
  XOR2_X1 Red_AddKeyXOR22_XORInst_8_0_U1 ( .A(Red_MCOutput2[8]), .B(Red_K1[8]), 
        .Z(Red_final[8]) );
  XOR2_X1 Red_AddKeyXOR22_XORInst_9_0_U1 ( .A(Red_MCOutput2[9]), .B(Red_K1[9]), 
        .Z(Red_final[9]) );
  DFF_X1 Red_StateReg2_s_current_state_reg_0_ ( .D(Red_final[0]), .CK(clk), 
        .Q(Red_StateRegOutput2[0]), .QN() );
  DFF_X1 Red_StateReg2_s_current_state_reg_1_ ( .D(Red_final[1]), .CK(clk), 
        .Q(Red_StateRegOutput2[1]), .QN() );
  DFF_X1 Red_StateReg2_s_current_state_reg_2_ ( .D(Red_final[2]), .CK(clk), 
        .Q(Red_StateRegOutput2[2]), .QN() );
  DFF_X1 Red_StateReg2_s_current_state_reg_3_ ( .D(Red_final[3]), .CK(clk), 
        .Q(Red_StateRegOutput2[3]), .QN() );
  DFF_X1 Red_StateReg2_s_current_state_reg_4_ ( .D(Red_final[4]), .CK(clk), 
        .Q(Red_StateRegOutput2[4]), .QN() );
  DFF_X1 Red_StateReg2_s_current_state_reg_5_ ( .D(Red_final[5]), .CK(clk), 
        .Q(Red_StateRegOutput2[5]), .QN() );
  DFF_X1 Red_StateReg2_s_current_state_reg_6_ ( .D(Red_final[6]), .CK(clk), 
        .Q(Red_StateRegOutput2[6]), .QN() );
  DFF_X1 Red_StateReg2_s_current_state_reg_7_ ( .D(Red_final[7]), .CK(clk), 
        .Q(Red_StateRegOutput2[7]), .QN() );
  DFF_X1 Red_StateReg2_s_current_state_reg_8_ ( .D(Red_final[8]), .CK(clk), 
        .Q(Red_StateRegOutput2[8]), .QN() );
  DFF_X1 Red_StateReg2_s_current_state_reg_9_ ( .D(Red_final[9]), .CK(clk), 
        .Q(Red_StateRegOutput2[9]), .QN() );
  DFF_X1 Red_StateReg2_s_current_state_reg_10_ ( .D(Red_final[10]), .CK(clk), 
        .Q(Red_StateRegOutput2[10]), .QN() );
  DFF_X1 Red_StateReg2_s_current_state_reg_11_ ( .D(Red_final[11]), .CK(clk), 
        .Q(Red_StateRegOutput2[11]), .QN() );
  DFF_X1 Red_StateReg2_s_current_state_reg_12_ ( .D(Red_final[12]), .CK(clk), 
        .Q(Red_StateRegOutput2[12]), .QN() );
  DFF_X1 Red_StateReg2_s_current_state_reg_13_ ( .D(Red_final[13]), .CK(clk), 
        .Q(Red_StateRegOutput2[13]), .QN() );
  DFF_X1 Red_StateReg2_s_current_state_reg_14_ ( .D(Red_final[14]), .CK(clk), 
        .Q(Red_StateRegOutput2[14]), .QN() );
  DFF_X1 Red_StateReg2_s_current_state_reg_15_ ( .D(Red_final[15]), .CK(clk), 
        .Q(Red_StateRegOutput2[15]), .QN() );
  XNOR2_X1 Red_SubCellInst2_LFInst_0_LFInst_0_U5 ( .A(
        Red_SubCellInst2_LFInst_0_LFInst_0_n15), .B(
        Red_SubCellInst2_LFInst_0_LFInst_0_n17), .ZN(Red_Feedback[0]) );
  NOR2_X1 Red_SubCellInst2_LFInst_0_LFInst_0_U4 ( .A1(PermutationOutput2[0]), 
        .A2(Red_SubCellInst2_LFInst_0_LFInst_0_n16), .ZN(
        Red_SubCellInst2_LFInst_0_LFInst_0_n17) );
  NOR2_X1 Red_SubCellInst2_LFInst_0_LFInst_0_U3 ( .A1(PermutationOutput2[3]), 
        .A2(PermutationOutput2[1]), .ZN(Red_SubCellInst2_LFInst_0_LFInst_0_n16) );
  NAND2_X1 Red_SubCellInst2_LFInst_0_LFInst_0_U2 ( .A1(
        Red_SubCellInst2_LFInst_0_LFInst_0_n14), .A2(PermutationOutput2[2]), 
        .ZN(Red_SubCellInst2_LFInst_0_LFInst_0_n15) );
  NAND2_X1 Red_SubCellInst2_LFInst_0_LFInst_0_U1 ( .A1(PermutationOutput2[1]), 
        .A2(PermutationOutput2[3]), .ZN(Red_SubCellInst2_LFInst_0_LFInst_0_n14) );
  NAND2_X1 Red_SubCellInst2_LFInst_1_LFInst_0_U7 ( .A1(
        Red_SubCellInst2_LFInst_1_LFInst_0_n17), .A2(
        Red_SubCellInst2_LFInst_1_LFInst_0_n21), .ZN(Red_Feedback[1]) );
  NAND2_X1 Red_SubCellInst2_LFInst_1_LFInst_0_U6 ( .A1(
        Red_SubCellInst2_LFInst_1_LFInst_0_n20), .A2(
        Red_SubCellInst2_LFInst_1_LFInst_0_n16), .ZN(
        Red_SubCellInst2_LFInst_1_LFInst_0_n21) );
  XOR2_X1 Red_SubCellInst2_LFInst_1_LFInst_0_U5 ( .A(PermutationOutput2[6]), 
        .B(Red_SubCellInst2_LFInst_1_LFInst_0_n19), .Z(
        Red_SubCellInst2_LFInst_1_LFInst_0_n20) );
  NOR2_X1 Red_SubCellInst2_LFInst_1_LFInst_0_U4 ( .A1(PermutationOutput2[4]), 
        .A2(Red_SubCellInst2_LFInst_1_LFInst_0_n18), .ZN(
        Red_SubCellInst2_LFInst_1_LFInst_0_n19) );
  NOR2_X1 Red_SubCellInst2_LFInst_1_LFInst_0_U3 ( .A1(PermutationOutput2[7]), 
        .A2(PermutationOutput2[5]), .ZN(Red_SubCellInst2_LFInst_1_LFInst_0_n18) );
  OR2_X1 Red_SubCellInst2_LFInst_1_LFInst_0_U2 ( .A1(PermutationOutput2[4]), 
        .A2(Red_SubCellInst2_LFInst_1_LFInst_0_n16), .ZN(
        Red_SubCellInst2_LFInst_1_LFInst_0_n17) );
  NAND2_X1 Red_SubCellInst2_LFInst_1_LFInst_0_U1 ( .A1(PermutationOutput2[7]), 
        .A2(PermutationOutput2[5]), .ZN(Red_SubCellInst2_LFInst_1_LFInst_0_n16) );
  XNOR2_X1 Red_SubCellInst2_LFInst_2_LFInst_0_U5 ( .A(
        Red_SubCellInst2_LFInst_2_LFInst_0_n15), .B(
        Red_SubCellInst2_LFInst_2_LFInst_0_n17), .ZN(Red_Feedback[2]) );
  NOR2_X1 Red_SubCellInst2_LFInst_2_LFInst_0_U4 ( .A1(PermutationOutput2[8]), 
        .A2(Red_SubCellInst2_LFInst_2_LFInst_0_n16), .ZN(
        Red_SubCellInst2_LFInst_2_LFInst_0_n17) );
  NOR2_X1 Red_SubCellInst2_LFInst_2_LFInst_0_U3 ( .A1(PermutationOutput2[11]), 
        .A2(PermutationOutput2[9]), .ZN(Red_SubCellInst2_LFInst_2_LFInst_0_n16) );
  NAND2_X1 Red_SubCellInst2_LFInst_2_LFInst_0_U2 ( .A1(
        Red_SubCellInst2_LFInst_2_LFInst_0_n14), .A2(PermutationOutput2[10]), 
        .ZN(Red_SubCellInst2_LFInst_2_LFInst_0_n15) );
  NAND2_X1 Red_SubCellInst2_LFInst_2_LFInst_0_U1 ( .A1(PermutationOutput2[9]), 
        .A2(PermutationOutput2[11]), .ZN(
        Red_SubCellInst2_LFInst_2_LFInst_0_n14) );
  XNOR2_X1 Red_SubCellInst2_LFInst_3_LFInst_0_U5 ( .A(
        Red_SubCellInst2_LFInst_3_LFInst_0_n15), .B(
        Red_SubCellInst2_LFInst_3_LFInst_0_n17), .ZN(Red_Feedback[3]) );
  NOR2_X1 Red_SubCellInst2_LFInst_3_LFInst_0_U4 ( .A1(PermutationOutput2[12]), 
        .A2(Red_SubCellInst2_LFInst_3_LFInst_0_n16), .ZN(
        Red_SubCellInst2_LFInst_3_LFInst_0_n17) );
  NOR2_X1 Red_SubCellInst2_LFInst_3_LFInst_0_U3 ( .A1(PermutationOutput2[15]), 
        .A2(PermutationOutput2[13]), .ZN(
        Red_SubCellInst2_LFInst_3_LFInst_0_n16) );
  NAND2_X1 Red_SubCellInst2_LFInst_3_LFInst_0_U2 ( .A1(
        Red_SubCellInst2_LFInst_3_LFInst_0_n14), .A2(PermutationOutput2[14]), 
        .ZN(Red_SubCellInst2_LFInst_3_LFInst_0_n15) );
  NAND2_X1 Red_SubCellInst2_LFInst_3_LFInst_0_U1 ( .A1(PermutationOutput2[13]), 
        .A2(PermutationOutput2[15]), .ZN(
        Red_SubCellInst2_LFInst_3_LFInst_0_n14) );
  AND2_X1 Red_SubCellInst2_LFInst_4_LFInst_0_U10 ( .A1(
        Red_SubCellInst2_LFInst_4_LFInst_0_n22), .A2(
        Red_SubCellInst2_LFInst_4_LFInst_0_n21), .ZN(Red_Feedback[4]) );
  NAND2_X1 Red_SubCellInst2_LFInst_4_LFInst_0_U9 ( .A1(
        Red_SubCellInst2_LFInst_4_LFInst_0_n20), .A2(
        Red_SubCellInst2_LFInst_4_LFInst_0_n19), .ZN(
        Red_SubCellInst2_LFInst_4_LFInst_0_n21) );
  INV_X1 Red_SubCellInst2_LFInst_4_LFInst_0_U8 ( .A(PermutationOutput2[18]), 
        .ZN(Red_SubCellInst2_LFInst_4_LFInst_0_n19) );
  NAND2_X1 Red_SubCellInst2_LFInst_4_LFInst_0_U7 ( .A1(
        Red_SubCellInst2_LFInst_4_LFInst_0_n18), .A2(PermutationOutput2[18]), 
        .ZN(Red_SubCellInst2_LFInst_4_LFInst_0_n22) );
  XNOR2_X1 Red_SubCellInst2_LFInst_4_LFInst_0_U6 ( .A(
        Red_SubCellInst2_LFInst_4_LFInst_0_n17), .B(
        Red_SubCellInst2_LFInst_4_LFInst_0_n20), .ZN(
        Red_SubCellInst2_LFInst_4_LFInst_0_n18) );
  NOR2_X1 Red_SubCellInst2_LFInst_4_LFInst_0_U5 ( .A1(
        Red_SubCellInst2_LFInst_4_LFInst_0_n16), .A2(
        Red_SubCellInst2_LFInst_4_LFInst_0_n15), .ZN(
        Red_SubCellInst2_LFInst_4_LFInst_0_n17) );
  INV_X1 Red_SubCellInst2_LFInst_4_LFInst_0_U4 ( .A(PermutationOutput2[17]), 
        .ZN(Red_SubCellInst2_LFInst_4_LFInst_0_n15) );
  INV_X1 Red_SubCellInst2_LFInst_4_LFInst_0_U3 ( .A(PermutationOutput2[19]), 
        .ZN(Red_SubCellInst2_LFInst_4_LFInst_0_n16) );
  OR2_X1 Red_SubCellInst2_LFInst_4_LFInst_0_U2 ( .A1(
        Red_SubCellInst2_LFInst_4_LFInst_0_n14), .A2(PermutationOutput2[16]), 
        .ZN(Red_SubCellInst2_LFInst_4_LFInst_0_n20) );
  AND2_X1 Red_SubCellInst2_LFInst_4_LFInst_0_U1 ( .A1(
        Red_SubCellInst2_LFInst_4_LFInst_0_n15), .A2(
        Red_SubCellInst2_LFInst_4_LFInst_0_n16), .ZN(
        Red_SubCellInst2_LFInst_4_LFInst_0_n14) );
  XNOR2_X1 Red_SubCellInst2_LFInst_5_LFInst_0_U5 ( .A(
        Red_SubCellInst2_LFInst_5_LFInst_0_n15), .B(
        Red_SubCellInst2_LFInst_5_LFInst_0_n17), .ZN(Red_Feedback[5]) );
  NOR2_X1 Red_SubCellInst2_LFInst_5_LFInst_0_U4 ( .A1(PermutationOutput2[20]), 
        .A2(Red_SubCellInst2_LFInst_5_LFInst_0_n16), .ZN(
        Red_SubCellInst2_LFInst_5_LFInst_0_n17) );
  NOR2_X1 Red_SubCellInst2_LFInst_5_LFInst_0_U3 ( .A1(PermutationOutput2[23]), 
        .A2(PermutationOutput2[21]), .ZN(
        Red_SubCellInst2_LFInst_5_LFInst_0_n16) );
  NAND2_X1 Red_SubCellInst2_LFInst_5_LFInst_0_U2 ( .A1(
        Red_SubCellInst2_LFInst_5_LFInst_0_n14), .A2(PermutationOutput2[22]), 
        .ZN(Red_SubCellInst2_LFInst_5_LFInst_0_n15) );
  NAND2_X1 Red_SubCellInst2_LFInst_5_LFInst_0_U1 ( .A1(PermutationOutput2[21]), 
        .A2(PermutationOutput2[23]), .ZN(
        Red_SubCellInst2_LFInst_5_LFInst_0_n14) );
  AND2_X1 Red_SubCellInst2_LFInst_6_LFInst_0_U10 ( .A1(
        Red_SubCellInst2_LFInst_6_LFInst_0_n22), .A2(
        Red_SubCellInst2_LFInst_6_LFInst_0_n21), .ZN(Red_Feedback[6]) );
  NAND2_X1 Red_SubCellInst2_LFInst_6_LFInst_0_U9 ( .A1(
        Red_SubCellInst2_LFInst_6_LFInst_0_n20), .A2(
        Red_SubCellInst2_LFInst_6_LFInst_0_n19), .ZN(
        Red_SubCellInst2_LFInst_6_LFInst_0_n21) );
  INV_X1 Red_SubCellInst2_LFInst_6_LFInst_0_U8 ( .A(PermutationOutput2[26]), 
        .ZN(Red_SubCellInst2_LFInst_6_LFInst_0_n19) );
  NAND2_X1 Red_SubCellInst2_LFInst_6_LFInst_0_U7 ( .A1(
        Red_SubCellInst2_LFInst_6_LFInst_0_n18), .A2(PermutationOutput2[26]), 
        .ZN(Red_SubCellInst2_LFInst_6_LFInst_0_n22) );
  XNOR2_X1 Red_SubCellInst2_LFInst_6_LFInst_0_U6 ( .A(
        Red_SubCellInst2_LFInst_6_LFInst_0_n17), .B(
        Red_SubCellInst2_LFInst_6_LFInst_0_n20), .ZN(
        Red_SubCellInst2_LFInst_6_LFInst_0_n18) );
  NOR2_X1 Red_SubCellInst2_LFInst_6_LFInst_0_U5 ( .A1(
        Red_SubCellInst2_LFInst_6_LFInst_0_n16), .A2(
        Red_SubCellInst2_LFInst_6_LFInst_0_n15), .ZN(
        Red_SubCellInst2_LFInst_6_LFInst_0_n17) );
  INV_X1 Red_SubCellInst2_LFInst_6_LFInst_0_U4 ( .A(PermutationOutput2[25]), 
        .ZN(Red_SubCellInst2_LFInst_6_LFInst_0_n15) );
  INV_X1 Red_SubCellInst2_LFInst_6_LFInst_0_U3 ( .A(PermutationOutput2[27]), 
        .ZN(Red_SubCellInst2_LFInst_6_LFInst_0_n16) );
  OR2_X1 Red_SubCellInst2_LFInst_6_LFInst_0_U2 ( .A1(
        Red_SubCellInst2_LFInst_6_LFInst_0_n14), .A2(PermutationOutput2[24]), 
        .ZN(Red_SubCellInst2_LFInst_6_LFInst_0_n20) );
  AND2_X1 Red_SubCellInst2_LFInst_6_LFInst_0_U1 ( .A1(
        Red_SubCellInst2_LFInst_6_LFInst_0_n15), .A2(
        Red_SubCellInst2_LFInst_6_LFInst_0_n16), .ZN(
        Red_SubCellInst2_LFInst_6_LFInst_0_n14) );
  AND2_X1 Red_SubCellInst2_LFInst_7_LFInst_0_U10 ( .A1(
        Red_SubCellInst2_LFInst_7_LFInst_0_n22), .A2(
        Red_SubCellInst2_LFInst_7_LFInst_0_n21), .ZN(Red_Feedback[7]) );
  NAND2_X1 Red_SubCellInst2_LFInst_7_LFInst_0_U9 ( .A1(
        Red_SubCellInst2_LFInst_7_LFInst_0_n20), .A2(
        Red_SubCellInst2_LFInst_7_LFInst_0_n19), .ZN(
        Red_SubCellInst2_LFInst_7_LFInst_0_n21) );
  INV_X1 Red_SubCellInst2_LFInst_7_LFInst_0_U8 ( .A(PermutationOutput2[30]), 
        .ZN(Red_SubCellInst2_LFInst_7_LFInst_0_n19) );
  NAND2_X1 Red_SubCellInst2_LFInst_7_LFInst_0_U7 ( .A1(
        Red_SubCellInst2_LFInst_7_LFInst_0_n18), .A2(PermutationOutput2[30]), 
        .ZN(Red_SubCellInst2_LFInst_7_LFInst_0_n22) );
  XNOR2_X1 Red_SubCellInst2_LFInst_7_LFInst_0_U6 ( .A(
        Red_SubCellInst2_LFInst_7_LFInst_0_n17), .B(
        Red_SubCellInst2_LFInst_7_LFInst_0_n20), .ZN(
        Red_SubCellInst2_LFInst_7_LFInst_0_n18) );
  NOR2_X1 Red_SubCellInst2_LFInst_7_LFInst_0_U5 ( .A1(
        Red_SubCellInst2_LFInst_7_LFInst_0_n16), .A2(
        Red_SubCellInst2_LFInst_7_LFInst_0_n15), .ZN(
        Red_SubCellInst2_LFInst_7_LFInst_0_n17) );
  INV_X1 Red_SubCellInst2_LFInst_7_LFInst_0_U4 ( .A(PermutationOutput2[29]), 
        .ZN(Red_SubCellInst2_LFInst_7_LFInst_0_n15) );
  INV_X1 Red_SubCellInst2_LFInst_7_LFInst_0_U3 ( .A(PermutationOutput2[31]), 
        .ZN(Red_SubCellInst2_LFInst_7_LFInst_0_n16) );
  OR2_X1 Red_SubCellInst2_LFInst_7_LFInst_0_U2 ( .A1(
        Red_SubCellInst2_LFInst_7_LFInst_0_n14), .A2(PermutationOutput2[28]), 
        .ZN(Red_SubCellInst2_LFInst_7_LFInst_0_n20) );
  AND2_X1 Red_SubCellInst2_LFInst_7_LFInst_0_U1 ( .A1(
        Red_SubCellInst2_LFInst_7_LFInst_0_n15), .A2(
        Red_SubCellInst2_LFInst_7_LFInst_0_n16), .ZN(
        Red_SubCellInst2_LFInst_7_LFInst_0_n14) );
  XNOR2_X1 Red_SubCellInst2_LFInst_8_LFInst_0_U5 ( .A(
        Red_SubCellInst2_LFInst_8_LFInst_0_n17), .B(
        Red_SubCellInst2_LFInst_8_LFInst_0_n15), .ZN(Red_Feedback[8]) );
  NAND2_X1 Red_SubCellInst2_LFInst_8_LFInst_0_U4 ( .A1(
        Red_SubCellInst2_LFInst_8_LFInst_0_n16), .A2(PermutationOutput2[34]), 
        .ZN(Red_SubCellInst2_LFInst_8_LFInst_0_n17) );
  NAND2_X1 Red_SubCellInst2_LFInst_8_LFInst_0_U3 ( .A1(PermutationOutput2[33]), 
        .A2(PermutationOutput2[35]), .ZN(
        Red_SubCellInst2_LFInst_8_LFInst_0_n16) );
  NOR2_X1 Red_SubCellInst2_LFInst_8_LFInst_0_U2 ( .A1(PermutationOutput2[32]), 
        .A2(Red_SubCellInst2_LFInst_8_LFInst_0_n14), .ZN(
        Red_SubCellInst2_LFInst_8_LFInst_0_n15) );
  NOR2_X1 Red_SubCellInst2_LFInst_8_LFInst_0_U1 ( .A1(PermutationOutput2[35]), 
        .A2(PermutationOutput2[33]), .ZN(
        Red_SubCellInst2_LFInst_8_LFInst_0_n14) );
  XNOR2_X1 Red_SubCellInst2_LFInst_9_LFInst_0_U5 ( .A(
        Red_SubCellInst2_LFInst_9_LFInst_0_n15), .B(
        Red_SubCellInst2_LFInst_9_LFInst_0_n17), .ZN(Red_Feedback[9]) );
  NOR2_X1 Red_SubCellInst2_LFInst_9_LFInst_0_U4 ( .A1(PermutationOutput2[36]), 
        .A2(Red_SubCellInst2_LFInst_9_LFInst_0_n16), .ZN(
        Red_SubCellInst2_LFInst_9_LFInst_0_n17) );
  NOR2_X1 Red_SubCellInst2_LFInst_9_LFInst_0_U3 ( .A1(PermutationOutput2[39]), 
        .A2(PermutationOutput2[37]), .ZN(
        Red_SubCellInst2_LFInst_9_LFInst_0_n16) );
  NAND2_X1 Red_SubCellInst2_LFInst_9_LFInst_0_U2 ( .A1(
        Red_SubCellInst2_LFInst_9_LFInst_0_n14), .A2(PermutationOutput2[38]), 
        .ZN(Red_SubCellInst2_LFInst_9_LFInst_0_n15) );
  NAND2_X1 Red_SubCellInst2_LFInst_9_LFInst_0_U1 ( .A1(PermutationOutput2[37]), 
        .A2(PermutationOutput2[39]), .ZN(
        Red_SubCellInst2_LFInst_9_LFInst_0_n14) );
  AND2_X1 Red_SubCellInst2_LFInst_10_LFInst_0_U10 ( .A1(
        Red_SubCellInst2_LFInst_10_LFInst_0_n22), .A2(
        Red_SubCellInst2_LFInst_10_LFInst_0_n21), .ZN(Red_Feedback[10]) );
  NAND2_X1 Red_SubCellInst2_LFInst_10_LFInst_0_U9 ( .A1(
        Red_SubCellInst2_LFInst_10_LFInst_0_n20), .A2(
        Red_SubCellInst2_LFInst_10_LFInst_0_n19), .ZN(
        Red_SubCellInst2_LFInst_10_LFInst_0_n21) );
  INV_X1 Red_SubCellInst2_LFInst_10_LFInst_0_U8 ( .A(PermutationOutput2[42]), 
        .ZN(Red_SubCellInst2_LFInst_10_LFInst_0_n19) );
  NAND2_X1 Red_SubCellInst2_LFInst_10_LFInst_0_U7 ( .A1(
        Red_SubCellInst2_LFInst_10_LFInst_0_n18), .A2(PermutationOutput2[42]), 
        .ZN(Red_SubCellInst2_LFInst_10_LFInst_0_n22) );
  XNOR2_X1 Red_SubCellInst2_LFInst_10_LFInst_0_U6 ( .A(
        Red_SubCellInst2_LFInst_10_LFInst_0_n17), .B(
        Red_SubCellInst2_LFInst_10_LFInst_0_n20), .ZN(
        Red_SubCellInst2_LFInst_10_LFInst_0_n18) );
  NOR2_X1 Red_SubCellInst2_LFInst_10_LFInst_0_U5 ( .A1(
        Red_SubCellInst2_LFInst_10_LFInst_0_n16), .A2(
        Red_SubCellInst2_LFInst_10_LFInst_0_n15), .ZN(
        Red_SubCellInst2_LFInst_10_LFInst_0_n17) );
  INV_X1 Red_SubCellInst2_LFInst_10_LFInst_0_U4 ( .A(PermutationOutput2[41]), 
        .ZN(Red_SubCellInst2_LFInst_10_LFInst_0_n15) );
  INV_X1 Red_SubCellInst2_LFInst_10_LFInst_0_U3 ( .A(PermutationOutput2[43]), 
        .ZN(Red_SubCellInst2_LFInst_10_LFInst_0_n16) );
  OR2_X1 Red_SubCellInst2_LFInst_10_LFInst_0_U2 ( .A1(
        Red_SubCellInst2_LFInst_10_LFInst_0_n14), .A2(PermutationOutput2[40]), 
        .ZN(Red_SubCellInst2_LFInst_10_LFInst_0_n20) );
  AND2_X1 Red_SubCellInst2_LFInst_10_LFInst_0_U1 ( .A1(
        Red_SubCellInst2_LFInst_10_LFInst_0_n15), .A2(
        Red_SubCellInst2_LFInst_10_LFInst_0_n16), .ZN(
        Red_SubCellInst2_LFInst_10_LFInst_0_n14) );
  XNOR2_X1 Red_SubCellInst2_LFInst_11_LFInst_0_U5 ( .A(
        Red_SubCellInst2_LFInst_11_LFInst_0_n15), .B(
        Red_SubCellInst2_LFInst_11_LFInst_0_n17), .ZN(Red_Feedback[11]) );
  NOR2_X1 Red_SubCellInst2_LFInst_11_LFInst_0_U4 ( .A1(PermutationOutput2[44]), 
        .A2(Red_SubCellInst2_LFInst_11_LFInst_0_n16), .ZN(
        Red_SubCellInst2_LFInst_11_LFInst_0_n17) );
  NOR2_X1 Red_SubCellInst2_LFInst_11_LFInst_0_U3 ( .A1(PermutationOutput2[47]), 
        .A2(PermutationOutput2[45]), .ZN(
        Red_SubCellInst2_LFInst_11_LFInst_0_n16) );
  NAND2_X1 Red_SubCellInst2_LFInst_11_LFInst_0_U2 ( .A1(
        Red_SubCellInst2_LFInst_11_LFInst_0_n14), .A2(PermutationOutput2[46]), 
        .ZN(Red_SubCellInst2_LFInst_11_LFInst_0_n15) );
  NAND2_X1 Red_SubCellInst2_LFInst_11_LFInst_0_U1 ( .A1(PermutationOutput2[45]), .A2(PermutationOutput2[47]), .ZN(Red_SubCellInst2_LFInst_11_LFInst_0_n14) );
  NAND2_X1 Red_SubCellInst2_LFInst_12_LFInst_0_U7 ( .A1(
        Red_SubCellInst2_LFInst_12_LFInst_0_n17), .A2(
        Red_SubCellInst2_LFInst_12_LFInst_0_n21), .ZN(Red_Feedback[12]) );
  NAND2_X1 Red_SubCellInst2_LFInst_12_LFInst_0_U6 ( .A1(
        Red_SubCellInst2_LFInst_12_LFInst_0_n20), .A2(
        Red_SubCellInst2_LFInst_12_LFInst_0_n16), .ZN(
        Red_SubCellInst2_LFInst_12_LFInst_0_n21) );
  XOR2_X1 Red_SubCellInst2_LFInst_12_LFInst_0_U5 ( .A(PermutationOutput2[50]), 
        .B(Red_SubCellInst2_LFInst_12_LFInst_0_n19), .Z(
        Red_SubCellInst2_LFInst_12_LFInst_0_n20) );
  NOR2_X1 Red_SubCellInst2_LFInst_12_LFInst_0_U4 ( .A1(PermutationOutput2[48]), 
        .A2(Red_SubCellInst2_LFInst_12_LFInst_0_n18), .ZN(
        Red_SubCellInst2_LFInst_12_LFInst_0_n19) );
  NOR2_X1 Red_SubCellInst2_LFInst_12_LFInst_0_U3 ( .A1(PermutationOutput2[51]), 
        .A2(PermutationOutput2[49]), .ZN(
        Red_SubCellInst2_LFInst_12_LFInst_0_n18) );
  OR2_X1 Red_SubCellInst2_LFInst_12_LFInst_0_U2 ( .A1(PermutationOutput2[48]), 
        .A2(Red_SubCellInst2_LFInst_12_LFInst_0_n16), .ZN(
        Red_SubCellInst2_LFInst_12_LFInst_0_n17) );
  NAND2_X1 Red_SubCellInst2_LFInst_12_LFInst_0_U1 ( .A1(PermutationOutput2[51]), .A2(PermutationOutput2[49]), .ZN(Red_SubCellInst2_LFInst_12_LFInst_0_n16) );
  XNOR2_X1 Red_SubCellInst2_LFInst_13_LFInst_0_U5 ( .A(
        Red_SubCellInst2_LFInst_13_LFInst_0_n17), .B(
        Red_SubCellInst2_LFInst_13_LFInst_0_n15), .ZN(Red_Feedback[13]) );
  NAND2_X1 Red_SubCellInst2_LFInst_13_LFInst_0_U4 ( .A1(
        Red_SubCellInst2_LFInst_13_LFInst_0_n16), .A2(PermutationOutput2[54]), 
        .ZN(Red_SubCellInst2_LFInst_13_LFInst_0_n17) );
  NAND2_X1 Red_SubCellInst2_LFInst_13_LFInst_0_U3 ( .A1(PermutationOutput2[53]), .A2(PermutationOutput2[55]), .ZN(Red_SubCellInst2_LFInst_13_LFInst_0_n16) );
  NOR2_X1 Red_SubCellInst2_LFInst_13_LFInst_0_U2 ( .A1(PermutationOutput2[52]), 
        .A2(Red_SubCellInst2_LFInst_13_LFInst_0_n14), .ZN(
        Red_SubCellInst2_LFInst_13_LFInst_0_n15) );
  NOR2_X1 Red_SubCellInst2_LFInst_13_LFInst_0_U1 ( .A1(PermutationOutput2[55]), 
        .A2(PermutationOutput2[53]), .ZN(
        Red_SubCellInst2_LFInst_13_LFInst_0_n14) );
  NAND2_X1 Red_SubCellInst2_LFInst_14_LFInst_0_U7 ( .A1(
        Red_SubCellInst2_LFInst_14_LFInst_0_n17), .A2(
        Red_SubCellInst2_LFInst_14_LFInst_0_n21), .ZN(Red_Feedback[14]) );
  NAND2_X1 Red_SubCellInst2_LFInst_14_LFInst_0_U6 ( .A1(
        Red_SubCellInst2_LFInst_14_LFInst_0_n20), .A2(
        Red_SubCellInst2_LFInst_14_LFInst_0_n16), .ZN(
        Red_SubCellInst2_LFInst_14_LFInst_0_n21) );
  XOR2_X1 Red_SubCellInst2_LFInst_14_LFInst_0_U5 ( .A(PermutationOutput2[58]), 
        .B(Red_SubCellInst2_LFInst_14_LFInst_0_n19), .Z(
        Red_SubCellInst2_LFInst_14_LFInst_0_n20) );
  NOR2_X1 Red_SubCellInst2_LFInst_14_LFInst_0_U4 ( .A1(PermutationOutput2[56]), 
        .A2(Red_SubCellInst2_LFInst_14_LFInst_0_n18), .ZN(
        Red_SubCellInst2_LFInst_14_LFInst_0_n19) );
  NOR2_X1 Red_SubCellInst2_LFInst_14_LFInst_0_U3 ( .A1(PermutationOutput2[59]), 
        .A2(PermutationOutput2[57]), .ZN(
        Red_SubCellInst2_LFInst_14_LFInst_0_n18) );
  OR2_X1 Red_SubCellInst2_LFInst_14_LFInst_0_U2 ( .A1(PermutationOutput2[56]), 
        .A2(Red_SubCellInst2_LFInst_14_LFInst_0_n16), .ZN(
        Red_SubCellInst2_LFInst_14_LFInst_0_n17) );
  NAND2_X1 Red_SubCellInst2_LFInst_14_LFInst_0_U1 ( .A1(PermutationOutput2[59]), .A2(PermutationOutput2[57]), .ZN(Red_SubCellInst2_LFInst_14_LFInst_0_n16) );
  NAND2_X1 Red_SubCellInst2_LFInst_15_LFInst_0_U7 ( .A1(
        Red_SubCellInst2_LFInst_15_LFInst_0_n17), .A2(
        Red_SubCellInst2_LFInst_15_LFInst_0_n21), .ZN(Red_Feedback[15]) );
  NAND2_X1 Red_SubCellInst2_LFInst_15_LFInst_0_U6 ( .A1(
        Red_SubCellInst2_LFInst_15_LFInst_0_n20), .A2(
        Red_SubCellInst2_LFInst_15_LFInst_0_n16), .ZN(
        Red_SubCellInst2_LFInst_15_LFInst_0_n21) );
  XOR2_X1 Red_SubCellInst2_LFInst_15_LFInst_0_U5 ( .A(PermutationOutput2[62]), 
        .B(Red_SubCellInst2_LFInst_15_LFInst_0_n19), .Z(
        Red_SubCellInst2_LFInst_15_LFInst_0_n20) );
  NOR2_X1 Red_SubCellInst2_LFInst_15_LFInst_0_U4 ( .A1(PermutationOutput2[60]), 
        .A2(Red_SubCellInst2_LFInst_15_LFInst_0_n18), .ZN(
        Red_SubCellInst2_LFInst_15_LFInst_0_n19) );
  NOR2_X1 Red_SubCellInst2_LFInst_15_LFInst_0_U3 ( .A1(PermutationOutput2[63]), 
        .A2(PermutationOutput2[61]), .ZN(
        Red_SubCellInst2_LFInst_15_LFInst_0_n18) );
  OR2_X1 Red_SubCellInst2_LFInst_15_LFInst_0_U2 ( .A1(PermutationOutput2[60]), 
        .A2(Red_SubCellInst2_LFInst_15_LFInst_0_n16), .ZN(
        Red_SubCellInst2_LFInst_15_LFInst_0_n17) );
  NAND2_X1 Red_SubCellInst2_LFInst_15_LFInst_0_U1 ( .A1(PermutationOutput2[63]), .A2(PermutationOutput2[61]), .ZN(Red_SubCellInst2_LFInst_15_LFInst_0_n16) );
  XNOR2_X1 Red_K0Inst_LFInst_0_LFInst_0_U3 ( .A(
        Red_K0Inst_LFInst_0_LFInst_0_n6), .B(Red_K0Inst_LFInst_0_LFInst_0_n5), 
        .ZN(Red_K0[0]) );
  XNOR2_X1 Red_K0Inst_LFInst_0_LFInst_0_U2 ( .A(Key[66]), .B(Key[67]), .ZN(
        Red_K0Inst_LFInst_0_LFInst_0_n5) );
  XOR2_X1 Red_K0Inst_LFInst_0_LFInst_0_U1 ( .A(Key[64]), .B(Key[65]), .Z(
        Red_K0Inst_LFInst_0_LFInst_0_n6) );
  XNOR2_X1 Red_K0Inst_LFInst_1_LFInst_0_U3 ( .A(
        Red_K0Inst_LFInst_1_LFInst_0_n6), .B(Red_K0Inst_LFInst_1_LFInst_0_n5), 
        .ZN(Red_K0[1]) );
  XNOR2_X1 Red_K0Inst_LFInst_1_LFInst_0_U2 ( .A(Key[70]), .B(Key[71]), .ZN(
        Red_K0Inst_LFInst_1_LFInst_0_n5) );
  XOR2_X1 Red_K0Inst_LFInst_1_LFInst_0_U1 ( .A(Key[68]), .B(Key[69]), .Z(
        Red_K0Inst_LFInst_1_LFInst_0_n6) );
  XNOR2_X1 Red_K0Inst_LFInst_2_LFInst_0_U3 ( .A(
        Red_K0Inst_LFInst_2_LFInst_0_n6), .B(Red_K0Inst_LFInst_2_LFInst_0_n5), 
        .ZN(Red_K0[2]) );
  XNOR2_X1 Red_K0Inst_LFInst_2_LFInst_0_U2 ( .A(Key[74]), .B(Key[75]), .ZN(
        Red_K0Inst_LFInst_2_LFInst_0_n5) );
  XOR2_X1 Red_K0Inst_LFInst_2_LFInst_0_U1 ( .A(Key[72]), .B(Key[73]), .Z(
        Red_K0Inst_LFInst_2_LFInst_0_n6) );
  XNOR2_X1 Red_K0Inst_LFInst_3_LFInst_0_U3 ( .A(
        Red_K0Inst_LFInst_3_LFInst_0_n6), .B(Red_K0Inst_LFInst_3_LFInst_0_n5), 
        .ZN(Red_K0[3]) );
  XNOR2_X1 Red_K0Inst_LFInst_3_LFInst_0_U2 ( .A(Key[78]), .B(Key[79]), .ZN(
        Red_K0Inst_LFInst_3_LFInst_0_n5) );
  XOR2_X1 Red_K0Inst_LFInst_3_LFInst_0_U1 ( .A(Key[76]), .B(Key[77]), .Z(
        Red_K0Inst_LFInst_3_LFInst_0_n6) );
  XNOR2_X1 Red_K0Inst_LFInst_4_LFInst_0_U3 ( .A(
        Red_K0Inst_LFInst_4_LFInst_0_n6), .B(Red_K0Inst_LFInst_4_LFInst_0_n5), 
        .ZN(Red_K0[4]) );
  XNOR2_X1 Red_K0Inst_LFInst_4_LFInst_0_U2 ( .A(Key[82]), .B(Key[83]), .ZN(
        Red_K0Inst_LFInst_4_LFInst_0_n5) );
  XOR2_X1 Red_K0Inst_LFInst_4_LFInst_0_U1 ( .A(Key[80]), .B(Key[81]), .Z(
        Red_K0Inst_LFInst_4_LFInst_0_n6) );
  XNOR2_X1 Red_K0Inst_LFInst_5_LFInst_0_U3 ( .A(
        Red_K0Inst_LFInst_5_LFInst_0_n6), .B(Red_K0Inst_LFInst_5_LFInst_0_n5), 
        .ZN(Red_K0[5]) );
  XNOR2_X1 Red_K0Inst_LFInst_5_LFInst_0_U2 ( .A(Key[86]), .B(Key[87]), .ZN(
        Red_K0Inst_LFInst_5_LFInst_0_n5) );
  XOR2_X1 Red_K0Inst_LFInst_5_LFInst_0_U1 ( .A(Key[84]), .B(Key[85]), .Z(
        Red_K0Inst_LFInst_5_LFInst_0_n6) );
  XNOR2_X1 Red_K0Inst_LFInst_6_LFInst_0_U3 ( .A(
        Red_K0Inst_LFInst_6_LFInst_0_n6), .B(Red_K0Inst_LFInst_6_LFInst_0_n5), 
        .ZN(Red_K0[6]) );
  XNOR2_X1 Red_K0Inst_LFInst_6_LFInst_0_U2 ( .A(Key[90]), .B(Key[91]), .ZN(
        Red_K0Inst_LFInst_6_LFInst_0_n5) );
  XOR2_X1 Red_K0Inst_LFInst_6_LFInst_0_U1 ( .A(Key[88]), .B(Key[89]), .Z(
        Red_K0Inst_LFInst_6_LFInst_0_n6) );
  XNOR2_X1 Red_K0Inst_LFInst_7_LFInst_0_U3 ( .A(
        Red_K0Inst_LFInst_7_LFInst_0_n6), .B(Red_K0Inst_LFInst_7_LFInst_0_n5), 
        .ZN(Red_K0[7]) );
  XNOR2_X1 Red_K0Inst_LFInst_7_LFInst_0_U2 ( .A(Key[94]), .B(Key[95]), .ZN(
        Red_K0Inst_LFInst_7_LFInst_0_n5) );
  XOR2_X1 Red_K0Inst_LFInst_7_LFInst_0_U1 ( .A(Key[92]), .B(Key[93]), .Z(
        Red_K0Inst_LFInst_7_LFInst_0_n6) );
  XNOR2_X1 Red_K0Inst_LFInst_8_LFInst_0_U3 ( .A(
        Red_K0Inst_LFInst_8_LFInst_0_n6), .B(Red_K0Inst_LFInst_8_LFInst_0_n5), 
        .ZN(Red_K0[8]) );
  XNOR2_X1 Red_K0Inst_LFInst_8_LFInst_0_U2 ( .A(Key[98]), .B(Key[99]), .ZN(
        Red_K0Inst_LFInst_8_LFInst_0_n5) );
  XOR2_X1 Red_K0Inst_LFInst_8_LFInst_0_U1 ( .A(Key[96]), .B(Key[97]), .Z(
        Red_K0Inst_LFInst_8_LFInst_0_n6) );
  XNOR2_X1 Red_K0Inst_LFInst_9_LFInst_0_U3 ( .A(
        Red_K0Inst_LFInst_9_LFInst_0_n6), .B(Red_K0Inst_LFInst_9_LFInst_0_n5), 
        .ZN(Red_K0[9]) );
  XNOR2_X1 Red_K0Inst_LFInst_9_LFInst_0_U2 ( .A(Key[102]), .B(Key[103]), .ZN(
        Red_K0Inst_LFInst_9_LFInst_0_n5) );
  XOR2_X1 Red_K0Inst_LFInst_9_LFInst_0_U1 ( .A(Key[100]), .B(Key[101]), .Z(
        Red_K0Inst_LFInst_9_LFInst_0_n6) );
  XNOR2_X1 Red_K0Inst_LFInst_10_LFInst_0_U3 ( .A(
        Red_K0Inst_LFInst_10_LFInst_0_n6), .B(Red_K0Inst_LFInst_10_LFInst_0_n5), .ZN(Red_K0[10]) );
  XNOR2_X1 Red_K0Inst_LFInst_10_LFInst_0_U2 ( .A(Key[106]), .B(Key[107]), .ZN(
        Red_K0Inst_LFInst_10_LFInst_0_n5) );
  XOR2_X1 Red_K0Inst_LFInst_10_LFInst_0_U1 ( .A(Key[104]), .B(Key[105]), .Z(
        Red_K0Inst_LFInst_10_LFInst_0_n6) );
  XNOR2_X1 Red_K0Inst_LFInst_11_LFInst_0_U3 ( .A(
        Red_K0Inst_LFInst_11_LFInst_0_n6), .B(Red_K0Inst_LFInst_11_LFInst_0_n5), .ZN(Red_K0[11]) );
  XNOR2_X1 Red_K0Inst_LFInst_11_LFInst_0_U2 ( .A(Key[110]), .B(Key[111]), .ZN(
        Red_K0Inst_LFInst_11_LFInst_0_n5) );
  XOR2_X1 Red_K0Inst_LFInst_11_LFInst_0_U1 ( .A(Key[108]), .B(Key[109]), .Z(
        Red_K0Inst_LFInst_11_LFInst_0_n6) );
  XNOR2_X1 Red_K0Inst_LFInst_12_LFInst_0_U3 ( .A(
        Red_K0Inst_LFInst_12_LFInst_0_n6), .B(Red_K0Inst_LFInst_12_LFInst_0_n5), .ZN(Red_K0[12]) );
  XNOR2_X1 Red_K0Inst_LFInst_12_LFInst_0_U2 ( .A(Key[114]), .B(Key[115]), .ZN(
        Red_K0Inst_LFInst_12_LFInst_0_n5) );
  XOR2_X1 Red_K0Inst_LFInst_12_LFInst_0_U1 ( .A(Key[112]), .B(Key[113]), .Z(
        Red_K0Inst_LFInst_12_LFInst_0_n6) );
  XNOR2_X1 Red_K0Inst_LFInst_13_LFInst_0_U3 ( .A(
        Red_K0Inst_LFInst_13_LFInst_0_n6), .B(Red_K0Inst_LFInst_13_LFInst_0_n5), .ZN(Red_K0[13]) );
  XNOR2_X1 Red_K0Inst_LFInst_13_LFInst_0_U2 ( .A(Key[118]), .B(Key[119]), .ZN(
        Red_K0Inst_LFInst_13_LFInst_0_n5) );
  XOR2_X1 Red_K0Inst_LFInst_13_LFInst_0_U1 ( .A(Key[116]), .B(Key[117]), .Z(
        Red_K0Inst_LFInst_13_LFInst_0_n6) );
  XNOR2_X1 Red_K0Inst_LFInst_14_LFInst_0_U3 ( .A(
        Red_K0Inst_LFInst_14_LFInst_0_n6), .B(Red_K0Inst_LFInst_14_LFInst_0_n5), .ZN(Red_K0[14]) );
  XNOR2_X1 Red_K0Inst_LFInst_14_LFInst_0_U2 ( .A(Key[122]), .B(Key[123]), .ZN(
        Red_K0Inst_LFInst_14_LFInst_0_n5) );
  XOR2_X1 Red_K0Inst_LFInst_14_LFInst_0_U1 ( .A(Key[120]), .B(Key[121]), .Z(
        Red_K0Inst_LFInst_14_LFInst_0_n6) );
  XNOR2_X1 Red_K0Inst_LFInst_15_LFInst_0_U3 ( .A(
        Red_K0Inst_LFInst_15_LFInst_0_n6), .B(Red_K0Inst_LFInst_15_LFInst_0_n5), .ZN(Red_K0[15]) );
  XNOR2_X1 Red_K0Inst_LFInst_15_LFInst_0_U2 ( .A(Key[126]), .B(Key[127]), .ZN(
        Red_K0Inst_LFInst_15_LFInst_0_n5) );
  XOR2_X1 Red_K0Inst_LFInst_15_LFInst_0_U1 ( .A(Key[124]), .B(Key[125]), .Z(
        Red_K0Inst_LFInst_15_LFInst_0_n6) );
  XNOR2_X1 Red_K1Inst_LFInst_0_LFInst_0_U3 ( .A(
        Red_K1Inst_LFInst_0_LFInst_0_n6), .B(Red_K1Inst_LFInst_0_LFInst_0_n5), 
        .ZN(Red_K1[0]) );
  XNOR2_X1 Red_K1Inst_LFInst_0_LFInst_0_U2 ( .A(Key[2]), .B(Key[3]), .ZN(
        Red_K1Inst_LFInst_0_LFInst_0_n5) );
  XOR2_X1 Red_K1Inst_LFInst_0_LFInst_0_U1 ( .A(Key[0]), .B(Key[1]), .Z(
        Red_K1Inst_LFInst_0_LFInst_0_n6) );
  XNOR2_X1 Red_K1Inst_LFInst_1_LFInst_0_U3 ( .A(
        Red_K1Inst_LFInst_1_LFInst_0_n6), .B(Red_K1Inst_LFInst_1_LFInst_0_n5), 
        .ZN(Red_K1[1]) );
  XNOR2_X1 Red_K1Inst_LFInst_1_LFInst_0_U2 ( .A(Key[6]), .B(Key[7]), .ZN(
        Red_K1Inst_LFInst_1_LFInst_0_n5) );
  XOR2_X1 Red_K1Inst_LFInst_1_LFInst_0_U1 ( .A(Key[4]), .B(Key[5]), .Z(
        Red_K1Inst_LFInst_1_LFInst_0_n6) );
  XNOR2_X1 Red_K1Inst_LFInst_2_LFInst_0_U3 ( .A(
        Red_K1Inst_LFInst_2_LFInst_0_n6), .B(Red_K1Inst_LFInst_2_LFInst_0_n5), 
        .ZN(Red_K1[2]) );
  XNOR2_X1 Red_K1Inst_LFInst_2_LFInst_0_U2 ( .A(Key[10]), .B(Key[11]), .ZN(
        Red_K1Inst_LFInst_2_LFInst_0_n5) );
  XOR2_X1 Red_K1Inst_LFInst_2_LFInst_0_U1 ( .A(Key[8]), .B(Key[9]), .Z(
        Red_K1Inst_LFInst_2_LFInst_0_n6) );
  XNOR2_X1 Red_K1Inst_LFInst_3_LFInst_0_U3 ( .A(
        Red_K1Inst_LFInst_3_LFInst_0_n6), .B(Red_K1Inst_LFInst_3_LFInst_0_n5), 
        .ZN(Red_K1[3]) );
  XNOR2_X1 Red_K1Inst_LFInst_3_LFInst_0_U2 ( .A(Key[14]), .B(Key[15]), .ZN(
        Red_K1Inst_LFInst_3_LFInst_0_n5) );
  XOR2_X1 Red_K1Inst_LFInst_3_LFInst_0_U1 ( .A(Key[12]), .B(Key[13]), .Z(
        Red_K1Inst_LFInst_3_LFInst_0_n6) );
  XNOR2_X1 Red_K1Inst_LFInst_4_LFInst_0_U3 ( .A(
        Red_K1Inst_LFInst_4_LFInst_0_n6), .B(Red_K1Inst_LFInst_4_LFInst_0_n5), 
        .ZN(Red_K1[4]) );
  XNOR2_X1 Red_K1Inst_LFInst_4_LFInst_0_U2 ( .A(Key[18]), .B(Key[19]), .ZN(
        Red_K1Inst_LFInst_4_LFInst_0_n5) );
  XOR2_X1 Red_K1Inst_LFInst_4_LFInst_0_U1 ( .A(Key[16]), .B(Key[17]), .Z(
        Red_K1Inst_LFInst_4_LFInst_0_n6) );
  XNOR2_X1 Red_K1Inst_LFInst_5_LFInst_0_U3 ( .A(
        Red_K1Inst_LFInst_5_LFInst_0_n6), .B(Red_K1Inst_LFInst_5_LFInst_0_n5), 
        .ZN(Red_K1[5]) );
  XNOR2_X1 Red_K1Inst_LFInst_5_LFInst_0_U2 ( .A(Key[22]), .B(Key[23]), .ZN(
        Red_K1Inst_LFInst_5_LFInst_0_n5) );
  XOR2_X1 Red_K1Inst_LFInst_5_LFInst_0_U1 ( .A(Key[20]), .B(Key[21]), .Z(
        Red_K1Inst_LFInst_5_LFInst_0_n6) );
  XNOR2_X1 Red_K1Inst_LFInst_6_LFInst_0_U3 ( .A(
        Red_K1Inst_LFInst_6_LFInst_0_n6), .B(Red_K1Inst_LFInst_6_LFInst_0_n5), 
        .ZN(Red_K1[6]) );
  XNOR2_X1 Red_K1Inst_LFInst_6_LFInst_0_U2 ( .A(Key[26]), .B(Key[27]), .ZN(
        Red_K1Inst_LFInst_6_LFInst_0_n5) );
  XOR2_X1 Red_K1Inst_LFInst_6_LFInst_0_U1 ( .A(Key[24]), .B(Key[25]), .Z(
        Red_K1Inst_LFInst_6_LFInst_0_n6) );
  XNOR2_X1 Red_K1Inst_LFInst_7_LFInst_0_U3 ( .A(
        Red_K1Inst_LFInst_7_LFInst_0_n6), .B(Red_K1Inst_LFInst_7_LFInst_0_n5), 
        .ZN(Red_K1[7]) );
  XNOR2_X1 Red_K1Inst_LFInst_7_LFInst_0_U2 ( .A(Key[30]), .B(Key[31]), .ZN(
        Red_K1Inst_LFInst_7_LFInst_0_n5) );
  XOR2_X1 Red_K1Inst_LFInst_7_LFInst_0_U1 ( .A(Key[28]), .B(Key[29]), .Z(
        Red_K1Inst_LFInst_7_LFInst_0_n6) );
  XNOR2_X1 Red_K1Inst_LFInst_8_LFInst_0_U3 ( .A(
        Red_K1Inst_LFInst_8_LFInst_0_n6), .B(Red_K1Inst_LFInst_8_LFInst_0_n5), 
        .ZN(Red_K1[8]) );
  XNOR2_X1 Red_K1Inst_LFInst_8_LFInst_0_U2 ( .A(Key[34]), .B(Key[35]), .ZN(
        Red_K1Inst_LFInst_8_LFInst_0_n5) );
  XOR2_X1 Red_K1Inst_LFInst_8_LFInst_0_U1 ( .A(Key[32]), .B(Key[33]), .Z(
        Red_K1Inst_LFInst_8_LFInst_0_n6) );
  XNOR2_X1 Red_K1Inst_LFInst_9_LFInst_0_U3 ( .A(
        Red_K1Inst_LFInst_9_LFInst_0_n6), .B(Red_K1Inst_LFInst_9_LFInst_0_n5), 
        .ZN(Red_K1[9]) );
  XNOR2_X1 Red_K1Inst_LFInst_9_LFInst_0_U2 ( .A(Key[38]), .B(Key[39]), .ZN(
        Red_K1Inst_LFInst_9_LFInst_0_n5) );
  XOR2_X1 Red_K1Inst_LFInst_9_LFInst_0_U1 ( .A(Key[36]), .B(Key[37]), .Z(
        Red_K1Inst_LFInst_9_LFInst_0_n6) );
  XNOR2_X1 Red_K1Inst_LFInst_10_LFInst_0_U3 ( .A(
        Red_K1Inst_LFInst_10_LFInst_0_n6), .B(Red_K1Inst_LFInst_10_LFInst_0_n5), .ZN(Red_K1[10]) );
  XNOR2_X1 Red_K1Inst_LFInst_10_LFInst_0_U2 ( .A(Key[42]), .B(Key[43]), .ZN(
        Red_K1Inst_LFInst_10_LFInst_0_n5) );
  XOR2_X1 Red_K1Inst_LFInst_10_LFInst_0_U1 ( .A(Key[40]), .B(Key[41]), .Z(
        Red_K1Inst_LFInst_10_LFInst_0_n6) );
  XNOR2_X1 Red_K1Inst_LFInst_11_LFInst_0_U3 ( .A(
        Red_K1Inst_LFInst_11_LFInst_0_n6), .B(Red_K1Inst_LFInst_11_LFInst_0_n5), .ZN(Red_K1[11]) );
  XNOR2_X1 Red_K1Inst_LFInst_11_LFInst_0_U2 ( .A(Key[46]), .B(Key[47]), .ZN(
        Red_K1Inst_LFInst_11_LFInst_0_n5) );
  XOR2_X1 Red_K1Inst_LFInst_11_LFInst_0_U1 ( .A(Key[44]), .B(Key[45]), .Z(
        Red_K1Inst_LFInst_11_LFInst_0_n6) );
  XNOR2_X1 Red_K1Inst_LFInst_12_LFInst_0_U3 ( .A(
        Red_K1Inst_LFInst_12_LFInst_0_n6), .B(Red_K1Inst_LFInst_12_LFInst_0_n5), .ZN(Red_K1[12]) );
  XNOR2_X1 Red_K1Inst_LFInst_12_LFInst_0_U2 ( .A(Key[50]), .B(Key[51]), .ZN(
        Red_K1Inst_LFInst_12_LFInst_0_n5) );
  XOR2_X1 Red_K1Inst_LFInst_12_LFInst_0_U1 ( .A(Key[48]), .B(Key[49]), .Z(
        Red_K1Inst_LFInst_12_LFInst_0_n6) );
  XNOR2_X1 Red_K1Inst_LFInst_13_LFInst_0_U3 ( .A(
        Red_K1Inst_LFInst_13_LFInst_0_n6), .B(Red_K1Inst_LFInst_13_LFInst_0_n5), .ZN(Red_K1[13]) );
  XNOR2_X1 Red_K1Inst_LFInst_13_LFInst_0_U2 ( .A(Key[54]), .B(Key[55]), .ZN(
        Red_K1Inst_LFInst_13_LFInst_0_n5) );
  XOR2_X1 Red_K1Inst_LFInst_13_LFInst_0_U1 ( .A(Key[52]), .B(Key[53]), .Z(
        Red_K1Inst_LFInst_13_LFInst_0_n6) );
  XNOR2_X1 Red_K1Inst_LFInst_14_LFInst_0_U3 ( .A(
        Red_K1Inst_LFInst_14_LFInst_0_n6), .B(Red_K1Inst_LFInst_14_LFInst_0_n5), .ZN(Red_K1[14]) );
  XNOR2_X1 Red_K1Inst_LFInst_14_LFInst_0_U2 ( .A(Key[58]), .B(Key[59]), .ZN(
        Red_K1Inst_LFInst_14_LFInst_0_n5) );
  XOR2_X1 Red_K1Inst_LFInst_14_LFInst_0_U1 ( .A(Key[56]), .B(Key[57]), .Z(
        Red_K1Inst_LFInst_14_LFInst_0_n6) );
  XNOR2_X1 Red_K1Inst_LFInst_15_LFInst_0_U3 ( .A(
        Red_K1Inst_LFInst_15_LFInst_0_n6), .B(Red_K1Inst_LFInst_15_LFInst_0_n5), .ZN(Red_K1[15]) );
  XNOR2_X1 Red_K1Inst_LFInst_15_LFInst_0_U2 ( .A(Key[62]), .B(Key[63]), .ZN(
        Red_K1Inst_LFInst_15_LFInst_0_n5) );
  XOR2_X1 Red_K1Inst_LFInst_15_LFInst_0_U1 ( .A(Key[60]), .B(Key[61]), .Z(
        Red_K1Inst_LFInst_15_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_0_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_0_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_0_LFInst_0_n5), .ZN(Red_SignaltoCheck[0]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_0_LFInst_0_U2 ( .A(AddRoundKeyOutput2[2]), 
        .B(AddRoundKeyOutput2[3]), .ZN(Red_ToCheckInst_LFInst_0_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_0_LFInst_0_U1 ( .A(AddRoundKeyOutput2[0]), 
        .B(AddRoundKeyOutput2[1]), .Z(Red_ToCheckInst_LFInst_0_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_1_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_1_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_1_LFInst_0_n5), .ZN(Red_SignaltoCheck[1]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_1_LFInst_0_U2 ( .A(AddRoundKeyOutput2[6]), 
        .B(AddRoundKeyOutput2[7]), .ZN(Red_ToCheckInst_LFInst_1_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_1_LFInst_0_U1 ( .A(AddRoundKeyOutput2[4]), 
        .B(AddRoundKeyOutput2[5]), .Z(Red_ToCheckInst_LFInst_1_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_2_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_2_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_2_LFInst_0_n5), .ZN(Red_SignaltoCheck[2]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_2_LFInst_0_U2 ( .A(AddRoundKeyOutput2[10]), 
        .B(AddRoundKeyOutput2[11]), .ZN(Red_ToCheckInst_LFInst_2_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_2_LFInst_0_U1 ( .A(AddRoundKeyOutput2[8]), 
        .B(AddRoundKeyOutput2[9]), .Z(Red_ToCheckInst_LFInst_2_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_3_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_3_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_3_LFInst_0_n5), .ZN(Red_SignaltoCheck[3]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_3_LFInst_0_U2 ( .A(AddRoundKeyOutput2[14]), 
        .B(AddRoundKeyOutput2[15]), .ZN(Red_ToCheckInst_LFInst_3_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_3_LFInst_0_U1 ( .A(AddRoundKeyOutput2[12]), 
        .B(AddRoundKeyOutput2[13]), .Z(Red_ToCheckInst_LFInst_3_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_4_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_4_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_4_LFInst_0_n5), .ZN(Red_SignaltoCheck[4]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_4_LFInst_0_U2 ( .A(AddRoundKeyOutput2[18]), 
        .B(AddRoundKeyOutput2[19]), .ZN(Red_ToCheckInst_LFInst_4_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_4_LFInst_0_U1 ( .A(AddRoundKeyOutput2[16]), 
        .B(AddRoundKeyOutput2[17]), .Z(Red_ToCheckInst_LFInst_4_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_5_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_5_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_5_LFInst_0_n5), .ZN(Red_SignaltoCheck[5]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_5_LFInst_0_U2 ( .A(AddRoundKeyOutput2[22]), 
        .B(AddRoundKeyOutput2[23]), .ZN(Red_ToCheckInst_LFInst_5_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_5_LFInst_0_U1 ( .A(AddRoundKeyOutput2[20]), 
        .B(AddRoundKeyOutput2[21]), .Z(Red_ToCheckInst_LFInst_5_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_6_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_6_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_6_LFInst_0_n5), .ZN(Red_SignaltoCheck[6]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_6_LFInst_0_U2 ( .A(AddRoundKeyOutput2[26]), 
        .B(AddRoundKeyOutput2[27]), .ZN(Red_ToCheckInst_LFInst_6_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_6_LFInst_0_U1 ( .A(AddRoundKeyOutput2[24]), 
        .B(AddRoundKeyOutput2[25]), .Z(Red_ToCheckInst_LFInst_6_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_7_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_7_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_7_LFInst_0_n5), .ZN(Red_SignaltoCheck[7]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_7_LFInst_0_U2 ( .A(AddRoundKeyOutput2[30]), 
        .B(AddRoundKeyOutput2[31]), .ZN(Red_ToCheckInst_LFInst_7_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_7_LFInst_0_U1 ( .A(AddRoundKeyOutput2[28]), 
        .B(AddRoundKeyOutput2[29]), .Z(Red_ToCheckInst_LFInst_7_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_8_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_8_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_8_LFInst_0_n5), .ZN(Red_SignaltoCheck[8]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_8_LFInst_0_U2 ( .A(AddRoundKeyOutput2[34]), 
        .B(AddRoundKeyOutput2[35]), .ZN(Red_ToCheckInst_LFInst_8_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_8_LFInst_0_U1 ( .A(AddRoundKeyOutput2[32]), 
        .B(AddRoundKeyOutput2[33]), .Z(Red_ToCheckInst_LFInst_8_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_9_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_9_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_9_LFInst_0_n5), .ZN(Red_SignaltoCheck[9]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_9_LFInst_0_U2 ( .A(AddRoundKeyOutput2[38]), 
        .B(AddRoundKeyOutput2[39]), .ZN(Red_ToCheckInst_LFInst_9_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_9_LFInst_0_U1 ( .A(AddRoundKeyOutput2[36]), 
        .B(AddRoundKeyOutput2[37]), .Z(Red_ToCheckInst_LFInst_9_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_10_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_10_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_10_LFInst_0_n5), .ZN(Red_SignaltoCheck[10]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_10_LFInst_0_U2 ( .A(AddRoundKeyOutput2[42]), 
        .B(AddRoundKeyOutput2[43]), .ZN(Red_ToCheckInst_LFInst_10_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_10_LFInst_0_U1 ( .A(AddRoundKeyOutput2[40]), 
        .B(AddRoundKeyOutput2[41]), .Z(Red_ToCheckInst_LFInst_10_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_11_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_11_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_11_LFInst_0_n5), .ZN(Red_SignaltoCheck[11]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_11_LFInst_0_U2 ( .A(AddRoundKeyOutput2[46]), 
        .B(AddRoundKeyOutput2[47]), .ZN(Red_ToCheckInst_LFInst_11_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_11_LFInst_0_U1 ( .A(AddRoundKeyOutput2[44]), 
        .B(AddRoundKeyOutput2[45]), .Z(Red_ToCheckInst_LFInst_11_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_12_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_12_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_12_LFInst_0_n5), .ZN(Red_SignaltoCheck[12]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_12_LFInst_0_U2 ( .A(AddRoundKeyOutput2[50]), 
        .B(AddRoundKeyOutput2[51]), .ZN(Red_ToCheckInst_LFInst_12_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_12_LFInst_0_U1 ( .A(AddRoundKeyOutput2[48]), 
        .B(AddRoundKeyOutput2[49]), .Z(Red_ToCheckInst_LFInst_12_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_13_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_13_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_13_LFInst_0_n5), .ZN(Red_SignaltoCheck[13]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_13_LFInst_0_U2 ( .A(AddRoundKeyOutput2[54]), 
        .B(AddRoundKeyOutput2[55]), .ZN(Red_ToCheckInst_LFInst_13_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_13_LFInst_0_U1 ( .A(AddRoundKeyOutput2[52]), 
        .B(AddRoundKeyOutput2[53]), .Z(Red_ToCheckInst_LFInst_13_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_14_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_14_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_14_LFInst_0_n5), .ZN(Red_SignaltoCheck[14]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_14_LFInst_0_U2 ( .A(AddRoundKeyOutput2[58]), 
        .B(AddRoundKeyOutput2[59]), .ZN(Red_ToCheckInst_LFInst_14_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_14_LFInst_0_U1 ( .A(AddRoundKeyOutput2[56]), 
        .B(AddRoundKeyOutput2[57]), .Z(Red_ToCheckInst_LFInst_14_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_15_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_15_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_15_LFInst_0_n5), .ZN(Red_SignaltoCheck[15]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_15_LFInst_0_U2 ( .A(AddRoundKeyOutput2[62]), 
        .B(AddRoundKeyOutput2[63]), .ZN(Red_ToCheckInst_LFInst_15_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_15_LFInst_0_U1 ( .A(AddRoundKeyOutput2[60]), 
        .B(AddRoundKeyOutput2[61]), .Z(Red_ToCheckInst_LFInst_15_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_16_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_16_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_16_LFInst_0_n5), .ZN(Red_SignaltoCheck[16]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_16_LFInst_0_U2 ( .A(AddRoundKeyOutput[2]), 
        .B(AddRoundKeyOutput[3]), .ZN(Red_ToCheckInst_LFInst_16_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_16_LFInst_0_U1 ( .A(AddRoundKeyOutput[0]), 
        .B(AddRoundKeyOutput[1]), .Z(Red_ToCheckInst_LFInst_16_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_17_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_17_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_17_LFInst_0_n5), .ZN(Red_SignaltoCheck[17]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_17_LFInst_0_U2 ( .A(AddRoundKeyOutput[6]), 
        .B(AddRoundKeyOutput[7]), .ZN(Red_ToCheckInst_LFInst_17_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_17_LFInst_0_U1 ( .A(AddRoundKeyOutput[4]), 
        .B(AddRoundKeyOutput[5]), .Z(Red_ToCheckInst_LFInst_17_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_18_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_18_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_18_LFInst_0_n5), .ZN(Red_SignaltoCheck[18]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_18_LFInst_0_U2 ( .A(AddRoundKeyOutput[10]), 
        .B(AddRoundKeyOutput[11]), .ZN(Red_ToCheckInst_LFInst_18_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_18_LFInst_0_U1 ( .A(AddRoundKeyOutput[8]), 
        .B(AddRoundKeyOutput[9]), .Z(Red_ToCheckInst_LFInst_18_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_19_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_19_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_19_LFInst_0_n5), .ZN(Red_SignaltoCheck[19]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_19_LFInst_0_U2 ( .A(AddRoundKeyOutput[14]), 
        .B(AddRoundKeyOutput[15]), .ZN(Red_ToCheckInst_LFInst_19_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_19_LFInst_0_U1 ( .A(AddRoundKeyOutput[12]), 
        .B(AddRoundKeyOutput[13]), .Z(Red_ToCheckInst_LFInst_19_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_20_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_20_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_20_LFInst_0_n5), .ZN(Red_SignaltoCheck[20]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_20_LFInst_0_U2 ( .A(AddRoundKeyOutput[18]), 
        .B(AddRoundKeyOutput[19]), .ZN(Red_ToCheckInst_LFInst_20_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_20_LFInst_0_U1 ( .A(AddRoundKeyOutput[16]), 
        .B(AddRoundKeyOutput[17]), .Z(Red_ToCheckInst_LFInst_20_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_21_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_21_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_21_LFInst_0_n5), .ZN(Red_SignaltoCheck[21]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_21_LFInst_0_U2 ( .A(AddRoundKeyOutput[22]), 
        .B(AddRoundKeyOutput[23]), .ZN(Red_ToCheckInst_LFInst_21_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_21_LFInst_0_U1 ( .A(AddRoundKeyOutput[20]), 
        .B(AddRoundKeyOutput[21]), .Z(Red_ToCheckInst_LFInst_21_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_22_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_22_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_22_LFInst_0_n5), .ZN(Red_SignaltoCheck[22]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_22_LFInst_0_U2 ( .A(AddRoundKeyOutput[26]), 
        .B(AddRoundKeyOutput[27]), .ZN(Red_ToCheckInst_LFInst_22_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_22_LFInst_0_U1 ( .A(AddRoundKeyOutput[24]), 
        .B(AddRoundKeyOutput[25]), .Z(Red_ToCheckInst_LFInst_22_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_23_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_23_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_23_LFInst_0_n5), .ZN(Red_SignaltoCheck[23]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_23_LFInst_0_U2 ( .A(AddRoundKeyOutput[30]), 
        .B(AddRoundKeyOutput[31]), .ZN(Red_ToCheckInst_LFInst_23_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_23_LFInst_0_U1 ( .A(AddRoundKeyOutput[28]), 
        .B(AddRoundKeyOutput[29]), .Z(Red_ToCheckInst_LFInst_23_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_24_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_24_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_24_LFInst_0_n5), .ZN(Red_SignaltoCheck[24]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_24_LFInst_0_U2 ( .A(AddRoundKeyOutput[34]), 
        .B(AddRoundKeyOutput[35]), .ZN(Red_ToCheckInst_LFInst_24_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_24_LFInst_0_U1 ( .A(AddRoundKeyOutput[32]), 
        .B(AddRoundKeyOutput[33]), .Z(Red_ToCheckInst_LFInst_24_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_25_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_25_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_25_LFInst_0_n5), .ZN(Red_SignaltoCheck[25]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_25_LFInst_0_U2 ( .A(AddRoundKeyOutput[38]), 
        .B(AddRoundKeyOutput[39]), .ZN(Red_ToCheckInst_LFInst_25_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_25_LFInst_0_U1 ( .A(AddRoundKeyOutput[36]), 
        .B(AddRoundKeyOutput[37]), .Z(Red_ToCheckInst_LFInst_25_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_26_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_26_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_26_LFInst_0_n5), .ZN(Red_SignaltoCheck[26]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_26_LFInst_0_U2 ( .A(AddRoundKeyOutput[42]), 
        .B(AddRoundKeyOutput[43]), .ZN(Red_ToCheckInst_LFInst_26_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_26_LFInst_0_U1 ( .A(AddRoundKeyOutput[40]), 
        .B(AddRoundKeyOutput[41]), .Z(Red_ToCheckInst_LFInst_26_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_27_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_27_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_27_LFInst_0_n5), .ZN(Red_SignaltoCheck[27]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_27_LFInst_0_U2 ( .A(AddRoundKeyOutput[46]), 
        .B(AddRoundKeyOutput[47]), .ZN(Red_ToCheckInst_LFInst_27_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_27_LFInst_0_U1 ( .A(AddRoundKeyOutput[44]), 
        .B(AddRoundKeyOutput[45]), .Z(Red_ToCheckInst_LFInst_27_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_28_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_28_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_28_LFInst_0_n5), .ZN(Red_SignaltoCheck[28]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_28_LFInst_0_U2 ( .A(AddRoundKeyOutput[50]), 
        .B(AddRoundKeyOutput[51]), .ZN(Red_ToCheckInst_LFInst_28_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_28_LFInst_0_U1 ( .A(AddRoundKeyOutput[48]), 
        .B(AddRoundKeyOutput[49]), .Z(Red_ToCheckInst_LFInst_28_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_29_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_29_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_29_LFInst_0_n5), .ZN(Red_SignaltoCheck[29]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_29_LFInst_0_U2 ( .A(AddRoundKeyOutput[54]), 
        .B(AddRoundKeyOutput[55]), .ZN(Red_ToCheckInst_LFInst_29_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_29_LFInst_0_U1 ( .A(AddRoundKeyOutput[52]), 
        .B(AddRoundKeyOutput[53]), .Z(Red_ToCheckInst_LFInst_29_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_30_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_30_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_30_LFInst_0_n5), .ZN(Red_SignaltoCheck[30]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_30_LFInst_0_U2 ( .A(AddRoundKeyOutput[58]), 
        .B(AddRoundKeyOutput[59]), .ZN(Red_ToCheckInst_LFInst_30_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_30_LFInst_0_U1 ( .A(AddRoundKeyOutput[56]), 
        .B(AddRoundKeyOutput[57]), .Z(Red_ToCheckInst_LFInst_30_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_31_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_31_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_31_LFInst_0_n5), .ZN(Red_SignaltoCheck[31]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_31_LFInst_0_U2 ( .A(AddRoundKeyOutput[62]), 
        .B(AddRoundKeyOutput[63]), .ZN(Red_ToCheckInst_LFInst_31_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_31_LFInst_0_U1 ( .A(AddRoundKeyOutput[60]), 
        .B(AddRoundKeyOutput[61]), .Z(Red_ToCheckInst_LFInst_31_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_32_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_32_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_32_LFInst_0_n5), .ZN(Red_SignaltoCheck[32]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_32_LFInst_0_U2 ( .A(Output[2]), .B(Output[3]), .ZN(Red_ToCheckInst_LFInst_32_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_32_LFInst_0_U1 ( .A(Output[0]), .B(Output[1]), 
        .Z(Red_ToCheckInst_LFInst_32_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_33_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_33_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_33_LFInst_0_n5), .ZN(Red_SignaltoCheck[33]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_33_LFInst_0_U2 ( .A(Output[6]), .B(Output[7]), .ZN(Red_ToCheckInst_LFInst_33_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_33_LFInst_0_U1 ( .A(Output[4]), .B(Output[5]), 
        .Z(Red_ToCheckInst_LFInst_33_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_34_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_34_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_34_LFInst_0_n5), .ZN(Red_SignaltoCheck[34]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_34_LFInst_0_U2 ( .A(Output[10]), .B(
        Output[11]), .ZN(Red_ToCheckInst_LFInst_34_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_34_LFInst_0_U1 ( .A(Output[8]), .B(Output[9]), 
        .Z(Red_ToCheckInst_LFInst_34_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_35_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_35_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_35_LFInst_0_n5), .ZN(Red_SignaltoCheck[35]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_35_LFInst_0_U2 ( .A(Output[14]), .B(
        Output[15]), .ZN(Red_ToCheckInst_LFInst_35_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_35_LFInst_0_U1 ( .A(Output[12]), .B(
        Output[13]), .Z(Red_ToCheckInst_LFInst_35_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_36_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_36_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_36_LFInst_0_n5), .ZN(Red_SignaltoCheck[36]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_36_LFInst_0_U2 ( .A(Output[18]), .B(
        Output[19]), .ZN(Red_ToCheckInst_LFInst_36_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_36_LFInst_0_U1 ( .A(Output[16]), .B(
        Output[17]), .Z(Red_ToCheckInst_LFInst_36_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_37_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_37_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_37_LFInst_0_n5), .ZN(Red_SignaltoCheck[37]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_37_LFInst_0_U2 ( .A(Output[22]), .B(
        Output[23]), .ZN(Red_ToCheckInst_LFInst_37_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_37_LFInst_0_U1 ( .A(Output[20]), .B(
        Output[21]), .Z(Red_ToCheckInst_LFInst_37_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_38_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_38_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_38_LFInst_0_n5), .ZN(Red_SignaltoCheck[38]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_38_LFInst_0_U2 ( .A(Output[26]), .B(
        Output[27]), .ZN(Red_ToCheckInst_LFInst_38_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_38_LFInst_0_U1 ( .A(Output[24]), .B(
        Output[25]), .Z(Red_ToCheckInst_LFInst_38_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_39_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_39_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_39_LFInst_0_n5), .ZN(Red_SignaltoCheck[39]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_39_LFInst_0_U2 ( .A(Output[30]), .B(
        Output[31]), .ZN(Red_ToCheckInst_LFInst_39_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_39_LFInst_0_U1 ( .A(Output[28]), .B(
        Output[29]), .Z(Red_ToCheckInst_LFInst_39_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_40_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_40_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_40_LFInst_0_n5), .ZN(Red_SignaltoCheck[40]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_40_LFInst_0_U2 ( .A(Output[34]), .B(
        Output[35]), .ZN(Red_ToCheckInst_LFInst_40_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_40_LFInst_0_U1 ( .A(Output[32]), .B(
        Output[33]), .Z(Red_ToCheckInst_LFInst_40_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_41_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_41_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_41_LFInst_0_n5), .ZN(Red_SignaltoCheck[41]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_41_LFInst_0_U2 ( .A(Output[38]), .B(
        Output[39]), .ZN(Red_ToCheckInst_LFInst_41_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_41_LFInst_0_U1 ( .A(Output[36]), .B(
        Output[37]), .Z(Red_ToCheckInst_LFInst_41_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_42_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_42_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_42_LFInst_0_n5), .ZN(Red_SignaltoCheck[42]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_42_LFInst_0_U2 ( .A(Output[42]), .B(
        Output[43]), .ZN(Red_ToCheckInst_LFInst_42_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_42_LFInst_0_U1 ( .A(Output[40]), .B(
        Output[41]), .Z(Red_ToCheckInst_LFInst_42_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_43_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_43_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_43_LFInst_0_n5), .ZN(Red_SignaltoCheck[43]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_43_LFInst_0_U2 ( .A(Output[46]), .B(
        Output[47]), .ZN(Red_ToCheckInst_LFInst_43_LFInst_0_n5) );
  XOR2_X1 Red_ToCheckInst_LFInst_43_LFInst_0_U1 ( .A(Output[44]), .B(
        Output[45]), .Z(Red_ToCheckInst_LFInst_43_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_44_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_44_LFInst_0_n5), .B(
        Red_ToCheckInst_LFInst_44_LFInst_0_n6), .ZN(Red_SignaltoCheck[44]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_44_LFInst_0_U2 ( .A(Output[48]), .B(
        Output[49]), .ZN(Red_ToCheckInst_LFInst_44_LFInst_0_n6) );
  XOR2_X1 Red_ToCheckInst_LFInst_44_LFInst_0_U1 ( .A(Output[51]), .B(
        Output[50]), .Z(Red_ToCheckInst_LFInst_44_LFInst_0_n5) );
  XNOR2_X1 Red_ToCheckInst_LFInst_45_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_45_LFInst_0_n5), .B(
        Red_ToCheckInst_LFInst_45_LFInst_0_n6), .ZN(Red_SignaltoCheck[45]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_45_LFInst_0_U2 ( .A(Output[52]), .B(
        Output[53]), .ZN(Red_ToCheckInst_LFInst_45_LFInst_0_n6) );
  XOR2_X1 Red_ToCheckInst_LFInst_45_LFInst_0_U1 ( .A(Output[55]), .B(
        Output[54]), .Z(Red_ToCheckInst_LFInst_45_LFInst_0_n5) );
  XNOR2_X1 Red_ToCheckInst_LFInst_46_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_46_LFInst_0_n5), .B(
        Red_ToCheckInst_LFInst_46_LFInst_0_n6), .ZN(Red_SignaltoCheck[46]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_46_LFInst_0_U2 ( .A(Output[56]), .B(
        Output[57]), .ZN(Red_ToCheckInst_LFInst_46_LFInst_0_n6) );
  XOR2_X1 Red_ToCheckInst_LFInst_46_LFInst_0_U1 ( .A(Output[59]), .B(
        Output[58]), .Z(Red_ToCheckInst_LFInst_46_LFInst_0_n5) );
  XNOR2_X1 Red_ToCheckInst_LFInst_47_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_47_LFInst_0_n5), .B(
        Red_ToCheckInst_LFInst_47_LFInst_0_n6), .ZN(Red_SignaltoCheck[47]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_47_LFInst_0_U2 ( .A(Output[60]), .B(
        Output[61]), .ZN(Red_ToCheckInst_LFInst_47_LFInst_0_n6) );
  XOR2_X1 Red_ToCheckInst_LFInst_47_LFInst_0_U1 ( .A(Output[63]), .B(
        Output[62]), .Z(Red_ToCheckInst_LFInst_47_LFInst_0_n5) );
  XNOR2_X1 Red_ToCheckInst_LFInst_48_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_48_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_48_LFInst_0_n5), .ZN(Red_SignaltoCheck[48]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_48_LFInst_0_U2 ( .A(PermutationOutput2[62]), 
        .B(PermutationOutput2[63]), .ZN(Red_ToCheckInst_LFInst_48_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_48_LFInst_0_U1 ( .A(PermutationOutput2[60]), 
        .B(PermutationOutput2[61]), .Z(Red_ToCheckInst_LFInst_48_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_49_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_49_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_49_LFInst_0_n5), .ZN(Red_SignaltoCheck[49]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_49_LFInst_0_U2 ( .A(PermutationOutput2[50]), 
        .B(PermutationOutput2[51]), .ZN(Red_ToCheckInst_LFInst_49_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_49_LFInst_0_U1 ( .A(PermutationOutput2[48]), 
        .B(PermutationOutput2[49]), .Z(Red_ToCheckInst_LFInst_49_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_50_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_50_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_50_LFInst_0_n5), .ZN(Red_SignaltoCheck[50]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_50_LFInst_0_U2 ( .A(PermutationOutput2[54]), 
        .B(PermutationOutput2[55]), .ZN(Red_ToCheckInst_LFInst_50_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_50_LFInst_0_U1 ( .A(PermutationOutput2[52]), 
        .B(PermutationOutput2[53]), .Z(Red_ToCheckInst_LFInst_50_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_51_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_51_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_51_LFInst_0_n5), .ZN(Red_SignaltoCheck[51]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_51_LFInst_0_U2 ( .A(PermutationOutput2[58]), 
        .B(PermutationOutput2[59]), .ZN(Red_ToCheckInst_LFInst_51_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_51_LFInst_0_U1 ( .A(PermutationOutput2[56]), 
        .B(PermutationOutput2[57]), .Z(Red_ToCheckInst_LFInst_51_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_52_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_52_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_52_LFInst_0_n5), .ZN(Red_SignaltoCheck[52]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_52_LFInst_0_U2 ( .A(PermutationOutput2[34]), 
        .B(PermutationOutput2[35]), .ZN(Red_ToCheckInst_LFInst_52_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_52_LFInst_0_U1 ( .A(PermutationOutput2[32]), 
        .B(PermutationOutput2[33]), .Z(Red_ToCheckInst_LFInst_52_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_53_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_53_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_53_LFInst_0_n5), .ZN(Red_SignaltoCheck[53]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_53_LFInst_0_U2 ( .A(PermutationOutput2[46]), 
        .B(PermutationOutput2[47]), .ZN(Red_ToCheckInst_LFInst_53_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_53_LFInst_0_U1 ( .A(PermutationOutput2[44]), 
        .B(PermutationOutput2[45]), .Z(Red_ToCheckInst_LFInst_53_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_54_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_54_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_54_LFInst_0_n5), .ZN(Red_SignaltoCheck[54]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_54_LFInst_0_U2 ( .A(PermutationOutput2[42]), 
        .B(PermutationOutput2[43]), .ZN(Red_ToCheckInst_LFInst_54_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_54_LFInst_0_U1 ( .A(PermutationOutput2[40]), 
        .B(PermutationOutput2[41]), .Z(Red_ToCheckInst_LFInst_54_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_55_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_55_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_55_LFInst_0_n5), .ZN(Red_SignaltoCheck[55]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_55_LFInst_0_U2 ( .A(PermutationOutput2[38]), 
        .B(PermutationOutput2[39]), .ZN(Red_ToCheckInst_LFInst_55_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_55_LFInst_0_U1 ( .A(PermutationOutput2[36]), 
        .B(PermutationOutput2[37]), .Z(Red_ToCheckInst_LFInst_55_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_56_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_56_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_56_LFInst_0_n5), .ZN(Red_SignaltoCheck[56]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_56_LFInst_0_U2 ( .A(PermutationOutput2[18]), 
        .B(PermutationOutput2[19]), .ZN(Red_ToCheckInst_LFInst_56_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_56_LFInst_0_U1 ( .A(PermutationOutput2[16]), 
        .B(PermutationOutput2[17]), .Z(Red_ToCheckInst_LFInst_56_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_57_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_57_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_57_LFInst_0_n5), .ZN(Red_SignaltoCheck[57]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_57_LFInst_0_U2 ( .A(PermutationOutput2[30]), 
        .B(PermutationOutput2[31]), .ZN(Red_ToCheckInst_LFInst_57_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_57_LFInst_0_U1 ( .A(PermutationOutput2[28]), 
        .B(PermutationOutput2[29]), .Z(Red_ToCheckInst_LFInst_57_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_58_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_58_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_58_LFInst_0_n5), .ZN(Red_SignaltoCheck[58]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_58_LFInst_0_U2 ( .A(PermutationOutput2[26]), 
        .B(PermutationOutput2[27]), .ZN(Red_ToCheckInst_LFInst_58_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_58_LFInst_0_U1 ( .A(PermutationOutput2[24]), 
        .B(PermutationOutput2[25]), .Z(Red_ToCheckInst_LFInst_58_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_59_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_59_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_59_LFInst_0_n5), .ZN(Red_SignaltoCheck[59]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_59_LFInst_0_U2 ( .A(PermutationOutput2[22]), 
        .B(PermutationOutput2[23]), .ZN(Red_ToCheckInst_LFInst_59_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_59_LFInst_0_U1 ( .A(PermutationOutput2[20]), 
        .B(PermutationOutput2[21]), .Z(Red_ToCheckInst_LFInst_59_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_60_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_60_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_60_LFInst_0_n5), .ZN(Red_SignaltoCheck[60]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_60_LFInst_0_U2 ( .A(PermutationOutput2[6]), 
        .B(PermutationOutput2[7]), .ZN(Red_ToCheckInst_LFInst_60_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_60_LFInst_0_U1 ( .A(PermutationOutput2[4]), 
        .B(PermutationOutput2[5]), .Z(Red_ToCheckInst_LFInst_60_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_61_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_61_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_61_LFInst_0_n5), .ZN(Red_SignaltoCheck[61]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_61_LFInst_0_U2 ( .A(PermutationOutput2[10]), 
        .B(PermutationOutput2[11]), .ZN(Red_ToCheckInst_LFInst_61_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_61_LFInst_0_U1 ( .A(PermutationOutput2[8]), 
        .B(PermutationOutput2[9]), .Z(Red_ToCheckInst_LFInst_61_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_62_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_62_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_62_LFInst_0_n5), .ZN(Red_SignaltoCheck[62]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_62_LFInst_0_U2 ( .A(PermutationOutput2[14]), 
        .B(PermutationOutput2[15]), .ZN(Red_ToCheckInst_LFInst_62_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_62_LFInst_0_U1 ( .A(PermutationOutput2[12]), 
        .B(PermutationOutput2[13]), .Z(Red_ToCheckInst_LFInst_62_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_63_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_63_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_63_LFInst_0_n5), .ZN(Red_SignaltoCheck[63]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_63_LFInst_0_U2 ( .A(PermutationOutput2[2]), 
        .B(PermutationOutput2[3]), .ZN(Red_ToCheckInst_LFInst_63_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_63_LFInst_0_U1 ( .A(PermutationOutput2[0]), 
        .B(PermutationOutput2[1]), .Z(Red_ToCheckInst_LFInst_63_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_64_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_64_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_64_LFInst_0_n5), .ZN(Red_SignaltoCheck[64]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_64_LFInst_0_U2 ( .A(PermutationOutput[62]), 
        .B(PermutationOutput[63]), .ZN(Red_ToCheckInst_LFInst_64_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_64_LFInst_0_U1 ( .A(PermutationOutput[60]), 
        .B(PermutationOutput[61]), .Z(Red_ToCheckInst_LFInst_64_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_65_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_65_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_65_LFInst_0_n5), .ZN(Red_SignaltoCheck[65]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_65_LFInst_0_U2 ( .A(PermutationOutput[50]), 
        .B(PermutationOutput[51]), .ZN(Red_ToCheckInst_LFInst_65_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_65_LFInst_0_U1 ( .A(PermutationOutput[48]), 
        .B(PermutationOutput[49]), .Z(Red_ToCheckInst_LFInst_65_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_66_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_66_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_66_LFInst_0_n5), .ZN(Red_SignaltoCheck[66]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_66_LFInst_0_U2 ( .A(PermutationOutput[54]), 
        .B(PermutationOutput[55]), .ZN(Red_ToCheckInst_LFInst_66_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_66_LFInst_0_U1 ( .A(PermutationOutput[52]), 
        .B(PermutationOutput[53]), .Z(Red_ToCheckInst_LFInst_66_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_67_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_67_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_67_LFInst_0_n5), .ZN(Red_SignaltoCheck[67]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_67_LFInst_0_U2 ( .A(PermutationOutput[58]), 
        .B(PermutationOutput[59]), .ZN(Red_ToCheckInst_LFInst_67_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_67_LFInst_0_U1 ( .A(PermutationOutput[56]), 
        .B(PermutationOutput[57]), .Z(Red_ToCheckInst_LFInst_67_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_68_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_68_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_68_LFInst_0_n5), .ZN(Red_SignaltoCheck[68]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_68_LFInst_0_U2 ( .A(PermutationOutput[34]), 
        .B(PermutationOutput[35]), .ZN(Red_ToCheckInst_LFInst_68_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_68_LFInst_0_U1 ( .A(PermutationOutput[32]), 
        .B(PermutationOutput[33]), .Z(Red_ToCheckInst_LFInst_68_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_69_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_69_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_69_LFInst_0_n5), .ZN(Red_SignaltoCheck[69]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_69_LFInst_0_U2 ( .A(PermutationOutput[46]), 
        .B(PermutationOutput[47]), .ZN(Red_ToCheckInst_LFInst_69_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_69_LFInst_0_U1 ( .A(PermutationOutput[44]), 
        .B(PermutationOutput[45]), .Z(Red_ToCheckInst_LFInst_69_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_70_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_70_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_70_LFInst_0_n5), .ZN(Red_SignaltoCheck[70]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_70_LFInst_0_U2 ( .A(PermutationOutput[42]), 
        .B(PermutationOutput[43]), .ZN(Red_ToCheckInst_LFInst_70_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_70_LFInst_0_U1 ( .A(PermutationOutput[40]), 
        .B(PermutationOutput[41]), .Z(Red_ToCheckInst_LFInst_70_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_71_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_71_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_71_LFInst_0_n5), .ZN(Red_SignaltoCheck[71]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_71_LFInst_0_U2 ( .A(PermutationOutput[38]), 
        .B(PermutationOutput[39]), .ZN(Red_ToCheckInst_LFInst_71_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_71_LFInst_0_U1 ( .A(PermutationOutput[36]), 
        .B(PermutationOutput[37]), .Z(Red_ToCheckInst_LFInst_71_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_72_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_72_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_72_LFInst_0_n5), .ZN(Red_SignaltoCheck[72]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_72_LFInst_0_U2 ( .A(PermutationOutput[18]), 
        .B(PermutationOutput[19]), .ZN(Red_ToCheckInst_LFInst_72_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_72_LFInst_0_U1 ( .A(PermutationOutput[16]), 
        .B(PermutationOutput[17]), .Z(Red_ToCheckInst_LFInst_72_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_73_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_73_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_73_LFInst_0_n5), .ZN(Red_SignaltoCheck[73]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_73_LFInst_0_U2 ( .A(PermutationOutput[30]), 
        .B(PermutationOutput[31]), .ZN(Red_ToCheckInst_LFInst_73_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_73_LFInst_0_U1 ( .A(PermutationOutput[28]), 
        .B(PermutationOutput[29]), .Z(Red_ToCheckInst_LFInst_73_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_74_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_74_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_74_LFInst_0_n5), .ZN(Red_SignaltoCheck[74]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_74_LFInst_0_U2 ( .A(PermutationOutput[26]), 
        .B(PermutationOutput[27]), .ZN(Red_ToCheckInst_LFInst_74_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_74_LFInst_0_U1 ( .A(PermutationOutput[24]), 
        .B(PermutationOutput[25]), .Z(Red_ToCheckInst_LFInst_74_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_75_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_75_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_75_LFInst_0_n5), .ZN(Red_SignaltoCheck[75]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_75_LFInst_0_U2 ( .A(PermutationOutput[22]), 
        .B(PermutationOutput[23]), .ZN(Red_ToCheckInst_LFInst_75_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_75_LFInst_0_U1 ( .A(PermutationOutput[20]), 
        .B(PermutationOutput[21]), .Z(Red_ToCheckInst_LFInst_75_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_76_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_76_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_76_LFInst_0_n5), .ZN(Red_SignaltoCheck[76]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_76_LFInst_0_U2 ( .A(PermutationOutput[6]), 
        .B(PermutationOutput[7]), .ZN(Red_ToCheckInst_LFInst_76_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_76_LFInst_0_U1 ( .A(PermutationOutput[4]), 
        .B(PermutationOutput[5]), .Z(Red_ToCheckInst_LFInst_76_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_77_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_77_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_77_LFInst_0_n5), .ZN(Red_SignaltoCheck[77]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_77_LFInst_0_U2 ( .A(PermutationOutput[10]), 
        .B(PermutationOutput[11]), .ZN(Red_ToCheckInst_LFInst_77_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_77_LFInst_0_U1 ( .A(PermutationOutput[8]), 
        .B(PermutationOutput[9]), .Z(Red_ToCheckInst_LFInst_77_LFInst_0_n6) );
  XNOR2_X1 Red_ToCheckInst_LFInst_78_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_78_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_78_LFInst_0_n5), .ZN(Red_SignaltoCheck[78]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_78_LFInst_0_U2 ( .A(PermutationOutput[14]), 
        .B(PermutationOutput[15]), .ZN(Red_ToCheckInst_LFInst_78_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_78_LFInst_0_U1 ( .A(PermutationOutput[12]), 
        .B(PermutationOutput[13]), .Z(Red_ToCheckInst_LFInst_78_LFInst_0_n6)
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_79_LFInst_0_U3 ( .A(
        Red_ToCheckInst_LFInst_79_LFInst_0_n6), .B(
        Red_ToCheckInst_LFInst_79_LFInst_0_n5), .ZN(Red_SignaltoCheck[79]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_79_LFInst_0_U2 ( .A(PermutationOutput[2]), 
        .B(PermutationOutput[3]), .ZN(Red_ToCheckInst_LFInst_79_LFInst_0_n5)
         );
  XOR2_X1 Red_ToCheckInst_LFInst_79_LFInst_0_U1 ( .A(PermutationOutput[0]), 
        .B(PermutationOutput[1]), .Z(Red_ToCheckInst_LFInst_79_LFInst_0_n6) );
  NOR2_X1 Check1_CheckInst_0_U159 ( .A1(Check1_CheckInst_0_n158), .A2(
        Check1_CheckInst_0_n157), .ZN(Error_0_) );
  NAND2_X1 Check1_CheckInst_0_U158 ( .A1(Check1_CheckInst_0_n156), .A2(
        Check1_CheckInst_0_n155), .ZN(Check1_CheckInst_0_n157) );
  NOR2_X1 Check1_CheckInst_0_U157 ( .A1(Check1_CheckInst_0_n154), .A2(
        Check1_CheckInst_0_n153), .ZN(Check1_CheckInst_0_n155) );
  NAND2_X1 Check1_CheckInst_0_U156 ( .A1(Check1_CheckInst_0_n152), .A2(
        Check1_CheckInst_0_n151), .ZN(Check1_CheckInst_0_n153) );
  NOR2_X1 Check1_CheckInst_0_U155 ( .A1(Check1_CheckInst_0_n150), .A2(
        Check1_CheckInst_0_n149), .ZN(Check1_CheckInst_0_n151) );
  NAND2_X1 Check1_CheckInst_0_U154 ( .A1(Check1_CheckInst_0_n148), .A2(
        Check1_CheckInst_0_n147), .ZN(Check1_CheckInst_0_n149) );
  NOR2_X1 Check1_CheckInst_0_U153 ( .A1(Check1_CheckInst_0_n146), .A2(
        Check1_CheckInst_0_n145), .ZN(Check1_CheckInst_0_n147) );
  XOR2_X1 Check1_CheckInst_0_U152 ( .A(Red_Feedback[9]), .B(
        Red_SignaltoCheck[41]), .Z(Check1_CheckInst_0_n145) );
  XOR2_X1 Check1_CheckInst_0_U151 ( .A(Red_Feedback[8]), .B(
        Red_SignaltoCheck[40]), .Z(Check1_CheckInst_0_n146) );
  XNOR2_X1 Check1_CheckInst_0_U150 ( .A(Red_Feedback[7]), .B(
        Red_SignaltoCheck[39]), .ZN(Check1_CheckInst_0_n148) );
  NAND2_X1 Check1_CheckInst_0_U149 ( .A1(Check1_CheckInst_0_n144), .A2(
        Check1_CheckInst_0_n143), .ZN(Check1_CheckInst_0_n150) );
  NOR2_X1 Check1_CheckInst_0_U148 ( .A1(Check1_CheckInst_0_n142), .A2(
        Check1_CheckInst_0_n141), .ZN(Check1_CheckInst_0_n143) );
  NAND2_X1 Check1_CheckInst_0_U147 ( .A1(Check1_CheckInst_0_n140), .A2(
        Check1_CheckInst_0_n139), .ZN(Check1_CheckInst_0_n141) );
  NOR2_X1 Check1_CheckInst_0_U146 ( .A1(Check1_CheckInst_0_n138), .A2(
        Check1_CheckInst_0_n137), .ZN(Check1_CheckInst_0_n139) );
  XOR2_X1 Check1_CheckInst_0_U145 ( .A(Red_StateRegOutput2[6]), .B(
        Red_SignaltoCheck[54]), .Z(Check1_CheckInst_0_n137) );
  XOR2_X1 Check1_CheckInst_0_U144 ( .A(Red_StateRegOutput2[8]), .B(
        Red_SignaltoCheck[56]), .Z(Check1_CheckInst_0_n138) );
  XNOR2_X1 Check1_CheckInst_0_U143 ( .A(Red_Feedback[11]), .B(
        Red_SignaltoCheck[43]), .ZN(Check1_CheckInst_0_n140) );
  NAND2_X1 Check1_CheckInst_0_U142 ( .A1(Check1_CheckInst_0_n136), .A2(
        Check1_CheckInst_0_n135), .ZN(Check1_CheckInst_0_n142) );
  NOR2_X1 Check1_CheckInst_0_U141 ( .A1(Check1_CheckInst_0_n134), .A2(
        Check1_CheckInst_0_n133), .ZN(Check1_CheckInst_0_n135) );
  NAND2_X1 Check1_CheckInst_0_U140 ( .A1(Check1_CheckInst_0_n132), .A2(
        Check1_CheckInst_0_n131), .ZN(Check1_CheckInst_0_n133) );
  NOR2_X1 Check1_CheckInst_0_U139 ( .A1(Check1_CheckInst_0_n130), .A2(
        Check1_CheckInst_0_n129), .ZN(Check1_CheckInst_0_n131) );
  XOR2_X1 Check1_CheckInst_0_U138 ( .A(Red_StateRegOutput2[10]), .B(
        Red_SignaltoCheck[58]), .Z(Check1_CheckInst_0_n129) );
  XOR2_X1 Check1_CheckInst_0_U137 ( .A(Red_StateRegOutput2[1]), .B(
        Red_SignaltoCheck[49]), .Z(Check1_CheckInst_0_n130) );
  XNOR2_X1 Check1_CheckInst_0_U136 ( .A(Red_StateRegOutput2[9]), .B(
        Red_SignaltoCheck[57]), .ZN(Check1_CheckInst_0_n132) );
  NAND2_X1 Check1_CheckInst_0_U135 ( .A1(Check1_CheckInst_0_n128), .A2(
        Check1_CheckInst_0_n127), .ZN(Check1_CheckInst_0_n134) );
  NOR2_X1 Check1_CheckInst_0_U134 ( .A1(Check1_CheckInst_0_n126), .A2(
        Check1_CheckInst_0_n125), .ZN(Check1_CheckInst_0_n127) );
  XOR2_X1 Check1_CheckInst_0_U133 ( .A(Red_StateRegOutput2[3]), .B(
        Red_SignaltoCheck[51]), .Z(Check1_CheckInst_0_n125) );
  XOR2_X1 Check1_CheckInst_0_U132 ( .A(Red_StateRegOutput2[2]), .B(
        Red_SignaltoCheck[50]), .Z(Check1_CheckInst_0_n126) );
  NOR2_X1 Check1_CheckInst_0_U131 ( .A1(Check1_CheckInst_0_n124), .A2(
        Check1_CheckInst_0_n123), .ZN(Check1_CheckInst_0_n128) );
  XOR2_X1 Check1_CheckInst_0_U130 ( .A(Red_StateRegOutput2[4]), .B(
        Red_SignaltoCheck[52]), .Z(Check1_CheckInst_0_n123) );
  XOR2_X1 Check1_CheckInst_0_U129 ( .A(Red_StateRegOutput2[5]), .B(
        Red_SignaltoCheck[53]), .Z(Check1_CheckInst_0_n124) );
  XNOR2_X1 Check1_CheckInst_0_U128 ( .A(Red_SignaltoCheck[55]), .B(
        Red_StateRegOutput2[7]), .ZN(Check1_CheckInst_0_n136) );
  XNOR2_X1 Check1_CheckInst_0_U127 ( .A(Red_SignaltoCheck[42]), .B(
        Red_Feedback[10]), .ZN(Check1_CheckInst_0_n144) );
  XNOR2_X1 Check1_CheckInst_0_U126 ( .A(Red_SignaltoCheck[48]), .B(
        Red_StateRegOutput2[0]), .ZN(Check1_CheckInst_0_n152) );
  NAND2_X1 Check1_CheckInst_0_U125 ( .A1(Check1_CheckInst_0_n122), .A2(
        Check1_CheckInst_0_n121), .ZN(Check1_CheckInst_0_n154) );
  NOR2_X1 Check1_CheckInst_0_U124 ( .A1(Check1_CheckInst_0_n120), .A2(
        Check1_CheckInst_0_n119), .ZN(Check1_CheckInst_0_n121) );
  NAND2_X1 Check1_CheckInst_0_U123 ( .A1(Check1_CheckInst_0_n118), .A2(
        Check1_CheckInst_0_n117), .ZN(Check1_CheckInst_0_n119) );
  NOR2_X1 Check1_CheckInst_0_U122 ( .A1(Check1_CheckInst_0_n116), .A2(
        Check1_CheckInst_0_n115), .ZN(Check1_CheckInst_0_n117) );
  XOR2_X1 Check1_CheckInst_0_U121 ( .A(Red_StateRegOutput[10]), .B(
        Red_SignaltoCheck[74]), .Z(Check1_CheckInst_0_n115) );
  XOR2_X1 Check1_CheckInst_0_U120 ( .A(Red_StateRegOutput[12]), .B(
        Red_SignaltoCheck[76]), .Z(Check1_CheckInst_0_n116) );
  XNOR2_X1 Check1_CheckInst_0_U119 ( .A(Red_StateRegOutput2[15]), .B(
        Red_SignaltoCheck[63]), .ZN(Check1_CheckInst_0_n118) );
  NAND2_X1 Check1_CheckInst_0_U118 ( .A1(Check1_CheckInst_0_n114), .A2(
        Check1_CheckInst_0_n113), .ZN(Check1_CheckInst_0_n120) );
  NOR2_X1 Check1_CheckInst_0_U117 ( .A1(Check1_CheckInst_0_n112), .A2(
        Check1_CheckInst_0_n111), .ZN(Check1_CheckInst_0_n113) );
  NAND2_X1 Check1_CheckInst_0_U116 ( .A1(Check1_CheckInst_0_n110), .A2(
        Check1_CheckInst_0_n109), .ZN(Check1_CheckInst_0_n111) );
  NOR2_X1 Check1_CheckInst_0_U115 ( .A1(Check1_CheckInst_0_n108), .A2(
        Check1_CheckInst_0_n107), .ZN(Check1_CheckInst_0_n109) );
  XOR2_X1 Check1_CheckInst_0_U114 ( .A(Red_StateRegOutput[14]), .B(
        Red_SignaltoCheck[78]), .Z(Check1_CheckInst_0_n107) );
  XOR2_X1 Check1_CheckInst_0_U113 ( .A(Red_StateRegOutput[5]), .B(
        Red_SignaltoCheck[69]), .Z(Check1_CheckInst_0_n108) );
  XNOR2_X1 Check1_CheckInst_0_U112 ( .A(Red_StateRegOutput[13]), .B(
        Red_SignaltoCheck[77]), .ZN(Check1_CheckInst_0_n110) );
  NAND2_X1 Check1_CheckInst_0_U111 ( .A1(Check1_CheckInst_0_n106), .A2(
        Check1_CheckInst_0_n105), .ZN(Check1_CheckInst_0_n112) );
  NOR2_X1 Check1_CheckInst_0_U110 ( .A1(Check1_CheckInst_0_n104), .A2(
        Check1_CheckInst_0_n103), .ZN(Check1_CheckInst_0_n105) );
  NAND2_X1 Check1_CheckInst_0_U109 ( .A1(Check1_CheckInst_0_n102), .A2(
        Check1_CheckInst_0_n101), .ZN(Check1_CheckInst_0_n103) );
  NOR2_X1 Check1_CheckInst_0_U108 ( .A1(Check1_CheckInst_0_n100), .A2(
        Check1_CheckInst_0_n99), .ZN(Check1_CheckInst_0_n101) );
  XOR2_X1 Check1_CheckInst_0_U107 ( .A(Red_StateRegOutput[8]), .B(
        Red_SignaltoCheck[72]), .Z(Check1_CheckInst_0_n99) );
  XOR2_X1 Check1_CheckInst_0_U106 ( .A(Red_StateRegOutput[9]), .B(
        Red_SignaltoCheck[73]), .Z(Check1_CheckInst_0_n100) );
  XNOR2_X1 Check1_CheckInst_0_U105 ( .A(Red_StateRegOutput[6]), .B(
        Red_SignaltoCheck[70]), .ZN(Check1_CheckInst_0_n102) );
  NAND2_X1 Check1_CheckInst_0_U104 ( .A1(Check1_CheckInst_0_n98), .A2(
        Check1_CheckInst_0_n97), .ZN(Check1_CheckInst_0_n104) );
  NOR2_X1 Check1_CheckInst_0_U103 ( .A1(Check1_CheckInst_0_n96), .A2(
        Check1_CheckInst_0_n95), .ZN(Check1_CheckInst_0_n97) );
  NOR2_X1 Check1_CheckInst_0_U102 ( .A1(Check1_CheckInst_0_n94), .A2(
        Check1_CheckInst_0_n93), .ZN(Check1_CheckInst_0_n98) );
  XNOR2_X1 Check1_CheckInst_0_U101 ( .A(Red_SignaltoCheck[71]), .B(
        Red_StateRegOutput[7]), .ZN(Check1_CheckInst_0_n106) );
  XNOR2_X1 Check1_CheckInst_0_U100 ( .A(Red_SignaltoCheck[75]), .B(
        Red_StateRegOutput[11]), .ZN(Check1_CheckInst_0_n114) );
  XNOR2_X1 Check1_CheckInst_0_U99 ( .A(Red_SignaltoCheck[62]), .B(
        Red_StateRegOutput2[14]), .ZN(Check1_CheckInst_0_n122) );
  NOR2_X1 Check1_CheckInst_0_U98 ( .A1(Check1_CheckInst_0_n92), .A2(
        Check1_CheckInst_0_n91), .ZN(Check1_CheckInst_0_n156) );
  NAND2_X1 Check1_CheckInst_0_U97 ( .A1(Check1_CheckInst_0_n90), .A2(
        Check1_CheckInst_0_n89), .ZN(Check1_CheckInst_0_n91) );
  NOR2_X1 Check1_CheckInst_0_U96 ( .A1(Check1_CheckInst_0_n88), .A2(
        Check1_CheckInst_0_n87), .ZN(Check1_CheckInst_0_n89) );
  NAND2_X1 Check1_CheckInst_0_U95 ( .A1(Check1_CheckInst_0_n86), .A2(
        Check1_CheckInst_0_n85), .ZN(Check1_CheckInst_0_n87) );
  NOR2_X1 Check1_CheckInst_0_U94 ( .A1(Check1_CheckInst_0_n84), .A2(
        Check1_CheckInst_0_n83), .ZN(Check1_CheckInst_0_n85) );
  NAND2_X1 Check1_CheckInst_0_U93 ( .A1(Check1_CheckInst_0_n82), .A2(
        Check1_CheckInst_0_n81), .ZN(Check1_CheckInst_0_n83) );
  NOR2_X1 Check1_CheckInst_0_U92 ( .A1(Check1_CheckInst_0_n80), .A2(
        Check1_CheckInst_0_n79), .ZN(Check1_CheckInst_0_n81) );
  XOR2_X1 Check1_CheckInst_0_U91 ( .A(Red_final[21]), .B(Red_SignaltoCheck[21]), .Z(Check1_CheckInst_0_n79) );
  XOR2_X1 Check1_CheckInst_0_U90 ( .A(Red_final[22]), .B(Red_SignaltoCheck[22]), .Z(Check1_CheckInst_0_n80) );
  NOR2_X1 Check1_CheckInst_0_U89 ( .A1(Check1_CheckInst_0_n78), .A2(
        Check1_CheckInst_0_n77), .ZN(Check1_CheckInst_0_n82) );
  XOR2_X1 Check1_CheckInst_0_U88 ( .A(Red_Feedback[3]), .B(
        Red_SignaltoCheck[35]), .Z(Check1_CheckInst_0_n77) );
  XOR2_X1 Check1_CheckInst_0_U87 ( .A(Red_Feedback[2]), .B(
        Red_SignaltoCheck[34]), .Z(Check1_CheckInst_0_n78) );
  NAND2_X1 Check1_CheckInst_0_U86 ( .A1(Check1_CheckInst_0_n76), .A2(
        Check1_CheckInst_0_n75), .ZN(Check1_CheckInst_0_n84) );
  XNOR2_X1 Check1_CheckInst_0_U85 ( .A(Red_Feedback[5]), .B(
        Red_SignaltoCheck[37]), .ZN(Check1_CheckInst_0_n75) );
  XNOR2_X1 Check1_CheckInst_0_U84 ( .A(Red_Feedback[6]), .B(
        Red_SignaltoCheck[38]), .ZN(Check1_CheckInst_0_n76) );
  NOR2_X1 Check1_CheckInst_0_U83 ( .A1(Check1_CheckInst_0_n74), .A2(
        Check1_CheckInst_0_n73), .ZN(Check1_CheckInst_0_n86) );
  XOR2_X1 Check1_CheckInst_0_U82 ( .A(Red_final[29]), .B(Red_SignaltoCheck[29]), .Z(Check1_CheckInst_0_n73) );
  XOR2_X1 Check1_CheckInst_0_U81 ( .A(Red_Feedback[4]), .B(
        Red_SignaltoCheck[36]), .Z(Check1_CheckInst_0_n74) );
  NAND2_X1 Check1_CheckInst_0_U80 ( .A1(Check1_CheckInst_0_n72), .A2(
        Check1_CheckInst_0_n71), .ZN(Check1_CheckInst_0_n88) );
  NOR2_X1 Check1_CheckInst_0_U79 ( .A1(Check1_CheckInst_0_n70), .A2(
        Check1_CheckInst_0_n69), .ZN(Check1_CheckInst_0_n71) );
  NAND2_X1 Check1_CheckInst_0_U78 ( .A1(Check1_CheckInst_0_n68), .A2(
        Check1_CheckInst_0_n67), .ZN(Check1_CheckInst_0_n69) );
  NOR2_X1 Check1_CheckInst_0_U77 ( .A1(Check1_CheckInst_0_n66), .A2(
        Check1_CheckInst_0_n65), .ZN(Check1_CheckInst_0_n67) );
  XOR2_X1 Check1_CheckInst_0_U76 ( .A(Red_Feedback[1]), .B(
        Red_SignaltoCheck[33]), .Z(Check1_CheckInst_0_n65) );
  XOR2_X1 Check1_CheckInst_0_U75 ( .A(Red_final[30]), .B(Red_SignaltoCheck[30]), .Z(Check1_CheckInst_0_n66) );
  NOR2_X1 Check1_CheckInst_0_U74 ( .A1(Check1_CheckInst_0_n64), .A2(
        Check1_CheckInst_0_n63), .ZN(Check1_CheckInst_0_n68) );
  XOR2_X1 Check1_CheckInst_0_U73 ( .A(Red_final[31]), .B(Red_SignaltoCheck[31]), .Z(Check1_CheckInst_0_n63) );
  XOR2_X1 Check1_CheckInst_0_U72 ( .A(Red_Feedback[0]), .B(
        Red_SignaltoCheck[32]), .Z(Check1_CheckInst_0_n64) );
  NAND2_X1 Check1_CheckInst_0_U71 ( .A1(Check1_CheckInst_0_n62), .A2(
        Check1_CheckInst_0_n61), .ZN(Check1_CheckInst_0_n70) );
  XNOR2_X1 Check1_CheckInst_0_U70 ( .A(Red_final[5]), .B(Red_SignaltoCheck[5]), 
        .ZN(Check1_CheckInst_0_n61) );
  XNOR2_X1 Check1_CheckInst_0_U69 ( .A(Red_final[4]), .B(Red_SignaltoCheck[4]), 
        .ZN(Check1_CheckInst_0_n62) );
  NOR2_X1 Check1_CheckInst_0_U68 ( .A1(Check1_CheckInst_0_n60), .A2(
        Check1_CheckInst_0_n59), .ZN(Check1_CheckInst_0_n72) );
  XOR2_X1 Check1_CheckInst_0_U67 ( .A(Red_final[7]), .B(Red_SignaltoCheck[7]), 
        .Z(Check1_CheckInst_0_n59) );
  XOR2_X1 Check1_CheckInst_0_U66 ( .A(Red_final[8]), .B(Red_SignaltoCheck[8]), 
        .Z(Check1_CheckInst_0_n60) );
  NOR2_X1 Check1_CheckInst_0_U65 ( .A1(Check1_CheckInst_0_n58), .A2(
        Check1_CheckInst_0_n57), .ZN(Check1_CheckInst_0_n90) );
  NAND2_X1 Check1_CheckInst_0_U64 ( .A1(Check1_CheckInst_0_n56), .A2(
        Check1_CheckInst_0_n55), .ZN(Check1_CheckInst_0_n57) );
  NOR2_X1 Check1_CheckInst_0_U63 ( .A1(Check1_CheckInst_0_n54), .A2(
        Check1_CheckInst_0_n53), .ZN(Check1_CheckInst_0_n55) );
  NAND2_X1 Check1_CheckInst_0_U62 ( .A1(Check1_CheckInst_0_n52), .A2(
        Check1_CheckInst_0_n51), .ZN(Check1_CheckInst_0_n53) );
  XNOR2_X1 Check1_CheckInst_0_U61 ( .A(Red_SignaltoCheck[0]), .B(Red_final[0]), 
        .ZN(Check1_CheckInst_0_n51) );
  XNOR2_X1 Check1_CheckInst_0_U60 ( .A(Red_final[6]), .B(Red_SignaltoCheck[6]), 
        .ZN(Check1_CheckInst_0_n52) );
  NAND2_X1 Check1_CheckInst_0_U59 ( .A1(Check1_CheckInst_0_n50), .A2(
        Check1_CheckInst_0_n49), .ZN(Check1_CheckInst_0_n54) );
  XNOR2_X1 Check1_CheckInst_0_U58 ( .A(Red_final[3]), .B(Red_SignaltoCheck[3]), 
        .ZN(Check1_CheckInst_0_n49) );
  XNOR2_X1 Check1_CheckInst_0_U57 ( .A(Red_SignaltoCheck[1]), .B(Red_final[1]), 
        .ZN(Check1_CheckInst_0_n50) );
  NOR2_X1 Check1_CheckInst_0_U56 ( .A1(Check1_CheckInst_0_n48), .A2(
        Check1_CheckInst_0_n47), .ZN(Check1_CheckInst_0_n56) );
  XOR2_X1 Check1_CheckInst_0_U55 ( .A(Red_StateRegOutput[15]), .B(
        Red_SignaltoCheck[79]), .Z(Check1_CheckInst_0_n47) );
  XOR2_X1 Check1_CheckInst_0_U54 ( .A(Red_final[2]), .B(Red_SignaltoCheck[2]), 
        .Z(Check1_CheckInst_0_n48) );
  NAND2_X1 Check1_CheckInst_0_U53 ( .A1(Check1_CheckInst_0_n46), .A2(
        Check1_CheckInst_0_n45), .ZN(Check1_CheckInst_0_n58) );
  XNOR2_X1 Check1_CheckInst_0_U52 ( .A(Red_final[15]), .B(
        Red_SignaltoCheck[15]), .ZN(Check1_CheckInst_0_n45) );
  XNOR2_X1 Check1_CheckInst_0_U51 ( .A(Red_final[14]), .B(
        Red_SignaltoCheck[14]), .ZN(Check1_CheckInst_0_n46) );
  NAND2_X1 Check1_CheckInst_0_U50 ( .A1(Check1_CheckInst_0_n44), .A2(
        Check1_CheckInst_0_n43), .ZN(Check1_CheckInst_0_n92) );
  NOR2_X1 Check1_CheckInst_0_U49 ( .A1(Check1_CheckInst_0_n42), .A2(
        Check1_CheckInst_0_n41), .ZN(Check1_CheckInst_0_n43) );
  NAND2_X1 Check1_CheckInst_0_U48 ( .A1(Check1_CheckInst_0_n40), .A2(
        Check1_CheckInst_0_n39), .ZN(Check1_CheckInst_0_n41) );
  NOR2_X1 Check1_CheckInst_0_U47 ( .A1(Check1_CheckInst_0_n38), .A2(
        Check1_CheckInst_0_n37), .ZN(Check1_CheckInst_0_n39) );
  XOR2_X1 Check1_CheckInst_0_U46 ( .A(Red_final[17]), .B(Red_SignaltoCheck[17]), .Z(Check1_CheckInst_0_n37) );
  XOR2_X1 Check1_CheckInst_0_U45 ( .A(Red_final[18]), .B(Red_SignaltoCheck[18]), .Z(Check1_CheckInst_0_n38) );
  NOR2_X1 Check1_CheckInst_0_U44 ( .A1(Check1_CheckInst_0_n36), .A2(
        Check1_CheckInst_0_n35), .ZN(Check1_CheckInst_0_n40) );
  XOR2_X1 Check1_CheckInst_0_U43 ( .A(Red_final[9]), .B(Red_SignaltoCheck[9]), 
        .Z(Check1_CheckInst_0_n35) );
  XOR2_X1 Check1_CheckInst_0_U42 ( .A(Red_final[16]), .B(Red_SignaltoCheck[16]), .Z(Check1_CheckInst_0_n36) );
  NAND2_X1 Check1_CheckInst_0_U41 ( .A1(Check1_CheckInst_0_n34), .A2(
        Check1_CheckInst_0_n33), .ZN(Check1_CheckInst_0_n42) );
  XNOR2_X1 Check1_CheckInst_0_U40 ( .A(Red_final[13]), .B(
        Red_SignaltoCheck[13]), .ZN(Check1_CheckInst_0_n33) );
  XNOR2_X1 Check1_CheckInst_0_U39 ( .A(Red_final[10]), .B(
        Red_SignaltoCheck[10]), .ZN(Check1_CheckInst_0_n34) );
  NOR2_X1 Check1_CheckInst_0_U38 ( .A1(Check1_CheckInst_0_n32), .A2(
        Check1_CheckInst_0_n31), .ZN(Check1_CheckInst_0_n44) );
  XOR2_X1 Check1_CheckInst_0_U37 ( .A(Red_final[11]), .B(Red_SignaltoCheck[11]), .Z(Check1_CheckInst_0_n31) );
  XOR2_X1 Check1_CheckInst_0_U36 ( .A(Red_final[12]), .B(Red_SignaltoCheck[12]), .Z(Check1_CheckInst_0_n32) );
  NAND2_X1 Check1_CheckInst_0_U35 ( .A1(Check1_CheckInst_0_n30), .A2(
        Check1_CheckInst_0_n29), .ZN(Check1_CheckInst_0_n158) );
  NOR2_X1 Check1_CheckInst_0_U34 ( .A1(Check1_CheckInst_0_n28), .A2(
        Check1_CheckInst_0_n27), .ZN(Check1_CheckInst_0_n29) );
  NAND2_X1 Check1_CheckInst_0_U33 ( .A1(Check1_CheckInst_0_n26), .A2(
        Check1_CheckInst_0_n25), .ZN(Check1_CheckInst_0_n27) );
  NOR2_X1 Check1_CheckInst_0_U32 ( .A1(Check1_CheckInst_0_n24), .A2(
        Check1_CheckInst_0_n23), .ZN(Check1_CheckInst_0_n25) );
  XOR2_X1 Check1_CheckInst_0_U31 ( .A(Red_final[19]), .B(Red_SignaltoCheck[19]), .Z(Check1_CheckInst_0_n23) );
  XOR2_X1 Check1_CheckInst_0_U30 ( .A(Red_final[26]), .B(Red_SignaltoCheck[26]), .Z(Check1_CheckInst_0_n24) );
  XNOR2_X1 Check1_CheckInst_0_U29 ( .A(Red_final[20]), .B(
        Red_SignaltoCheck[20]), .ZN(Check1_CheckInst_0_n26) );
  NAND2_X1 Check1_CheckInst_0_U28 ( .A1(Check1_CheckInst_0_n22), .A2(
        Check1_CheckInst_0_n21), .ZN(Check1_CheckInst_0_n28) );
  NOR2_X1 Check1_CheckInst_0_U27 ( .A1(Check1_CheckInst_0_n20), .A2(
        Check1_CheckInst_0_n19), .ZN(Check1_CheckInst_0_n21) );
  NAND2_X1 Check1_CheckInst_0_U26 ( .A1(Check1_CheckInst_0_n18), .A2(
        Check1_CheckInst_0_n17), .ZN(Check1_CheckInst_0_n19) );
  NOR2_X1 Check1_CheckInst_0_U25 ( .A1(Check1_CheckInst_0_n16), .A2(
        Check1_CheckInst_0_n15), .ZN(Check1_CheckInst_0_n17) );
  XOR2_X1 Check1_CheckInst_0_U24 ( .A(Red_final[25]), .B(Red_SignaltoCheck[25]), .Z(Check1_CheckInst_0_n15) );
  XOR2_X1 Check1_CheckInst_0_U23 ( .A(Red_final[24]), .B(Red_SignaltoCheck[24]), .Z(Check1_CheckInst_0_n16) );
  XNOR2_X1 Check1_CheckInst_0_U22 ( .A(Red_final[28]), .B(
        Red_SignaltoCheck[28]), .ZN(Check1_CheckInst_0_n18) );
  NAND2_X1 Check1_CheckInst_0_U21 ( .A1(Check1_CheckInst_0_n14), .A2(
        Check1_CheckInst_0_n13), .ZN(Check1_CheckInst_0_n20) );
  NOR2_X1 Check1_CheckInst_0_U20 ( .A1(Check1_CheckInst_0_n12), .A2(
        Check1_CheckInst_0_n11), .ZN(Check1_CheckInst_0_n13) );
  NAND2_X1 Check1_CheckInst_0_U19 ( .A1(Check1_CheckInst_0_n10), .A2(
        Check1_CheckInst_0_n9), .ZN(Check1_CheckInst_0_n11) );
  NOR2_X1 Check1_CheckInst_0_U18 ( .A1(Check1_CheckInst_0_n8), .A2(
        Check1_CheckInst_0_n7), .ZN(Check1_CheckInst_0_n9) );
  XOR2_X1 Check1_CheckInst_0_U17 ( .A(Red_StateRegOutput[1]), .B(
        Red_SignaltoCheck[65]), .Z(Check1_CheckInst_0_n7) );
  XOR2_X1 Check1_CheckInst_0_U16 ( .A(Red_StateRegOutput[3]), .B(
        Red_SignaltoCheck[67]), .Z(Check1_CheckInst_0_n8) );
  XNOR2_X1 Check1_CheckInst_0_U15 ( .A(Red_StateRegOutput[2]), .B(
        Red_SignaltoCheck[66]), .ZN(Check1_CheckInst_0_n10) );
  NAND2_X1 Check1_CheckInst_0_U14 ( .A1(Check1_CheckInst_0_n6), .A2(
        Check1_CheckInst_0_n5), .ZN(Check1_CheckInst_0_n12) );
  NOR2_X1 Check1_CheckInst_0_U13 ( .A1(Check1_CheckInst_0_n4), .A2(
        Check1_CheckInst_0_n3), .ZN(Check1_CheckInst_0_n5) );
  XOR2_X1 Check1_CheckInst_0_U12 ( .A(Red_StateRegOutput[4]), .B(
        Red_SignaltoCheck[68]), .Z(Check1_CheckInst_0_n3) );
  XOR2_X1 Check1_CheckInst_0_U11 ( .A(Red_StateRegOutput2[11]), .B(
        Red_SignaltoCheck[59]), .Z(Check1_CheckInst_0_n4) );
  NOR2_X1 Check1_CheckInst_0_U10 ( .A1(Check1_CheckInst_0_n2), .A2(
        Check1_CheckInst_0_n1), .ZN(Check1_CheckInst_0_n6) );
  XOR2_X1 Check1_CheckInst_0_U9 ( .A(Red_StateRegOutput2[13]), .B(
        Red_SignaltoCheck[61]), .Z(Check1_CheckInst_0_n1) );
  XOR2_X1 Check1_CheckInst_0_U8 ( .A(Red_StateRegOutput2[12]), .B(
        Red_SignaltoCheck[60]), .Z(Check1_CheckInst_0_n2) );
  XNOR2_X1 Check1_CheckInst_0_U7 ( .A(Red_SignaltoCheck[64]), .B(
        Red_StateRegOutput[0]), .ZN(Check1_CheckInst_0_n14) );
  XNOR2_X1 Check1_CheckInst_0_U6 ( .A(Red_SignaltoCheck[27]), .B(Red_final[27]), .ZN(Check1_CheckInst_0_n22) );
  XNOR2_X1 Check1_CheckInst_0_U5 ( .A(Red_SignaltoCheck[23]), .B(Red_final[23]), .ZN(Check1_CheckInst_0_n30) );
  XOR2_X1 Check1_CheckInst_0_U4 ( .A(Red_Feedback[15]), .B(
        Red_SignaltoCheck[47]), .Z(Check1_CheckInst_0_n94) );
  XOR2_X1 Check1_CheckInst_0_U3 ( .A(Red_Feedback[13]), .B(
        Red_SignaltoCheck[45]), .Z(Check1_CheckInst_0_n93) );
  XOR2_X1 Check1_CheckInst_0_U2 ( .A(Red_Feedback[14]), .B(
        Red_SignaltoCheck[46]), .Z(Check1_CheckInst_0_n96) );
  XOR2_X1 Check1_CheckInst_0_U1 ( .A(Red_Feedback[12]), .B(
        Red_SignaltoCheck[44]), .Z(Check1_CheckInst_0_n95) );
endmodule

