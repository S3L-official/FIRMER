module LED64Enc ( clk, rst, Plaintext, Key, Ciphertext, ErrorFlag );
  input [63:0] Plaintext;
  input [63:0] Key;
  output [63:0] Ciphertext;
  (* FIRMER="clock" *)input clk;
  output ErrorFlag;
  wire   Error [0] , AddKeyXOR_XORInst_0_0_n2 , AddKeyXOR_XORInst_0_2_n2 ,
         AddKeyXOR_XORInst_1_0_n2 , AddKeyXOR_XORInst_1_2_n2 ,
         AddKeyXOR_XORInst_2_0_n2 , AddKeyXOR_XORInst_2_2_n2 ,
         AddKeyXOR_XORInst_3_0_n2 , AddKeyXOR_XORInst_3_2_n2 ,
         AddKeyXOR_XORInst_4_0_n2 , AddKeyXOR_XORInst_4_2_n2 ,
         AddKeyXOR_XORInst_5_0_n2 , AddKeyXOR_XORInst_5_2_n2 ,
         AddKeyXOR_XORInst_6_0_n2 , AddKeyXOR_XORInst_6_2_n2 ,
         AddKeyXOR_XORInst_7_0_n2 , AddKeyXOR_XORInst_7_2_n2 ,
         AddKeyXOR_XORInst_8_0_n2 , AddKeyXOR_XORInst_8_2_n2 ,
         AddKeyXOR_XORInst_9_0_n2 , AddKeyXOR_XORInst_9_2_n2 ,
         AddKeyXOR_XORInst_10_0_n2 , AddKeyXOR_XORInst_10_2_n2 ,
         AddKeyXOR_XORInst_11_0_n2 , AddKeyXOR_XORInst_11_2_n2 ,
         AddKeyXOR_XORInst_12_0_n2 , AddKeyXOR_XORInst_12_2_n2 ,
         AddKeyXOR_XORInst_13_0_n2 , AddKeyXOR_XORInst_13_2_n2 ,
         AddKeyXOR_XORInst_14_0_n2 , AddKeyXOR_XORInst_14_2_n2 ,
         AddKeyXOR_XORInst_15_0_n2 , AddKeyXOR_XORInst_15_2_n2 ,
         SubCellInst_LFInst_0_LFInst_0_n6 ,
         SubCellInst_LFInst_0_LFInst_0_n5 ,
         SubCellInst_LFInst_0_LFInst_0_n4 ,
         SubCellInst_LFInst_0_LFInst_1_n18 ,
         SubCellInst_LFInst_0_LFInst_1_n17 ,
         SubCellInst_LFInst_0_LFInst_1_n16 ,
         SubCellInst_LFInst_0_LFInst_1_n15 ,
         SubCellInst_LFInst_0_LFInst_1_n14 ,
         SubCellInst_LFInst_0_LFInst_1_n13 ,
         SubCellInst_LFInst_0_LFInst_1_n12 ,
         SubCellInst_LFInst_0_LFInst_1_n11 ,
         SubCellInst_LFInst_0_LFInst_1_n10 ,
         SubCellInst_LFInst_0_LFInst_2_n22 ,
         SubCellInst_LFInst_0_LFInst_2_n21 ,
         SubCellInst_LFInst_0_LFInst_2_n20 ,
         SubCellInst_LFInst_0_LFInst_2_n19 ,
         SubCellInst_LFInst_0_LFInst_2_n18 ,
         SubCellInst_LFInst_0_LFInst_2_n17 ,
         SubCellInst_LFInst_0_LFInst_2_n16 ,
         SubCellInst_LFInst_0_LFInst_2_n15 ,
         SubCellInst_LFInst_0_LFInst_3_n16 ,
         SubCellInst_LFInst_0_LFInst_3_n15 ,
         SubCellInst_LFInst_0_LFInst_3_n14 ,
         SubCellInst_LFInst_0_LFInst_3_n13 ,
         SubCellInst_LFInst_0_LFInst_3_n12 ,
         SubCellInst_LFInst_0_LFInst_3_n11 ,
         SubCellInst_LFInst_1_LFInst_0_n6 ,
         SubCellInst_LFInst_1_LFInst_0_n5 ,
         SubCellInst_LFInst_1_LFInst_0_n4 ,
         SubCellInst_LFInst_1_LFInst_1_n18 ,
         SubCellInst_LFInst_1_LFInst_1_n17 ,
         SubCellInst_LFInst_1_LFInst_1_n16 ,
         SubCellInst_LFInst_1_LFInst_1_n15 ,
         SubCellInst_LFInst_1_LFInst_1_n14 ,
         SubCellInst_LFInst_1_LFInst_1_n13 ,
         SubCellInst_LFInst_1_LFInst_1_n12 ,
         SubCellInst_LFInst_1_LFInst_1_n11 ,
         SubCellInst_LFInst_1_LFInst_1_n10 ,
         SubCellInst_LFInst_1_LFInst_2_n22 ,
         SubCellInst_LFInst_1_LFInst_2_n21 ,
         SubCellInst_LFInst_1_LFInst_2_n20 ,
         SubCellInst_LFInst_1_LFInst_2_n19 ,
         SubCellInst_LFInst_1_LFInst_2_n18 ,
         SubCellInst_LFInst_1_LFInst_2_n17 ,
         SubCellInst_LFInst_1_LFInst_2_n16 ,
         SubCellInst_LFInst_1_LFInst_2_n15 ,
         SubCellInst_LFInst_1_LFInst_3_n16 ,
         SubCellInst_LFInst_1_LFInst_3_n15 ,
         SubCellInst_LFInst_1_LFInst_3_n14 ,
         SubCellInst_LFInst_1_LFInst_3_n13 ,
         SubCellInst_LFInst_1_LFInst_3_n12 ,
         SubCellInst_LFInst_1_LFInst_3_n11 ,
         SubCellInst_LFInst_2_LFInst_0_n6 ,
         SubCellInst_LFInst_2_LFInst_0_n5 ,
         SubCellInst_LFInst_2_LFInst_0_n4 ,
         SubCellInst_LFInst_2_LFInst_1_n18 ,
         SubCellInst_LFInst_2_LFInst_1_n17 ,
         SubCellInst_LFInst_2_LFInst_1_n16 ,
         SubCellInst_LFInst_2_LFInst_1_n15 ,
         SubCellInst_LFInst_2_LFInst_1_n14 ,
         SubCellInst_LFInst_2_LFInst_1_n13 ,
         SubCellInst_LFInst_2_LFInst_1_n12 ,
         SubCellInst_LFInst_2_LFInst_1_n11 ,
         SubCellInst_LFInst_2_LFInst_1_n10 ,
         SubCellInst_LFInst_2_LFInst_2_n22 ,
         SubCellInst_LFInst_2_LFInst_2_n21 ,
         SubCellInst_LFInst_2_LFInst_2_n20 ,
         SubCellInst_LFInst_2_LFInst_2_n19 ,
         SubCellInst_LFInst_2_LFInst_2_n18 ,
         SubCellInst_LFInst_2_LFInst_2_n17 ,
         SubCellInst_LFInst_2_LFInst_2_n16 ,
         SubCellInst_LFInst_2_LFInst_2_n15 ,
         SubCellInst_LFInst_2_LFInst_3_n16 ,
         SubCellInst_LFInst_2_LFInst_3_n15 ,
         SubCellInst_LFInst_2_LFInst_3_n14 ,
         SubCellInst_LFInst_2_LFInst_3_n13 ,
         SubCellInst_LFInst_2_LFInst_3_n12 ,
         SubCellInst_LFInst_2_LFInst_3_n11 ,
         SubCellInst_LFInst_3_LFInst_0_n6 ,
         SubCellInst_LFInst_3_LFInst_0_n5 ,
         SubCellInst_LFInst_3_LFInst_0_n4 ,
         SubCellInst_LFInst_3_LFInst_1_n18 ,
         SubCellInst_LFInst_3_LFInst_1_n17 ,
         SubCellInst_LFInst_3_LFInst_1_n16 ,
         SubCellInst_LFInst_3_LFInst_1_n15 ,
         SubCellInst_LFInst_3_LFInst_1_n14 ,
         SubCellInst_LFInst_3_LFInst_1_n13 ,
         SubCellInst_LFInst_3_LFInst_1_n12 ,
         SubCellInst_LFInst_3_LFInst_1_n11 ,
         SubCellInst_LFInst_3_LFInst_1_n10 ,
         SubCellInst_LFInst_3_LFInst_2_n22 ,
         SubCellInst_LFInst_3_LFInst_2_n21 ,
         SubCellInst_LFInst_3_LFInst_2_n20 ,
         SubCellInst_LFInst_3_LFInst_2_n19 ,
         SubCellInst_LFInst_3_LFInst_2_n18 ,
         SubCellInst_LFInst_3_LFInst_2_n17 ,
         SubCellInst_LFInst_3_LFInst_2_n16 ,
         SubCellInst_LFInst_3_LFInst_2_n15 ,
         SubCellInst_LFInst_3_LFInst_3_n16 ,
         SubCellInst_LFInst_3_LFInst_3_n15 ,
         SubCellInst_LFInst_3_LFInst_3_n14 ,
         SubCellInst_LFInst_3_LFInst_3_n13 ,
         SubCellInst_LFInst_3_LFInst_3_n12 ,
         SubCellInst_LFInst_3_LFInst_3_n11 ,
         SubCellInst_LFInst_4_LFInst_0_n6 ,
         SubCellInst_LFInst_4_LFInst_0_n5 ,
         SubCellInst_LFInst_4_LFInst_0_n4 ,
         SubCellInst_LFInst_4_LFInst_1_n18 ,
         SubCellInst_LFInst_4_LFInst_1_n17 ,
         SubCellInst_LFInst_4_LFInst_1_n16 ,
         SubCellInst_LFInst_4_LFInst_1_n15 ,
         SubCellInst_LFInst_4_LFInst_1_n14 ,
         SubCellInst_LFInst_4_LFInst_1_n13 ,
         SubCellInst_LFInst_4_LFInst_1_n12 ,
         SubCellInst_LFInst_4_LFInst_1_n11 ,
         SubCellInst_LFInst_4_LFInst_1_n10 ,
         SubCellInst_LFInst_4_LFInst_2_n22 ,
         SubCellInst_LFInst_4_LFInst_2_n21 ,
         SubCellInst_LFInst_4_LFInst_2_n20 ,
         SubCellInst_LFInst_4_LFInst_2_n19 ,
         SubCellInst_LFInst_4_LFInst_2_n18 ,
         SubCellInst_LFInst_4_LFInst_2_n17 ,
         SubCellInst_LFInst_4_LFInst_2_n16 ,
         SubCellInst_LFInst_4_LFInst_2_n15 ,
         SubCellInst_LFInst_4_LFInst_3_n16 ,
         SubCellInst_LFInst_4_LFInst_3_n15 ,
         SubCellInst_LFInst_4_LFInst_3_n14 ,
         SubCellInst_LFInst_4_LFInst_3_n13 ,
         SubCellInst_LFInst_4_LFInst_3_n12 ,
         SubCellInst_LFInst_4_LFInst_3_n11 ,
         SubCellInst_LFInst_5_LFInst_0_n6 ,
         SubCellInst_LFInst_5_LFInst_0_n5 ,
         SubCellInst_LFInst_5_LFInst_0_n4 ,
         SubCellInst_LFInst_5_LFInst_1_n18 ,
         SubCellInst_LFInst_5_LFInst_1_n17 ,
         SubCellInst_LFInst_5_LFInst_1_n16 ,
         SubCellInst_LFInst_5_LFInst_1_n15 ,
         SubCellInst_LFInst_5_LFInst_1_n14 ,
         SubCellInst_LFInst_5_LFInst_1_n13 ,
         SubCellInst_LFInst_5_LFInst_1_n12 ,
         SubCellInst_LFInst_5_LFInst_1_n11 ,
         SubCellInst_LFInst_5_LFInst_1_n10 ,
         SubCellInst_LFInst_5_LFInst_2_n22 ,
         SubCellInst_LFInst_5_LFInst_2_n21 ,
         SubCellInst_LFInst_5_LFInst_2_n20 ,
         SubCellInst_LFInst_5_LFInst_2_n19 ,
         SubCellInst_LFInst_5_LFInst_2_n18 ,
         SubCellInst_LFInst_5_LFInst_2_n17 ,
         SubCellInst_LFInst_5_LFInst_2_n16 ,
         SubCellInst_LFInst_5_LFInst_2_n15 ,
         SubCellInst_LFInst_5_LFInst_3_n16 ,
         SubCellInst_LFInst_5_LFInst_3_n15 ,
         SubCellInst_LFInst_5_LFInst_3_n14 ,
         SubCellInst_LFInst_5_LFInst_3_n13 ,
         SubCellInst_LFInst_5_LFInst_3_n12 ,
         SubCellInst_LFInst_5_LFInst_3_n11 ,
         SubCellInst_LFInst_6_LFInst_0_n6 ,
         SubCellInst_LFInst_6_LFInst_0_n5 ,
         SubCellInst_LFInst_6_LFInst_0_n4 ,
         SubCellInst_LFInst_6_LFInst_1_n18 ,
         SubCellInst_LFInst_6_LFInst_1_n17 ,
         SubCellInst_LFInst_6_LFInst_1_n16 ,
         SubCellInst_LFInst_6_LFInst_1_n15 ,
         SubCellInst_LFInst_6_LFInst_1_n14 ,
         SubCellInst_LFInst_6_LFInst_1_n13 ,
         SubCellInst_LFInst_6_LFInst_1_n12 ,
         SubCellInst_LFInst_6_LFInst_1_n11 ,
         SubCellInst_LFInst_6_LFInst_1_n10 ,
         SubCellInst_LFInst_6_LFInst_2_n22 ,
         SubCellInst_LFInst_6_LFInst_2_n21 ,
         SubCellInst_LFInst_6_LFInst_2_n20 ,
         SubCellInst_LFInst_6_LFInst_2_n19 ,
         SubCellInst_LFInst_6_LFInst_2_n18 ,
         SubCellInst_LFInst_6_LFInst_2_n17 ,
         SubCellInst_LFInst_6_LFInst_2_n16 ,
         SubCellInst_LFInst_6_LFInst_2_n15 ,
         SubCellInst_LFInst_6_LFInst_3_n16 ,
         SubCellInst_LFInst_6_LFInst_3_n15 ,
         SubCellInst_LFInst_6_LFInst_3_n14 ,
         SubCellInst_LFInst_6_LFInst_3_n13 ,
         SubCellInst_LFInst_6_LFInst_3_n12 ,
         SubCellInst_LFInst_6_LFInst_3_n11 ,
         SubCellInst_LFInst_7_LFInst_0_n6 ,
         SubCellInst_LFInst_7_LFInst_0_n5 ,
         SubCellInst_LFInst_7_LFInst_0_n4 ,
         SubCellInst_LFInst_7_LFInst_1_n18 ,
         SubCellInst_LFInst_7_LFInst_1_n17 ,
         SubCellInst_LFInst_7_LFInst_1_n16 ,
         SubCellInst_LFInst_7_LFInst_1_n15 ,
         SubCellInst_LFInst_7_LFInst_1_n14 ,
         SubCellInst_LFInst_7_LFInst_1_n13 ,
         SubCellInst_LFInst_7_LFInst_1_n12 ,
         SubCellInst_LFInst_7_LFInst_1_n11 ,
         SubCellInst_LFInst_7_LFInst_1_n10 ,
         SubCellInst_LFInst_7_LFInst_2_n22 ,
         SubCellInst_LFInst_7_LFInst_2_n21 ,
         SubCellInst_LFInst_7_LFInst_2_n20 ,
         SubCellInst_LFInst_7_LFInst_2_n19 ,
         SubCellInst_LFInst_7_LFInst_2_n18 ,
         SubCellInst_LFInst_7_LFInst_2_n17 ,
         SubCellInst_LFInst_7_LFInst_2_n16 ,
         SubCellInst_LFInst_7_LFInst_2_n15 ,
         SubCellInst_LFInst_7_LFInst_3_n16 ,
         SubCellInst_LFInst_7_LFInst_3_n15 ,
         SubCellInst_LFInst_7_LFInst_3_n14 ,
         SubCellInst_LFInst_7_LFInst_3_n13 ,
         SubCellInst_LFInst_7_LFInst_3_n12 ,
         SubCellInst_LFInst_7_LFInst_3_n11 ,
         SubCellInst_LFInst_8_LFInst_0_n6 ,
         SubCellInst_LFInst_8_LFInst_0_n5 ,
         SubCellInst_LFInst_8_LFInst_0_n4 ,
         SubCellInst_LFInst_8_LFInst_1_n18 ,
         SubCellInst_LFInst_8_LFInst_1_n17 ,
         SubCellInst_LFInst_8_LFInst_1_n16 ,
         SubCellInst_LFInst_8_LFInst_1_n15 ,
         SubCellInst_LFInst_8_LFInst_1_n14 ,
         SubCellInst_LFInst_8_LFInst_1_n13 ,
         SubCellInst_LFInst_8_LFInst_1_n12 ,
         SubCellInst_LFInst_8_LFInst_1_n11 ,
         SubCellInst_LFInst_8_LFInst_1_n10 ,
         SubCellInst_LFInst_8_LFInst_2_n22 ,
         SubCellInst_LFInst_8_LFInst_2_n21 ,
         SubCellInst_LFInst_8_LFInst_2_n20 ,
         SubCellInst_LFInst_8_LFInst_2_n19 ,
         SubCellInst_LFInst_8_LFInst_2_n18 ,
         SubCellInst_LFInst_8_LFInst_2_n17 ,
         SubCellInst_LFInst_8_LFInst_2_n16 ,
         SubCellInst_LFInst_8_LFInst_2_n15 ,
         SubCellInst_LFInst_8_LFInst_3_n16 ,
         SubCellInst_LFInst_8_LFInst_3_n15 ,
         SubCellInst_LFInst_8_LFInst_3_n14 ,
         SubCellInst_LFInst_8_LFInst_3_n13 ,
         SubCellInst_LFInst_8_LFInst_3_n12 ,
         SubCellInst_LFInst_8_LFInst_3_n11 ,
         SubCellInst_LFInst_9_LFInst_0_n6 ,
         SubCellInst_LFInst_9_LFInst_0_n5 ,
         SubCellInst_LFInst_9_LFInst_0_n4 ,
         SubCellInst_LFInst_9_LFInst_1_n18 ,
         SubCellInst_LFInst_9_LFInst_1_n17 ,
         SubCellInst_LFInst_9_LFInst_1_n16 ,
         SubCellInst_LFInst_9_LFInst_1_n15 ,
         SubCellInst_LFInst_9_LFInst_1_n14 ,
         SubCellInst_LFInst_9_LFInst_1_n13 ,
         SubCellInst_LFInst_9_LFInst_1_n12 ,
         SubCellInst_LFInst_9_LFInst_1_n11 ,
         SubCellInst_LFInst_9_LFInst_1_n10 ,
         SubCellInst_LFInst_9_LFInst_2_n22 ,
         SubCellInst_LFInst_9_LFInst_2_n21 ,
         SubCellInst_LFInst_9_LFInst_2_n20 ,
         SubCellInst_LFInst_9_LFInst_2_n19 ,
         SubCellInst_LFInst_9_LFInst_2_n18 ,
         SubCellInst_LFInst_9_LFInst_2_n17 ,
         SubCellInst_LFInst_9_LFInst_2_n16 ,
         SubCellInst_LFInst_9_LFInst_2_n15 ,
         SubCellInst_LFInst_9_LFInst_3_n16 ,
         SubCellInst_LFInst_9_LFInst_3_n15 ,
         SubCellInst_LFInst_9_LFInst_3_n14 ,
         SubCellInst_LFInst_9_LFInst_3_n13 ,
         SubCellInst_LFInst_9_LFInst_3_n12 ,
         SubCellInst_LFInst_9_LFInst_3_n11 ,
         SubCellInst_LFInst_10_LFInst_0_n6 ,
         SubCellInst_LFInst_10_LFInst_0_n5 ,
         SubCellInst_LFInst_10_LFInst_0_n4 ,
         SubCellInst_LFInst_10_LFInst_1_n18 ,
         SubCellInst_LFInst_10_LFInst_1_n17 ,
         SubCellInst_LFInst_10_LFInst_1_n16 ,
         SubCellInst_LFInst_10_LFInst_1_n15 ,
         SubCellInst_LFInst_10_LFInst_1_n14 ,
         SubCellInst_LFInst_10_LFInst_1_n13 ,
         SubCellInst_LFInst_10_LFInst_1_n12 ,
         SubCellInst_LFInst_10_LFInst_1_n11 ,
         SubCellInst_LFInst_10_LFInst_1_n10 ,
         SubCellInst_LFInst_10_LFInst_2_n22 ,
         SubCellInst_LFInst_10_LFInst_2_n21 ,
         SubCellInst_LFInst_10_LFInst_2_n20 ,
         SubCellInst_LFInst_10_LFInst_2_n19 ,
         SubCellInst_LFInst_10_LFInst_2_n18 ,
         SubCellInst_LFInst_10_LFInst_2_n17 ,
         SubCellInst_LFInst_10_LFInst_2_n16 ,
         SubCellInst_LFInst_10_LFInst_2_n15 ,
         SubCellInst_LFInst_10_LFInst_3_n16 ,
         SubCellInst_LFInst_10_LFInst_3_n15 ,
         SubCellInst_LFInst_10_LFInst_3_n14 ,
         SubCellInst_LFInst_10_LFInst_3_n13 ,
         SubCellInst_LFInst_10_LFInst_3_n12 ,
         SubCellInst_LFInst_10_LFInst_3_n11 ,
         SubCellInst_LFInst_11_LFInst_0_n6 ,
         SubCellInst_LFInst_11_LFInst_0_n5 ,
         SubCellInst_LFInst_11_LFInst_0_n4 ,
         SubCellInst_LFInst_11_LFInst_1_n18 ,
         SubCellInst_LFInst_11_LFInst_1_n17 ,
         SubCellInst_LFInst_11_LFInst_1_n16 ,
         SubCellInst_LFInst_11_LFInst_1_n15 ,
         SubCellInst_LFInst_11_LFInst_1_n14 ,
         SubCellInst_LFInst_11_LFInst_1_n13 ,
         SubCellInst_LFInst_11_LFInst_1_n12 ,
         SubCellInst_LFInst_11_LFInst_1_n11 ,
         SubCellInst_LFInst_11_LFInst_1_n10 ,
         SubCellInst_LFInst_11_LFInst_2_n22 ,
         SubCellInst_LFInst_11_LFInst_2_n21 ,
         SubCellInst_LFInst_11_LFInst_2_n20 ,
         SubCellInst_LFInst_11_LFInst_2_n19 ,
         SubCellInst_LFInst_11_LFInst_2_n18 ,
         SubCellInst_LFInst_11_LFInst_2_n17 ,
         SubCellInst_LFInst_11_LFInst_2_n16 ,
         SubCellInst_LFInst_11_LFInst_2_n15 ,
         SubCellInst_LFInst_11_LFInst_3_n16 ,
         SubCellInst_LFInst_11_LFInst_3_n15 ,
         SubCellInst_LFInst_11_LFInst_3_n14 ,
         SubCellInst_LFInst_11_LFInst_3_n13 ,
         SubCellInst_LFInst_11_LFInst_3_n12 ,
         SubCellInst_LFInst_11_LFInst_3_n11 ,
         SubCellInst_LFInst_12_LFInst_0_n6 ,
         SubCellInst_LFInst_12_LFInst_0_n5 ,
         SubCellInst_LFInst_12_LFInst_0_n4 ,
         SubCellInst_LFInst_12_LFInst_1_n18 ,
         SubCellInst_LFInst_12_LFInst_1_n17 ,
         SubCellInst_LFInst_12_LFInst_1_n16 ,
         SubCellInst_LFInst_12_LFInst_1_n15 ,
         SubCellInst_LFInst_12_LFInst_1_n14 ,
         SubCellInst_LFInst_12_LFInst_1_n13 ,
         SubCellInst_LFInst_12_LFInst_1_n12 ,
         SubCellInst_LFInst_12_LFInst_1_n11 ,
         SubCellInst_LFInst_12_LFInst_1_n10 ,
         SubCellInst_LFInst_12_LFInst_2_n22 ,
         SubCellInst_LFInst_12_LFInst_2_n21 ,
         SubCellInst_LFInst_12_LFInst_2_n20 ,
         SubCellInst_LFInst_12_LFInst_2_n19 ,
         SubCellInst_LFInst_12_LFInst_2_n18 ,
         SubCellInst_LFInst_12_LFInst_2_n17 ,
         SubCellInst_LFInst_12_LFInst_2_n16 ,
         SubCellInst_LFInst_12_LFInst_2_n15 ,
         SubCellInst_LFInst_12_LFInst_3_n16 ,
         SubCellInst_LFInst_12_LFInst_3_n15 ,
         SubCellInst_LFInst_12_LFInst_3_n14 ,
         SubCellInst_LFInst_12_LFInst_3_n13 ,
         SubCellInst_LFInst_12_LFInst_3_n12 ,
         SubCellInst_LFInst_12_LFInst_3_n11 ,
         SubCellInst_LFInst_13_LFInst_0_n6 ,
         SubCellInst_LFInst_13_LFInst_0_n5 ,
         SubCellInst_LFInst_13_LFInst_0_n4 ,
         SubCellInst_LFInst_13_LFInst_1_n18 ,
         SubCellInst_LFInst_13_LFInst_1_n17 ,
         SubCellInst_LFInst_13_LFInst_1_n16 ,
         SubCellInst_LFInst_13_LFInst_1_n15 ,
         SubCellInst_LFInst_13_LFInst_1_n14 ,
         SubCellInst_LFInst_13_LFInst_1_n13 ,
         SubCellInst_LFInst_13_LFInst_1_n12 ,
         SubCellInst_LFInst_13_LFInst_1_n11 ,
         SubCellInst_LFInst_13_LFInst_1_n10 ,
         SubCellInst_LFInst_13_LFInst_2_n22 ,
         SubCellInst_LFInst_13_LFInst_2_n21 ,
         SubCellInst_LFInst_13_LFInst_2_n20 ,
         SubCellInst_LFInst_13_LFInst_2_n19 ,
         SubCellInst_LFInst_13_LFInst_2_n18 ,
         SubCellInst_LFInst_13_LFInst_2_n17 ,
         SubCellInst_LFInst_13_LFInst_2_n16 ,
         SubCellInst_LFInst_13_LFInst_2_n15 ,
         SubCellInst_LFInst_13_LFInst_3_n16 ,
         SubCellInst_LFInst_13_LFInst_3_n15 ,
         SubCellInst_LFInst_13_LFInst_3_n14 ,
         SubCellInst_LFInst_13_LFInst_3_n13 ,
         SubCellInst_LFInst_13_LFInst_3_n12 ,
         SubCellInst_LFInst_13_LFInst_3_n11 ,
         SubCellInst_LFInst_14_LFInst_0_n6 ,
         SubCellInst_LFInst_14_LFInst_0_n5 ,
         SubCellInst_LFInst_14_LFInst_0_n4 ,
         SubCellInst_LFInst_14_LFInst_1_n18 ,
         SubCellInst_LFInst_14_LFInst_1_n17 ,
         SubCellInst_LFInst_14_LFInst_1_n16 ,
         SubCellInst_LFInst_14_LFInst_1_n15 ,
         SubCellInst_LFInst_14_LFInst_1_n14 ,
         SubCellInst_LFInst_14_LFInst_1_n13 ,
         SubCellInst_LFInst_14_LFInst_1_n12 ,
         SubCellInst_LFInst_14_LFInst_1_n11 ,
         SubCellInst_LFInst_14_LFInst_1_n10 ,
         SubCellInst_LFInst_14_LFInst_2_n22 ,
         SubCellInst_LFInst_14_LFInst_2_n21 ,
         SubCellInst_LFInst_14_LFInst_2_n20 ,
         SubCellInst_LFInst_14_LFInst_2_n19 ,
         SubCellInst_LFInst_14_LFInst_2_n18 ,
         SubCellInst_LFInst_14_LFInst_2_n17 ,
         SubCellInst_LFInst_14_LFInst_2_n16 ,
         SubCellInst_LFInst_14_LFInst_2_n15 ,
         SubCellInst_LFInst_14_LFInst_3_n16 ,
         SubCellInst_LFInst_14_LFInst_3_n15 ,
         SubCellInst_LFInst_14_LFInst_3_n14 ,
         SubCellInst_LFInst_14_LFInst_3_n13 ,
         SubCellInst_LFInst_14_LFInst_3_n12 ,
         SubCellInst_LFInst_14_LFInst_3_n11 ,
         SubCellInst_LFInst_15_LFInst_0_n6 ,
         SubCellInst_LFInst_15_LFInst_0_n5 ,
         SubCellInst_LFInst_15_LFInst_0_n4 ,
         SubCellInst_LFInst_15_LFInst_1_n18 ,
         SubCellInst_LFInst_15_LFInst_1_n17 ,
         SubCellInst_LFInst_15_LFInst_1_n16 ,
         SubCellInst_LFInst_15_LFInst_1_n15 ,
         SubCellInst_LFInst_15_LFInst_1_n14 ,
         SubCellInst_LFInst_15_LFInst_1_n13 ,
         SubCellInst_LFInst_15_LFInst_1_n12 ,
         SubCellInst_LFInst_15_LFInst_1_n11 ,
         SubCellInst_LFInst_15_LFInst_1_n10 ,
         SubCellInst_LFInst_15_LFInst_2_n22 ,
         SubCellInst_LFInst_15_LFInst_2_n21 ,
         SubCellInst_LFInst_15_LFInst_2_n20 ,
         SubCellInst_LFInst_15_LFInst_2_n19 ,
         SubCellInst_LFInst_15_LFInst_2_n18 ,
         SubCellInst_LFInst_15_LFInst_2_n17 ,
         SubCellInst_LFInst_15_LFInst_2_n16 ,
         SubCellInst_LFInst_15_LFInst_2_n15 ,
         SubCellInst_LFInst_15_LFInst_3_n16 ,
         SubCellInst_LFInst_15_LFInst_3_n15 ,
         SubCellInst_LFInst_15_LFInst_3_n14 ,
         SubCellInst_LFInst_15_LFInst_3_n13 ,
         SubCellInst_LFInst_15_LFInst_3_n12 ,
         SubCellInst_LFInst_15_LFInst_3_n11 , MCInst_MC0_v0_2Inst_0_n2 ,
         MCInst_MC0_v1_2Inst_0_n2 , MCInst_MC0_v2_3Inst_0_n4 ,
         MCInst_MC0_v2_3Inst_0_n3 , MCInst_MC0_v3_3Inst_0_n2 ,
         MCInst_MC0_v0_2Inst_1_n2 , MCInst_MC0_v2_1Inst_1_n2 ,
         MCInst_MC0_v2_2Inst_1_n4 , MCInst_MC0_v2_2Inst_1_n3 ,
         MCInst_MC0_v3_3Inst_1_n2 , MCInst_MC0_v1_1Inst_2_n2 ,
         MCInst_MC0_v1_2Inst_2_n2 , MCInst_MC0_v2_1Inst_2_n2 ,
         MCInst_MC0_v2_2Inst_2_n2 , MCInst_MC0_v3_1Inst_2_n2 ,
         MCInst_MC0_v1_2Inst_3_n4 , MCInst_MC0_v1_2Inst_3_n3 ,
         MCInst_MC0_v2_2Inst_3_n2 , MCInst_MC0_v2_3Inst_3_n2 ,
         MCInst_MC0_r0Inst_XORInst_0_0_n5 ,
         MCInst_MC0_r0Inst_XORInst_0_0_n4 ,
         MCInst_MC0_r0Inst_XORInst_0_1_n5 ,
         MCInst_MC0_r0Inst_XORInst_0_1_n4 ,
         MCInst_MC0_r0Inst_XORInst_0_2_n5 ,
         MCInst_MC0_r0Inst_XORInst_0_2_n4 ,
         MCInst_MC0_r0Inst_XORInst_0_3_n5 ,
         MCInst_MC0_r0Inst_XORInst_0_3_n4 ,
         MCInst_MC0_r1Inst_XORInst_0_0_n5 ,
         MCInst_MC0_r1Inst_XORInst_0_0_n4 ,
         MCInst_MC0_r1Inst_XORInst_0_1_n5 ,
         MCInst_MC0_r1Inst_XORInst_0_1_n4 ,
         MCInst_MC0_r1Inst_XORInst_0_2_n5 ,
         MCInst_MC0_r1Inst_XORInst_0_2_n4 ,
         MCInst_MC0_r1Inst_XORInst_0_3_n5 ,
         MCInst_MC0_r1Inst_XORInst_0_3_n4 ,
         MCInst_MC0_r2Inst_XORInst_0_0_n5 ,
         MCInst_MC0_r2Inst_XORInst_0_0_n4 ,
         MCInst_MC0_r2Inst_XORInst_0_1_n5 ,
         MCInst_MC0_r2Inst_XORInst_0_1_n4 ,
         MCInst_MC0_r2Inst_XORInst_0_2_n5 ,
         MCInst_MC0_r2Inst_XORInst_0_2_n4 ,
         MCInst_MC0_r2Inst_XORInst_0_3_n5 ,
         MCInst_MC0_r2Inst_XORInst_0_3_n4 ,
         MCInst_MC0_r3Inst_XORInst_0_0_n5 ,
         MCInst_MC0_r3Inst_XORInst_0_0_n4 ,
         MCInst_MC0_r3Inst_XORInst_0_1_n5 ,
         MCInst_MC0_r3Inst_XORInst_0_1_n4 ,
         MCInst_MC0_r3Inst_XORInst_0_2_n5 ,
         MCInst_MC0_r3Inst_XORInst_0_2_n4 ,
         MCInst_MC0_r3Inst_XORInst_0_3_n5 ,
         MCInst_MC0_r3Inst_XORInst_0_3_n4 , MCInst_MC1_v0_2Inst_0_n2 ,
         MCInst_MC1_v1_2Inst_0_n2 , MCInst_MC1_v2_3Inst_0_n4 ,
         MCInst_MC1_v2_3Inst_0_n3 , MCInst_MC1_v3_3Inst_0_n2 ,
         MCInst_MC1_v0_2Inst_1_n2 , MCInst_MC1_v2_1Inst_1_n2 ,
         MCInst_MC1_v2_2Inst_1_n4 , MCInst_MC1_v2_2Inst_1_n3 ,
         MCInst_MC1_v3_3Inst_1_n2 , MCInst_MC1_v1_1Inst_2_n2 ,
         MCInst_MC1_v1_2Inst_2_n2 , MCInst_MC1_v2_1Inst_2_n2 ,
         MCInst_MC1_v2_2Inst_2_n2 , MCInst_MC1_v3_1Inst_2_n2 ,
         MCInst_MC1_v1_2Inst_3_n4 , MCInst_MC1_v1_2Inst_3_n3 ,
         MCInst_MC1_v2_2Inst_3_n2 , MCInst_MC1_v2_3Inst_3_n2 ,
         MCInst_MC1_r0Inst_XORInst_0_0_n5 ,
         MCInst_MC1_r0Inst_XORInst_0_0_n4 ,
         MCInst_MC1_r0Inst_XORInst_0_1_n5 ,
         MCInst_MC1_r0Inst_XORInst_0_1_n4 ,
         MCInst_MC1_r0Inst_XORInst_0_2_n5 ,
         MCInst_MC1_r0Inst_XORInst_0_2_n4 ,
         MCInst_MC1_r0Inst_XORInst_0_3_n5 ,
         MCInst_MC1_r0Inst_XORInst_0_3_n4 ,
         MCInst_MC1_r1Inst_XORInst_0_0_n5 ,
         MCInst_MC1_r1Inst_XORInst_0_0_n4 ,
         MCInst_MC1_r1Inst_XORInst_0_1_n5 ,
         MCInst_MC1_r1Inst_XORInst_0_1_n4 ,
         MCInst_MC1_r1Inst_XORInst_0_2_n5 ,
         MCInst_MC1_r1Inst_XORInst_0_2_n4 ,
         MCInst_MC1_r1Inst_XORInst_0_3_n5 ,
         MCInst_MC1_r1Inst_XORInst_0_3_n4 ,
         MCInst_MC1_r2Inst_XORInst_0_0_n5 ,
         MCInst_MC1_r2Inst_XORInst_0_0_n4 ,
         MCInst_MC1_r2Inst_XORInst_0_1_n5 ,
         MCInst_MC1_r2Inst_XORInst_0_1_n4 ,
         MCInst_MC1_r2Inst_XORInst_0_2_n5 ,
         MCInst_MC1_r2Inst_XORInst_0_2_n4 ,
         MCInst_MC1_r2Inst_XORInst_0_3_n5 ,
         MCInst_MC1_r2Inst_XORInst_0_3_n4 ,
         MCInst_MC1_r3Inst_XORInst_0_0_n5 ,
         MCInst_MC1_r3Inst_XORInst_0_0_n4 ,
         MCInst_MC1_r3Inst_XORInst_0_1_n5 ,
         MCInst_MC1_r3Inst_XORInst_0_1_n4 ,
         MCInst_MC1_r3Inst_XORInst_0_2_n5 ,
         MCInst_MC1_r3Inst_XORInst_0_2_n4 ,
         MCInst_MC1_r3Inst_XORInst_0_3_n5 ,
         MCInst_MC1_r3Inst_XORInst_0_3_n4 , MCInst_MC2_v0_2Inst_0_n2 ,
         MCInst_MC2_v1_2Inst_0_n2 , MCInst_MC2_v2_3Inst_0_n4 ,
         MCInst_MC2_v2_3Inst_0_n3 , MCInst_MC2_v3_3Inst_0_n2 ,
         MCInst_MC2_v0_2Inst_1_n2 , MCInst_MC2_v2_1Inst_1_n2 ,
         MCInst_MC2_v2_2Inst_1_n4 , MCInst_MC2_v2_2Inst_1_n3 ,
         MCInst_MC2_v3_3Inst_1_n2 , MCInst_MC2_v1_1Inst_2_n2 ,
         MCInst_MC2_v1_2Inst_2_n2 , MCInst_MC2_v2_1Inst_2_n2 ,
         MCInst_MC2_v2_2Inst_2_n2 , MCInst_MC2_v3_1Inst_2_n2 ,
         MCInst_MC2_v1_2Inst_3_n4 , MCInst_MC2_v1_2Inst_3_n3 ,
         MCInst_MC2_v2_2Inst_3_n2 , MCInst_MC2_v2_3Inst_3_n2 ,
         MCInst_MC2_r0Inst_XORInst_0_0_n5 ,
         MCInst_MC2_r0Inst_XORInst_0_0_n4 ,
         MCInst_MC2_r0Inst_XORInst_0_1_n5 ,
         MCInst_MC2_r0Inst_XORInst_0_1_n4 ,
         MCInst_MC2_r0Inst_XORInst_0_2_n5 ,
         MCInst_MC2_r0Inst_XORInst_0_2_n4 ,
         MCInst_MC2_r0Inst_XORInst_0_3_n5 ,
         MCInst_MC2_r0Inst_XORInst_0_3_n4 ,
         MCInst_MC2_r1Inst_XORInst_0_0_n5 ,
         MCInst_MC2_r1Inst_XORInst_0_0_n4 ,
         MCInst_MC2_r1Inst_XORInst_0_1_n5 ,
         MCInst_MC2_r1Inst_XORInst_0_1_n4 ,
         MCInst_MC2_r1Inst_XORInst_0_2_n5 ,
         MCInst_MC2_r1Inst_XORInst_0_2_n4 ,
         MCInst_MC2_r1Inst_XORInst_0_3_n5 ,
         MCInst_MC2_r1Inst_XORInst_0_3_n4 ,
         MCInst_MC2_r2Inst_XORInst_0_0_n5 ,
         MCInst_MC2_r2Inst_XORInst_0_0_n4 ,
         MCInst_MC2_r2Inst_XORInst_0_1_n5 ,
         MCInst_MC2_r2Inst_XORInst_0_1_n4 ,
         MCInst_MC2_r2Inst_XORInst_0_2_n5 ,
         MCInst_MC2_r2Inst_XORInst_0_2_n4 ,
         MCInst_MC2_r2Inst_XORInst_0_3_n5 ,
         MCInst_MC2_r2Inst_XORInst_0_3_n4 ,
         MCInst_MC2_r3Inst_XORInst_0_0_n5 ,
         MCInst_MC2_r3Inst_XORInst_0_0_n4 ,
         MCInst_MC2_r3Inst_XORInst_0_1_n5 ,
         MCInst_MC2_r3Inst_XORInst_0_1_n4 ,
         MCInst_MC2_r3Inst_XORInst_0_2_n5 ,
         MCInst_MC2_r3Inst_XORInst_0_2_n4 ,
         MCInst_MC2_r3Inst_XORInst_0_3_n5 ,
         MCInst_MC2_r3Inst_XORInst_0_3_n4 , MCInst_MC3_v0_2Inst_0_n2 ,
         MCInst_MC3_v1_2Inst_0_n2 , MCInst_MC3_v2_3Inst_0_n4 ,
         MCInst_MC3_v2_3Inst_0_n3 , MCInst_MC3_v3_3Inst_0_n2 ,
         MCInst_MC3_v0_2Inst_1_n2 , MCInst_MC3_v2_1Inst_1_n2 ,
         MCInst_MC3_v2_2Inst_1_n4 , MCInst_MC3_v2_2Inst_1_n3 ,
         MCInst_MC3_v3_3Inst_1_n2 , MCInst_MC3_v1_1Inst_2_n2 ,
         MCInst_MC3_v1_2Inst_2_n2 , MCInst_MC3_v2_1Inst_2_n2 ,
         MCInst_MC3_v2_2Inst_2_n2 , MCInst_MC3_v3_1Inst_2_n2 ,
         MCInst_MC3_v1_2Inst_3_n4 , MCInst_MC3_v1_2Inst_3_n3 ,
         MCInst_MC3_v2_2Inst_3_n2 , MCInst_MC3_v2_3Inst_3_n2 ,
         MCInst_MC3_r0Inst_XORInst_0_0_n5 ,
         MCInst_MC3_r0Inst_XORInst_0_0_n4 ,
         MCInst_MC3_r0Inst_XORInst_0_1_n5 ,
         MCInst_MC3_r0Inst_XORInst_0_1_n4 ,
         MCInst_MC3_r0Inst_XORInst_0_2_n5 ,
         MCInst_MC3_r0Inst_XORInst_0_2_n4 ,
         MCInst_MC3_r0Inst_XORInst_0_3_n5 ,
         MCInst_MC3_r0Inst_XORInst_0_3_n4 ,
         MCInst_MC3_r1Inst_XORInst_0_0_n5 ,
         MCInst_MC3_r1Inst_XORInst_0_0_n4 ,
         MCInst_MC3_r1Inst_XORInst_0_1_n5 ,
         MCInst_MC3_r1Inst_XORInst_0_1_n4 ,
         MCInst_MC3_r1Inst_XORInst_0_2_n5 ,
         MCInst_MC3_r1Inst_XORInst_0_2_n4 ,
         MCInst_MC3_r1Inst_XORInst_0_3_n5 ,
         MCInst_MC3_r1Inst_XORInst_0_3_n4 ,
         MCInst_MC3_r2Inst_XORInst_0_0_n5 ,
         MCInst_MC3_r2Inst_XORInst_0_0_n4 ,
         MCInst_MC3_r2Inst_XORInst_0_1_n5 ,
         MCInst_MC3_r2Inst_XORInst_0_1_n4 ,
         MCInst_MC3_r2Inst_XORInst_0_2_n5 ,
         MCInst_MC3_r2Inst_XORInst_0_2_n4 ,
         MCInst_MC3_r2Inst_XORInst_0_3_n5 ,
         MCInst_MC3_r2Inst_XORInst_0_3_n4 ,
         MCInst_MC3_r3Inst_XORInst_0_0_n5 ,
         MCInst_MC3_r3Inst_XORInst_0_0_n4 ,
         MCInst_MC3_r3Inst_XORInst_0_1_n5 ,
         MCInst_MC3_r3Inst_XORInst_0_1_n4 ,
         MCInst_MC3_r3Inst_XORInst_0_2_n5 ,
         MCInst_MC3_r3Inst_XORInst_0_2_n4 ,
         MCInst_MC3_r3Inst_XORInst_0_3_n5 ,
         MCInst_MC3_r3Inst_XORInst_0_3_n4 ,
         SubCellInst2_LFInst_0_LFInst_0_n6 ,
         SubCellInst2_LFInst_0_LFInst_0_n5 ,
         SubCellInst2_LFInst_0_LFInst_0_n4 ,
         SubCellInst2_LFInst_0_LFInst_1_n18 ,
         SubCellInst2_LFInst_0_LFInst_1_n17 ,
         SubCellInst2_LFInst_0_LFInst_1_n16 ,
         SubCellInst2_LFInst_0_LFInst_1_n15 ,
         SubCellInst2_LFInst_0_LFInst_1_n14 ,
         SubCellInst2_LFInst_0_LFInst_1_n13 ,
         SubCellInst2_LFInst_0_LFInst_1_n12 ,
         SubCellInst2_LFInst_0_LFInst_1_n11 ,
         SubCellInst2_LFInst_0_LFInst_1_n10 ,
         SubCellInst2_LFInst_0_LFInst_2_n22 ,
         SubCellInst2_LFInst_0_LFInst_2_n21 ,
         SubCellInst2_LFInst_0_LFInst_2_n20 ,
         SubCellInst2_LFInst_0_LFInst_2_n19 ,
         SubCellInst2_LFInst_0_LFInst_2_n18 ,
         SubCellInst2_LFInst_0_LFInst_2_n17 ,
         SubCellInst2_LFInst_0_LFInst_2_n16 ,
         SubCellInst2_LFInst_0_LFInst_2_n15 ,
         SubCellInst2_LFInst_0_LFInst_3_n16 ,
         SubCellInst2_LFInst_0_LFInst_3_n15 ,
         SubCellInst2_LFInst_0_LFInst_3_n14 ,
         SubCellInst2_LFInst_0_LFInst_3_n13 ,
         SubCellInst2_LFInst_0_LFInst_3_n12 ,
         SubCellInst2_LFInst_0_LFInst_3_n11 ,
         SubCellInst2_LFInst_1_LFInst_0_n6 ,
         SubCellInst2_LFInst_1_LFInst_0_n5 ,
         SubCellInst2_LFInst_1_LFInst_0_n4 ,
         SubCellInst2_LFInst_1_LFInst_1_n18 ,
         SubCellInst2_LFInst_1_LFInst_1_n17 ,
         SubCellInst2_LFInst_1_LFInst_1_n16 ,
         SubCellInst2_LFInst_1_LFInst_1_n15 ,
         SubCellInst2_LFInst_1_LFInst_1_n14 ,
         SubCellInst2_LFInst_1_LFInst_1_n13 ,
         SubCellInst2_LFInst_1_LFInst_1_n12 ,
         SubCellInst2_LFInst_1_LFInst_1_n11 ,
         SubCellInst2_LFInst_1_LFInst_1_n10 ,
         SubCellInst2_LFInst_1_LFInst_2_n22 ,
         SubCellInst2_LFInst_1_LFInst_2_n21 ,
         SubCellInst2_LFInst_1_LFInst_2_n20 ,
         SubCellInst2_LFInst_1_LFInst_2_n19 ,
         SubCellInst2_LFInst_1_LFInst_2_n18 ,
         SubCellInst2_LFInst_1_LFInst_2_n17 ,
         SubCellInst2_LFInst_1_LFInst_2_n16 ,
         SubCellInst2_LFInst_1_LFInst_2_n15 ,
         SubCellInst2_LFInst_1_LFInst_3_n16 ,
         SubCellInst2_LFInst_1_LFInst_3_n15 ,
         SubCellInst2_LFInst_1_LFInst_3_n14 ,
         SubCellInst2_LFInst_1_LFInst_3_n13 ,
         SubCellInst2_LFInst_1_LFInst_3_n12 ,
         SubCellInst2_LFInst_1_LFInst_3_n11 ,
         SubCellInst2_LFInst_2_LFInst_0_n6 ,
         SubCellInst2_LFInst_2_LFInst_0_n5 ,
         SubCellInst2_LFInst_2_LFInst_0_n4 ,
         SubCellInst2_LFInst_2_LFInst_1_n18 ,
         SubCellInst2_LFInst_2_LFInst_1_n17 ,
         SubCellInst2_LFInst_2_LFInst_1_n16 ,
         SubCellInst2_LFInst_2_LFInst_1_n15 ,
         SubCellInst2_LFInst_2_LFInst_1_n14 ,
         SubCellInst2_LFInst_2_LFInst_1_n13 ,
         SubCellInst2_LFInst_2_LFInst_1_n12 ,
         SubCellInst2_LFInst_2_LFInst_1_n11 ,
         SubCellInst2_LFInst_2_LFInst_1_n10 ,
         SubCellInst2_LFInst_2_LFInst_2_n22 ,
         SubCellInst2_LFInst_2_LFInst_2_n21 ,
         SubCellInst2_LFInst_2_LFInst_2_n20 ,
         SubCellInst2_LFInst_2_LFInst_2_n19 ,
         SubCellInst2_LFInst_2_LFInst_2_n18 ,
         SubCellInst2_LFInst_2_LFInst_2_n17 ,
         SubCellInst2_LFInst_2_LFInst_2_n16 ,
         SubCellInst2_LFInst_2_LFInst_2_n15 ,
         SubCellInst2_LFInst_2_LFInst_3_n16 ,
         SubCellInst2_LFInst_2_LFInst_3_n15 ,
         SubCellInst2_LFInst_2_LFInst_3_n14 ,
         SubCellInst2_LFInst_2_LFInst_3_n13 ,
         SubCellInst2_LFInst_2_LFInst_3_n12 ,
         SubCellInst2_LFInst_2_LFInst_3_n11 ,
         SubCellInst2_LFInst_3_LFInst_0_n6 ,
         SubCellInst2_LFInst_3_LFInst_0_n5 ,
         SubCellInst2_LFInst_3_LFInst_0_n4 ,
         SubCellInst2_LFInst_3_LFInst_1_n18 ,
         SubCellInst2_LFInst_3_LFInst_1_n17 ,
         SubCellInst2_LFInst_3_LFInst_1_n16 ,
         SubCellInst2_LFInst_3_LFInst_1_n15 ,
         SubCellInst2_LFInst_3_LFInst_1_n14 ,
         SubCellInst2_LFInst_3_LFInst_1_n13 ,
         SubCellInst2_LFInst_3_LFInst_1_n12 ,
         SubCellInst2_LFInst_3_LFInst_1_n11 ,
         SubCellInst2_LFInst_3_LFInst_1_n10 ,
         SubCellInst2_LFInst_3_LFInst_2_n22 ,
         SubCellInst2_LFInst_3_LFInst_2_n21 ,
         SubCellInst2_LFInst_3_LFInst_2_n20 ,
         SubCellInst2_LFInst_3_LFInst_2_n19 ,
         SubCellInst2_LFInst_3_LFInst_2_n18 ,
         SubCellInst2_LFInst_3_LFInst_2_n17 ,
         SubCellInst2_LFInst_3_LFInst_2_n16 ,
         SubCellInst2_LFInst_3_LFInst_2_n15 ,
         SubCellInst2_LFInst_3_LFInst_3_n16 ,
         SubCellInst2_LFInst_3_LFInst_3_n15 ,
         SubCellInst2_LFInst_3_LFInst_3_n14 ,
         SubCellInst2_LFInst_3_LFInst_3_n13 ,
         SubCellInst2_LFInst_3_LFInst_3_n12 ,
         SubCellInst2_LFInst_3_LFInst_3_n11 ,
         SubCellInst2_LFInst_4_LFInst_0_n6 ,
         SubCellInst2_LFInst_4_LFInst_0_n5 ,
         SubCellInst2_LFInst_4_LFInst_0_n4 ,
         SubCellInst2_LFInst_4_LFInst_1_n18 ,
         SubCellInst2_LFInst_4_LFInst_1_n17 ,
         SubCellInst2_LFInst_4_LFInst_1_n16 ,
         SubCellInst2_LFInst_4_LFInst_1_n15 ,
         SubCellInst2_LFInst_4_LFInst_1_n14 ,
         SubCellInst2_LFInst_4_LFInst_1_n13 ,
         SubCellInst2_LFInst_4_LFInst_1_n12 ,
         SubCellInst2_LFInst_4_LFInst_1_n11 ,
         SubCellInst2_LFInst_4_LFInst_1_n10 ,
         SubCellInst2_LFInst_4_LFInst_2_n22 ,
         SubCellInst2_LFInst_4_LFInst_2_n21 ,
         SubCellInst2_LFInst_4_LFInst_2_n20 ,
         SubCellInst2_LFInst_4_LFInst_2_n19 ,
         SubCellInst2_LFInst_4_LFInst_2_n18 ,
         SubCellInst2_LFInst_4_LFInst_2_n17 ,
         SubCellInst2_LFInst_4_LFInst_2_n16 ,
         SubCellInst2_LFInst_4_LFInst_2_n15 ,
         SubCellInst2_LFInst_4_LFInst_3_n16 ,
         SubCellInst2_LFInst_4_LFInst_3_n15 ,
         SubCellInst2_LFInst_4_LFInst_3_n14 ,
         SubCellInst2_LFInst_4_LFInst_3_n13 ,
         SubCellInst2_LFInst_4_LFInst_3_n12 ,
         SubCellInst2_LFInst_4_LFInst_3_n11 ,
         SubCellInst2_LFInst_5_LFInst_0_n6 ,
         SubCellInst2_LFInst_5_LFInst_0_n5 ,
         SubCellInst2_LFInst_5_LFInst_0_n4 ,
         SubCellInst2_LFInst_5_LFInst_1_n18 ,
         SubCellInst2_LFInst_5_LFInst_1_n17 ,
         SubCellInst2_LFInst_5_LFInst_1_n16 ,
         SubCellInst2_LFInst_5_LFInst_1_n15 ,
         SubCellInst2_LFInst_5_LFInst_1_n14 ,
         SubCellInst2_LFInst_5_LFInst_1_n13 ,
         SubCellInst2_LFInst_5_LFInst_1_n12 ,
         SubCellInst2_LFInst_5_LFInst_1_n11 ,
         SubCellInst2_LFInst_5_LFInst_1_n10 ,
         SubCellInst2_LFInst_5_LFInst_2_n22 ,
         SubCellInst2_LFInst_5_LFInst_2_n21 ,
         SubCellInst2_LFInst_5_LFInst_2_n20 ,
         SubCellInst2_LFInst_5_LFInst_2_n19 ,
         SubCellInst2_LFInst_5_LFInst_2_n18 ,
         SubCellInst2_LFInst_5_LFInst_2_n17 ,
         SubCellInst2_LFInst_5_LFInst_2_n16 ,
         SubCellInst2_LFInst_5_LFInst_2_n15 ,
         SubCellInst2_LFInst_5_LFInst_3_n16 ,
         SubCellInst2_LFInst_5_LFInst_3_n15 ,
         SubCellInst2_LFInst_5_LFInst_3_n14 ,
         SubCellInst2_LFInst_5_LFInst_3_n13 ,
         SubCellInst2_LFInst_5_LFInst_3_n12 ,
         SubCellInst2_LFInst_5_LFInst_3_n11 ,
         SubCellInst2_LFInst_6_LFInst_0_n6 ,
         SubCellInst2_LFInst_6_LFInst_0_n5 ,
         SubCellInst2_LFInst_6_LFInst_0_n4 ,
         SubCellInst2_LFInst_6_LFInst_1_n18 ,
         SubCellInst2_LFInst_6_LFInst_1_n17 ,
         SubCellInst2_LFInst_6_LFInst_1_n16 ,
         SubCellInst2_LFInst_6_LFInst_1_n15 ,
         SubCellInst2_LFInst_6_LFInst_1_n14 ,
         SubCellInst2_LFInst_6_LFInst_1_n13 ,
         SubCellInst2_LFInst_6_LFInst_1_n12 ,
         SubCellInst2_LFInst_6_LFInst_1_n11 ,
         SubCellInst2_LFInst_6_LFInst_1_n10 ,
         SubCellInst2_LFInst_6_LFInst_2_n22 ,
         SubCellInst2_LFInst_6_LFInst_2_n21 ,
         SubCellInst2_LFInst_6_LFInst_2_n20 ,
         SubCellInst2_LFInst_6_LFInst_2_n19 ,
         SubCellInst2_LFInst_6_LFInst_2_n18 ,
         SubCellInst2_LFInst_6_LFInst_2_n17 ,
         SubCellInst2_LFInst_6_LFInst_2_n16 ,
         SubCellInst2_LFInst_6_LFInst_2_n15 ,
         SubCellInst2_LFInst_6_LFInst_3_n16 ,
         SubCellInst2_LFInst_6_LFInst_3_n15 ,
         SubCellInst2_LFInst_6_LFInst_3_n14 ,
         SubCellInst2_LFInst_6_LFInst_3_n13 ,
         SubCellInst2_LFInst_6_LFInst_3_n12 ,
         SubCellInst2_LFInst_6_LFInst_3_n11 ,
         SubCellInst2_LFInst_7_LFInst_0_n6 ,
         SubCellInst2_LFInst_7_LFInst_0_n5 ,
         SubCellInst2_LFInst_7_LFInst_0_n4 ,
         SubCellInst2_LFInst_7_LFInst_1_n18 ,
         SubCellInst2_LFInst_7_LFInst_1_n17 ,
         SubCellInst2_LFInst_7_LFInst_1_n16 ,
         SubCellInst2_LFInst_7_LFInst_1_n15 ,
         SubCellInst2_LFInst_7_LFInst_1_n14 ,
         SubCellInst2_LFInst_7_LFInst_1_n13 ,
         SubCellInst2_LFInst_7_LFInst_1_n12 ,
         SubCellInst2_LFInst_7_LFInst_1_n11 ,
         SubCellInst2_LFInst_7_LFInst_1_n10 ,
         SubCellInst2_LFInst_7_LFInst_2_n22 ,
         SubCellInst2_LFInst_7_LFInst_2_n21 ,
         SubCellInst2_LFInst_7_LFInst_2_n20 ,
         SubCellInst2_LFInst_7_LFInst_2_n19 ,
         SubCellInst2_LFInst_7_LFInst_2_n18 ,
         SubCellInst2_LFInst_7_LFInst_2_n17 ,
         SubCellInst2_LFInst_7_LFInst_2_n16 ,
         SubCellInst2_LFInst_7_LFInst_2_n15 ,
         SubCellInst2_LFInst_7_LFInst_3_n16 ,
         SubCellInst2_LFInst_7_LFInst_3_n15 ,
         SubCellInst2_LFInst_7_LFInst_3_n14 ,
         SubCellInst2_LFInst_7_LFInst_3_n13 ,
         SubCellInst2_LFInst_7_LFInst_3_n12 ,
         SubCellInst2_LFInst_7_LFInst_3_n11 ,
         SubCellInst2_LFInst_8_LFInst_0_n6 ,
         SubCellInst2_LFInst_8_LFInst_0_n5 ,
         SubCellInst2_LFInst_8_LFInst_0_n4 ,
         SubCellInst2_LFInst_8_LFInst_1_n18 ,
         SubCellInst2_LFInst_8_LFInst_1_n17 ,
         SubCellInst2_LFInst_8_LFInst_1_n16 ,
         SubCellInst2_LFInst_8_LFInst_1_n15 ,
         SubCellInst2_LFInst_8_LFInst_1_n14 ,
         SubCellInst2_LFInst_8_LFInst_1_n13 ,
         SubCellInst2_LFInst_8_LFInst_1_n12 ,
         SubCellInst2_LFInst_8_LFInst_1_n11 ,
         SubCellInst2_LFInst_8_LFInst_1_n10 ,
         SubCellInst2_LFInst_8_LFInst_2_n22 ,
         SubCellInst2_LFInst_8_LFInst_2_n21 ,
         SubCellInst2_LFInst_8_LFInst_2_n20 ,
         SubCellInst2_LFInst_8_LFInst_2_n19 ,
         SubCellInst2_LFInst_8_LFInst_2_n18 ,
         SubCellInst2_LFInst_8_LFInst_2_n17 ,
         SubCellInst2_LFInst_8_LFInst_2_n16 ,
         SubCellInst2_LFInst_8_LFInst_2_n15 ,
         SubCellInst2_LFInst_8_LFInst_3_n16 ,
         SubCellInst2_LFInst_8_LFInst_3_n15 ,
         SubCellInst2_LFInst_8_LFInst_3_n14 ,
         SubCellInst2_LFInst_8_LFInst_3_n13 ,
         SubCellInst2_LFInst_8_LFInst_3_n12 ,
         SubCellInst2_LFInst_8_LFInst_3_n11 ,
         SubCellInst2_LFInst_9_LFInst_0_n6 ,
         SubCellInst2_LFInst_9_LFInst_0_n5 ,
         SubCellInst2_LFInst_9_LFInst_0_n4 ,
         SubCellInst2_LFInst_9_LFInst_1_n18 ,
         SubCellInst2_LFInst_9_LFInst_1_n17 ,
         SubCellInst2_LFInst_9_LFInst_1_n16 ,
         SubCellInst2_LFInst_9_LFInst_1_n15 ,
         SubCellInst2_LFInst_9_LFInst_1_n14 ,
         SubCellInst2_LFInst_9_LFInst_1_n13 ,
         SubCellInst2_LFInst_9_LFInst_1_n12 ,
         SubCellInst2_LFInst_9_LFInst_1_n11 ,
         SubCellInst2_LFInst_9_LFInst_1_n10 ,
         SubCellInst2_LFInst_9_LFInst_2_n22 ,
         SubCellInst2_LFInst_9_LFInst_2_n21 ,
         SubCellInst2_LFInst_9_LFInst_2_n20 ,
         SubCellInst2_LFInst_9_LFInst_2_n19 ,
         SubCellInst2_LFInst_9_LFInst_2_n18 ,
         SubCellInst2_LFInst_9_LFInst_2_n17 ,
         SubCellInst2_LFInst_9_LFInst_2_n16 ,
         SubCellInst2_LFInst_9_LFInst_2_n15 ,
         SubCellInst2_LFInst_9_LFInst_3_n16 ,
         SubCellInst2_LFInst_9_LFInst_3_n15 ,
         SubCellInst2_LFInst_9_LFInst_3_n14 ,
         SubCellInst2_LFInst_9_LFInst_3_n13 ,
         SubCellInst2_LFInst_9_LFInst_3_n12 ,
         SubCellInst2_LFInst_9_LFInst_3_n11 ,
         SubCellInst2_LFInst_10_LFInst_0_n6 ,
         SubCellInst2_LFInst_10_LFInst_0_n5 ,
         SubCellInst2_LFInst_10_LFInst_0_n4 ,
         SubCellInst2_LFInst_10_LFInst_1_n18 ,
         SubCellInst2_LFInst_10_LFInst_1_n17 ,
         SubCellInst2_LFInst_10_LFInst_1_n16 ,
         SubCellInst2_LFInst_10_LFInst_1_n15 ,
         SubCellInst2_LFInst_10_LFInst_1_n14 ,
         SubCellInst2_LFInst_10_LFInst_1_n13 ,
         SubCellInst2_LFInst_10_LFInst_1_n12 ,
         SubCellInst2_LFInst_10_LFInst_1_n11 ,
         SubCellInst2_LFInst_10_LFInst_1_n10 ,
         SubCellInst2_LFInst_10_LFInst_2_n22 ,
         SubCellInst2_LFInst_10_LFInst_2_n21 ,
         SubCellInst2_LFInst_10_LFInst_2_n20 ,
         SubCellInst2_LFInst_10_LFInst_2_n19 ,
         SubCellInst2_LFInst_10_LFInst_2_n18 ,
         SubCellInst2_LFInst_10_LFInst_2_n17 ,
         SubCellInst2_LFInst_10_LFInst_2_n16 ,
         SubCellInst2_LFInst_10_LFInst_2_n15 ,
         SubCellInst2_LFInst_10_LFInst_3_n16 ,
         SubCellInst2_LFInst_10_LFInst_3_n15 ,
         SubCellInst2_LFInst_10_LFInst_3_n14 ,
         SubCellInst2_LFInst_10_LFInst_3_n13 ,
         SubCellInst2_LFInst_10_LFInst_3_n12 ,
         SubCellInst2_LFInst_10_LFInst_3_n11 ,
         SubCellInst2_LFInst_11_LFInst_0_n6 ,
         SubCellInst2_LFInst_11_LFInst_0_n5 ,
         SubCellInst2_LFInst_11_LFInst_0_n4 ,
         SubCellInst2_LFInst_11_LFInst_1_n18 ,
         SubCellInst2_LFInst_11_LFInst_1_n17 ,
         SubCellInst2_LFInst_11_LFInst_1_n16 ,
         SubCellInst2_LFInst_11_LFInst_1_n15 ,
         SubCellInst2_LFInst_11_LFInst_1_n14 ,
         SubCellInst2_LFInst_11_LFInst_1_n13 ,
         SubCellInst2_LFInst_11_LFInst_1_n12 ,
         SubCellInst2_LFInst_11_LFInst_1_n11 ,
         SubCellInst2_LFInst_11_LFInst_1_n10 ,
         SubCellInst2_LFInst_11_LFInst_2_n22 ,
         SubCellInst2_LFInst_11_LFInst_2_n21 ,
         SubCellInst2_LFInst_11_LFInst_2_n20 ,
         SubCellInst2_LFInst_11_LFInst_2_n19 ,
         SubCellInst2_LFInst_11_LFInst_2_n18 ,
         SubCellInst2_LFInst_11_LFInst_2_n17 ,
         SubCellInst2_LFInst_11_LFInst_2_n16 ,
         SubCellInst2_LFInst_11_LFInst_2_n15 ,
         SubCellInst2_LFInst_11_LFInst_3_n16 ,
         SubCellInst2_LFInst_11_LFInst_3_n15 ,
         SubCellInst2_LFInst_11_LFInst_3_n14 ,
         SubCellInst2_LFInst_11_LFInst_3_n13 ,
         SubCellInst2_LFInst_11_LFInst_3_n12 ,
         SubCellInst2_LFInst_11_LFInst_3_n11 ,
         SubCellInst2_LFInst_12_LFInst_0_n6 ,
         SubCellInst2_LFInst_12_LFInst_0_n5 ,
         SubCellInst2_LFInst_12_LFInst_0_n4 ,
         SubCellInst2_LFInst_12_LFInst_1_n18 ,
         SubCellInst2_LFInst_12_LFInst_1_n17 ,
         SubCellInst2_LFInst_12_LFInst_1_n16 ,
         SubCellInst2_LFInst_12_LFInst_1_n15 ,
         SubCellInst2_LFInst_12_LFInst_1_n14 ,
         SubCellInst2_LFInst_12_LFInst_1_n13 ,
         SubCellInst2_LFInst_12_LFInst_1_n12 ,
         SubCellInst2_LFInst_12_LFInst_1_n11 ,
         SubCellInst2_LFInst_12_LFInst_1_n10 ,
         SubCellInst2_LFInst_12_LFInst_2_n22 ,
         SubCellInst2_LFInst_12_LFInst_2_n21 ,
         SubCellInst2_LFInst_12_LFInst_2_n20 ,
         SubCellInst2_LFInst_12_LFInst_2_n19 ,
         SubCellInst2_LFInst_12_LFInst_2_n18 ,
         SubCellInst2_LFInst_12_LFInst_2_n17 ,
         SubCellInst2_LFInst_12_LFInst_2_n16 ,
         SubCellInst2_LFInst_12_LFInst_2_n15 ,
         SubCellInst2_LFInst_12_LFInst_3_n16 ,
         SubCellInst2_LFInst_12_LFInst_3_n15 ,
         SubCellInst2_LFInst_12_LFInst_3_n14 ,
         SubCellInst2_LFInst_12_LFInst_3_n13 ,
         SubCellInst2_LFInst_12_LFInst_3_n12 ,
         SubCellInst2_LFInst_12_LFInst_3_n11 ,
         SubCellInst2_LFInst_13_LFInst_0_n6 ,
         SubCellInst2_LFInst_13_LFInst_0_n5 ,
         SubCellInst2_LFInst_13_LFInst_0_n4 ,
         SubCellInst2_LFInst_13_LFInst_1_n18 ,
         SubCellInst2_LFInst_13_LFInst_1_n17 ,
         SubCellInst2_LFInst_13_LFInst_1_n16 ,
         SubCellInst2_LFInst_13_LFInst_1_n15 ,
         SubCellInst2_LFInst_13_LFInst_1_n14 ,
         SubCellInst2_LFInst_13_LFInst_1_n13 ,
         SubCellInst2_LFInst_13_LFInst_1_n12 ,
         SubCellInst2_LFInst_13_LFInst_1_n11 ,
         SubCellInst2_LFInst_13_LFInst_1_n10 ,
         SubCellInst2_LFInst_13_LFInst_2_n22 ,
         SubCellInst2_LFInst_13_LFInst_2_n21 ,
         SubCellInst2_LFInst_13_LFInst_2_n20 ,
         SubCellInst2_LFInst_13_LFInst_2_n19 ,
         SubCellInst2_LFInst_13_LFInst_2_n18 ,
         SubCellInst2_LFInst_13_LFInst_2_n17 ,
         SubCellInst2_LFInst_13_LFInst_2_n16 ,
         SubCellInst2_LFInst_13_LFInst_2_n15 ,
         SubCellInst2_LFInst_13_LFInst_3_n16 ,
         SubCellInst2_LFInst_13_LFInst_3_n15 ,
         SubCellInst2_LFInst_13_LFInst_3_n14 ,
         SubCellInst2_LFInst_13_LFInst_3_n13 ,
         SubCellInst2_LFInst_13_LFInst_3_n12 ,
         SubCellInst2_LFInst_13_LFInst_3_n11 ,
         SubCellInst2_LFInst_14_LFInst_0_n6 ,
         SubCellInst2_LFInst_14_LFInst_0_n5 ,
         SubCellInst2_LFInst_14_LFInst_0_n4 ,
         SubCellInst2_LFInst_14_LFInst_1_n18 ,
         SubCellInst2_LFInst_14_LFInst_1_n17 ,
         SubCellInst2_LFInst_14_LFInst_1_n16 ,
         SubCellInst2_LFInst_14_LFInst_1_n15 ,
         SubCellInst2_LFInst_14_LFInst_1_n14 ,
         SubCellInst2_LFInst_14_LFInst_1_n13 ,
         SubCellInst2_LFInst_14_LFInst_1_n12 ,
         SubCellInst2_LFInst_14_LFInst_1_n11 ,
         SubCellInst2_LFInst_14_LFInst_1_n10 ,
         SubCellInst2_LFInst_14_LFInst_2_n22 ,
         SubCellInst2_LFInst_14_LFInst_2_n21 ,
         SubCellInst2_LFInst_14_LFInst_2_n20 ,
         SubCellInst2_LFInst_14_LFInst_2_n19 ,
         SubCellInst2_LFInst_14_LFInst_2_n18 ,
         SubCellInst2_LFInst_14_LFInst_2_n17 ,
         SubCellInst2_LFInst_14_LFInst_2_n16 ,
         SubCellInst2_LFInst_14_LFInst_2_n15 ,
         SubCellInst2_LFInst_14_LFInst_3_n16 ,
         SubCellInst2_LFInst_14_LFInst_3_n15 ,
         SubCellInst2_LFInst_14_LFInst_3_n14 ,
         SubCellInst2_LFInst_14_LFInst_3_n13 ,
         SubCellInst2_LFInst_14_LFInst_3_n12 ,
         SubCellInst2_LFInst_14_LFInst_3_n11 ,
         SubCellInst2_LFInst_15_LFInst_0_n6 ,
         SubCellInst2_LFInst_15_LFInst_0_n5 ,
         SubCellInst2_LFInst_15_LFInst_0_n4 ,
         SubCellInst2_LFInst_15_LFInst_1_n18 ,
         SubCellInst2_LFInst_15_LFInst_1_n17 ,
         SubCellInst2_LFInst_15_LFInst_1_n16 ,
         SubCellInst2_LFInst_15_LFInst_1_n15 ,
         SubCellInst2_LFInst_15_LFInst_1_n14 ,
         SubCellInst2_LFInst_15_LFInst_1_n13 ,
         SubCellInst2_LFInst_15_LFInst_1_n12 ,
         SubCellInst2_LFInst_15_LFInst_1_n11 ,
         SubCellInst2_LFInst_15_LFInst_1_n10 ,
         SubCellInst2_LFInst_15_LFInst_2_n22 ,
         SubCellInst2_LFInst_15_LFInst_2_n21 ,
         SubCellInst2_LFInst_15_LFInst_2_n20 ,
         SubCellInst2_LFInst_15_LFInst_2_n19 ,
         SubCellInst2_LFInst_15_LFInst_2_n18 ,
         SubCellInst2_LFInst_15_LFInst_2_n17 ,
         SubCellInst2_LFInst_15_LFInst_2_n16 ,
         SubCellInst2_LFInst_15_LFInst_2_n15 ,
         SubCellInst2_LFInst_15_LFInst_3_n16 ,
         SubCellInst2_LFInst_15_LFInst_3_n15 ,
         SubCellInst2_LFInst_15_LFInst_3_n14 ,
         SubCellInst2_LFInst_15_LFInst_3_n13 ,
         SubCellInst2_LFInst_15_LFInst_3_n12 ,
         SubCellInst2_LFInst_15_LFInst_3_n11 , MCInst2_MC0_v0_2Inst_0_n2 ,
         MCInst2_MC0_v1_2Inst_0_n2 , MCInst2_MC0_v2_3Inst_0_n4 ,
         MCInst2_MC0_v2_3Inst_0_n3 , MCInst2_MC0_v3_3Inst_0_n2 ,
         MCInst2_MC0_v0_2Inst_1_n2 , MCInst2_MC0_v2_1Inst_1_n2 ,
         MCInst2_MC0_v2_2Inst_1_n4 , MCInst2_MC0_v2_2Inst_1_n3 ,
         MCInst2_MC0_v3_3Inst_1_n2 , MCInst2_MC0_v1_1Inst_2_n2 ,
         MCInst2_MC0_v1_2Inst_2_n2 , MCInst2_MC0_v2_1Inst_2_n2 ,
         MCInst2_MC0_v2_2Inst_2_n2 , MCInst2_MC0_v3_1Inst_2_n2 ,
         MCInst2_MC0_v1_2Inst_3_n4 , MCInst2_MC0_v1_2Inst_3_n3 ,
         MCInst2_MC0_v2_2Inst_3_n2 , MCInst2_MC0_v2_3Inst_3_n2 ,
         MCInst2_MC0_r0Inst_XORInst_0_0_n5 ,
         MCInst2_MC0_r0Inst_XORInst_0_0_n4 ,
         MCInst2_MC0_r0Inst_XORInst_0_1_n5 ,
         MCInst2_MC0_r0Inst_XORInst_0_1_n4 ,
         MCInst2_MC0_r0Inst_XORInst_0_2_n5 ,
         MCInst2_MC0_r0Inst_XORInst_0_2_n4 ,
         MCInst2_MC0_r0Inst_XORInst_0_3_n5 ,
         MCInst2_MC0_r0Inst_XORInst_0_3_n4 ,
         MCInst2_MC0_r1Inst_XORInst_0_0_n5 ,
         MCInst2_MC0_r1Inst_XORInst_0_0_n4 ,
         MCInst2_MC0_r1Inst_XORInst_0_1_n5 ,
         MCInst2_MC0_r1Inst_XORInst_0_1_n4 ,
         MCInst2_MC0_r1Inst_XORInst_0_2_n5 ,
         MCInst2_MC0_r1Inst_XORInst_0_2_n4 ,
         MCInst2_MC0_r1Inst_XORInst_0_3_n5 ,
         MCInst2_MC0_r1Inst_XORInst_0_3_n4 ,
         MCInst2_MC0_r2Inst_XORInst_0_0_n5 ,
         MCInst2_MC0_r2Inst_XORInst_0_0_n4 ,
         MCInst2_MC0_r2Inst_XORInst_0_1_n5 ,
         MCInst2_MC0_r2Inst_XORInst_0_1_n4 ,
         MCInst2_MC0_r2Inst_XORInst_0_2_n5 ,
         MCInst2_MC0_r2Inst_XORInst_0_2_n4 ,
         MCInst2_MC0_r2Inst_XORInst_0_3_n5 ,
         MCInst2_MC0_r2Inst_XORInst_0_3_n4 ,
         MCInst2_MC0_r3Inst_XORInst_0_0_n5 ,
         MCInst2_MC0_r3Inst_XORInst_0_0_n4 ,
         MCInst2_MC0_r3Inst_XORInst_0_1_n5 ,
         MCInst2_MC0_r3Inst_XORInst_0_1_n4 ,
         MCInst2_MC0_r3Inst_XORInst_0_2_n5 ,
         MCInst2_MC0_r3Inst_XORInst_0_2_n4 ,
         MCInst2_MC0_r3Inst_XORInst_0_3_n5 ,
         MCInst2_MC0_r3Inst_XORInst_0_3_n4 , MCInst2_MC1_v0_2Inst_0_n2 ,
         MCInst2_MC1_v1_2Inst_0_n2 , MCInst2_MC1_v2_3Inst_0_n4 ,
         MCInst2_MC1_v2_3Inst_0_n3 , MCInst2_MC1_v3_3Inst_0_n2 ,
         MCInst2_MC1_v0_2Inst_1_n2 , MCInst2_MC1_v2_1Inst_1_n2 ,
         MCInst2_MC1_v2_2Inst_1_n4 , MCInst2_MC1_v2_2Inst_1_n3 ,
         MCInst2_MC1_v3_3Inst_1_n2 , MCInst2_MC1_v1_1Inst_2_n2 ,
         MCInst2_MC1_v1_2Inst_2_n2 , MCInst2_MC1_v2_1Inst_2_n2 ,
         MCInst2_MC1_v2_2Inst_2_n2 , MCInst2_MC1_v3_1Inst_2_n2 ,
         MCInst2_MC1_v1_2Inst_3_n4 , MCInst2_MC1_v1_2Inst_3_n3 ,
         MCInst2_MC1_v2_2Inst_3_n2 , MCInst2_MC1_v2_3Inst_3_n2 ,
         MCInst2_MC1_r0Inst_XORInst_0_0_n5 ,
         MCInst2_MC1_r0Inst_XORInst_0_0_n4 ,
         MCInst2_MC1_r0Inst_XORInst_0_1_n5 ,
         MCInst2_MC1_r0Inst_XORInst_0_1_n4 ,
         MCInst2_MC1_r0Inst_XORInst_0_2_n5 ,
         MCInst2_MC1_r0Inst_XORInst_0_2_n4 ,
         MCInst2_MC1_r0Inst_XORInst_0_3_n5 ,
         MCInst2_MC1_r0Inst_XORInst_0_3_n4 ,
         MCInst2_MC1_r1Inst_XORInst_0_0_n5 ,
         MCInst2_MC1_r1Inst_XORInst_0_0_n4 ,
         MCInst2_MC1_r1Inst_XORInst_0_1_n5 ,
         MCInst2_MC1_r1Inst_XORInst_0_1_n4 ,
         MCInst2_MC1_r1Inst_XORInst_0_2_n5 ,
         MCInst2_MC1_r1Inst_XORInst_0_2_n4 ,
         MCInst2_MC1_r1Inst_XORInst_0_3_n5 ,
         MCInst2_MC1_r1Inst_XORInst_0_3_n4 ,
         MCInst2_MC1_r2Inst_XORInst_0_0_n5 ,
         MCInst2_MC1_r2Inst_XORInst_0_0_n4 ,
         MCInst2_MC1_r2Inst_XORInst_0_1_n5 ,
         MCInst2_MC1_r2Inst_XORInst_0_1_n4 ,
         MCInst2_MC1_r2Inst_XORInst_0_2_n5 ,
         MCInst2_MC1_r2Inst_XORInst_0_2_n4 ,
         MCInst2_MC1_r2Inst_XORInst_0_3_n5 ,
         MCInst2_MC1_r2Inst_XORInst_0_3_n4 ,
         MCInst2_MC1_r3Inst_XORInst_0_0_n5 ,
         MCInst2_MC1_r3Inst_XORInst_0_0_n4 ,
         MCInst2_MC1_r3Inst_XORInst_0_1_n5 ,
         MCInst2_MC1_r3Inst_XORInst_0_1_n4 ,
         MCInst2_MC1_r3Inst_XORInst_0_2_n5 ,
         MCInst2_MC1_r3Inst_XORInst_0_2_n4 ,
         MCInst2_MC1_r3Inst_XORInst_0_3_n5 ,
         MCInst2_MC1_r3Inst_XORInst_0_3_n4 , MCInst2_MC2_v0_2Inst_0_n2 ,
         MCInst2_MC2_v1_2Inst_0_n2 , MCInst2_MC2_v2_3Inst_0_n4 ,
         MCInst2_MC2_v2_3Inst_0_n3 , MCInst2_MC2_v3_3Inst_0_n2 ,
         MCInst2_MC2_v0_2Inst_1_n2 , MCInst2_MC2_v2_1Inst_1_n2 ,
         MCInst2_MC2_v2_2Inst_1_n4 , MCInst2_MC2_v2_2Inst_1_n3 ,
         MCInst2_MC2_v3_3Inst_1_n2 , MCInst2_MC2_v1_1Inst_2_n2 ,
         MCInst2_MC2_v1_2Inst_2_n2 , MCInst2_MC2_v2_1Inst_2_n2 ,
         MCInst2_MC2_v2_2Inst_2_n2 , MCInst2_MC2_v3_1Inst_2_n2 ,
         MCInst2_MC2_v1_2Inst_3_n4 , MCInst2_MC2_v1_2Inst_3_n3 ,
         MCInst2_MC2_v2_2Inst_3_n2 , MCInst2_MC2_v2_3Inst_3_n2 ,
         MCInst2_MC2_r0Inst_XORInst_0_0_n5 ,
         MCInst2_MC2_r0Inst_XORInst_0_0_n4 ,
         MCInst2_MC2_r0Inst_XORInst_0_1_n5 ,
         MCInst2_MC2_r0Inst_XORInst_0_1_n4 ,
         MCInst2_MC2_r0Inst_XORInst_0_2_n5 ,
         MCInst2_MC2_r0Inst_XORInst_0_2_n4 ,
         MCInst2_MC2_r0Inst_XORInst_0_3_n5 ,
         MCInst2_MC2_r0Inst_XORInst_0_3_n4 ,
         MCInst2_MC2_r1Inst_XORInst_0_0_n5 ,
         MCInst2_MC2_r1Inst_XORInst_0_0_n4 ,
         MCInst2_MC2_r1Inst_XORInst_0_1_n5 ,
         MCInst2_MC2_r1Inst_XORInst_0_1_n4 ,
         MCInst2_MC2_r1Inst_XORInst_0_2_n5 ,
         MCInst2_MC2_r1Inst_XORInst_0_2_n4 ,
         MCInst2_MC2_r1Inst_XORInst_0_3_n5 ,
         MCInst2_MC2_r1Inst_XORInst_0_3_n4 ,
         MCInst2_MC2_r2Inst_XORInst_0_0_n5 ,
         MCInst2_MC2_r2Inst_XORInst_0_0_n4 ,
         MCInst2_MC2_r2Inst_XORInst_0_1_n5 ,
         MCInst2_MC2_r2Inst_XORInst_0_1_n4 ,
         MCInst2_MC2_r2Inst_XORInst_0_2_n5 ,
         MCInst2_MC2_r2Inst_XORInst_0_2_n4 ,
         MCInst2_MC2_r2Inst_XORInst_0_3_n5 ,
         MCInst2_MC2_r2Inst_XORInst_0_3_n4 ,
         MCInst2_MC2_r3Inst_XORInst_0_0_n5 ,
         MCInst2_MC2_r3Inst_XORInst_0_0_n4 ,
         MCInst2_MC2_r3Inst_XORInst_0_1_n5 ,
         MCInst2_MC2_r3Inst_XORInst_0_1_n4 ,
         MCInst2_MC2_r3Inst_XORInst_0_2_n5 ,
         MCInst2_MC2_r3Inst_XORInst_0_2_n4 ,
         MCInst2_MC2_r3Inst_XORInst_0_3_n5 ,
         MCInst2_MC2_r3Inst_XORInst_0_3_n4 , MCInst2_MC3_v0_2Inst_0_n2 ,
         MCInst2_MC3_v1_2Inst_0_n2 , MCInst2_MC3_v2_3Inst_0_n4 ,
         MCInst2_MC3_v2_3Inst_0_n3 , MCInst2_MC3_v3_3Inst_0_n2 ,
         MCInst2_MC3_v0_2Inst_1_n2 , MCInst2_MC3_v2_1Inst_1_n2 ,
         MCInst2_MC3_v2_2Inst_1_n4 , MCInst2_MC3_v2_2Inst_1_n3 ,
         MCInst2_MC3_v3_3Inst_1_n2 , MCInst2_MC3_v1_1Inst_2_n2 ,
         MCInst2_MC3_v1_2Inst_2_n2 , MCInst2_MC3_v2_1Inst_2_n2 ,
         MCInst2_MC3_v2_2Inst_2_n2 , MCInst2_MC3_v3_1Inst_2_n2 ,
         MCInst2_MC3_v1_2Inst_3_n4 , MCInst2_MC3_v1_2Inst_3_n3 ,
         MCInst2_MC3_v2_2Inst_3_n2 , MCInst2_MC3_v2_3Inst_3_n2 ,
         MCInst2_MC3_r0Inst_XORInst_0_0_n5 ,
         MCInst2_MC3_r0Inst_XORInst_0_0_n4 ,
         MCInst2_MC3_r0Inst_XORInst_0_1_n5 ,
         MCInst2_MC3_r0Inst_XORInst_0_1_n4 ,
         MCInst2_MC3_r0Inst_XORInst_0_2_n5 ,
         MCInst2_MC3_r0Inst_XORInst_0_2_n4 ,
         MCInst2_MC3_r0Inst_XORInst_0_3_n5 ,
         MCInst2_MC3_r0Inst_XORInst_0_3_n4 ,
         MCInst2_MC3_r1Inst_XORInst_0_0_n5 ,
         MCInst2_MC3_r1Inst_XORInst_0_0_n4 ,
         MCInst2_MC3_r1Inst_XORInst_0_1_n5 ,
         MCInst2_MC3_r1Inst_XORInst_0_1_n4 ,
         MCInst2_MC3_r1Inst_XORInst_0_2_n5 ,
         MCInst2_MC3_r1Inst_XORInst_0_2_n4 ,
         MCInst2_MC3_r1Inst_XORInst_0_3_n5 ,
         MCInst2_MC3_r1Inst_XORInst_0_3_n4 ,
         MCInst2_MC3_r2Inst_XORInst_0_0_n5 ,
         MCInst2_MC3_r2Inst_XORInst_0_0_n4 ,
         MCInst2_MC3_r2Inst_XORInst_0_1_n5 ,
         MCInst2_MC3_r2Inst_XORInst_0_1_n4 ,
         MCInst2_MC3_r2Inst_XORInst_0_2_n5 ,
         MCInst2_MC3_r2Inst_XORInst_0_2_n4 ,
         MCInst2_MC3_r2Inst_XORInst_0_3_n5 ,
         MCInst2_MC3_r2Inst_XORInst_0_3_n4 ,
         MCInst2_MC3_r3Inst_XORInst_0_0_n5 ,
         MCInst2_MC3_r3Inst_XORInst_0_0_n4 ,
         MCInst2_MC3_r3Inst_XORInst_0_1_n5 ,
         MCInst2_MC3_r3Inst_XORInst_0_1_n4 ,
         MCInst2_MC3_r3Inst_XORInst_0_2_n5 ,
         MCInst2_MC3_r3Inst_XORInst_0_2_n4 ,
         MCInst2_MC3_r3Inst_XORInst_0_3_n5 ,
         MCInst2_MC3_r3Inst_XORInst_0_3_n4 ,
         SubCellInst3_LFInst_0_LFInst_0_n6 ,
         SubCellInst3_LFInst_0_LFInst_0_n5 ,
         SubCellInst3_LFInst_0_LFInst_0_n4 ,
         SubCellInst3_LFInst_0_LFInst_1_n18 ,
         SubCellInst3_LFInst_0_LFInst_1_n17 ,
         SubCellInst3_LFInst_0_LFInst_1_n16 ,
         SubCellInst3_LFInst_0_LFInst_1_n15 ,
         SubCellInst3_LFInst_0_LFInst_1_n14 ,
         SubCellInst3_LFInst_0_LFInst_1_n13 ,
         SubCellInst3_LFInst_0_LFInst_1_n12 ,
         SubCellInst3_LFInst_0_LFInst_1_n11 ,
         SubCellInst3_LFInst_0_LFInst_1_n10 ,
         SubCellInst3_LFInst_0_LFInst_2_n22 ,
         SubCellInst3_LFInst_0_LFInst_2_n21 ,
         SubCellInst3_LFInst_0_LFInst_2_n20 ,
         SubCellInst3_LFInst_0_LFInst_2_n19 ,
         SubCellInst3_LFInst_0_LFInst_2_n18 ,
         SubCellInst3_LFInst_0_LFInst_2_n17 ,
         SubCellInst3_LFInst_0_LFInst_2_n16 ,
         SubCellInst3_LFInst_0_LFInst_2_n15 ,
         SubCellInst3_LFInst_0_LFInst_3_n16 ,
         SubCellInst3_LFInst_0_LFInst_3_n15 ,
         SubCellInst3_LFInst_0_LFInst_3_n14 ,
         SubCellInst3_LFInst_0_LFInst_3_n13 ,
         SubCellInst3_LFInst_0_LFInst_3_n12 ,
         SubCellInst3_LFInst_0_LFInst_3_n11 ,
         SubCellInst3_LFInst_1_LFInst_0_n6 ,
         SubCellInst3_LFInst_1_LFInst_0_n5 ,
         SubCellInst3_LFInst_1_LFInst_0_n4 ,
         SubCellInst3_LFInst_1_LFInst_1_n18 ,
         SubCellInst3_LFInst_1_LFInst_1_n17 ,
         SubCellInst3_LFInst_1_LFInst_1_n16 ,
         SubCellInst3_LFInst_1_LFInst_1_n15 ,
         SubCellInst3_LFInst_1_LFInst_1_n14 ,
         SubCellInst3_LFInst_1_LFInst_1_n13 ,
         SubCellInst3_LFInst_1_LFInst_1_n12 ,
         SubCellInst3_LFInst_1_LFInst_1_n11 ,
         SubCellInst3_LFInst_1_LFInst_1_n10 ,
         SubCellInst3_LFInst_1_LFInst_2_n22 ,
         SubCellInst3_LFInst_1_LFInst_2_n21 ,
         SubCellInst3_LFInst_1_LFInst_2_n20 ,
         SubCellInst3_LFInst_1_LFInst_2_n19 ,
         SubCellInst3_LFInst_1_LFInst_2_n18 ,
         SubCellInst3_LFInst_1_LFInst_2_n17 ,
         SubCellInst3_LFInst_1_LFInst_2_n16 ,
         SubCellInst3_LFInst_1_LFInst_2_n15 ,
         SubCellInst3_LFInst_1_LFInst_3_n16 ,
         SubCellInst3_LFInst_1_LFInst_3_n15 ,
         SubCellInst3_LFInst_1_LFInst_3_n14 ,
         SubCellInst3_LFInst_1_LFInst_3_n13 ,
         SubCellInst3_LFInst_1_LFInst_3_n12 ,
         SubCellInst3_LFInst_1_LFInst_3_n11 ,
         SubCellInst3_LFInst_2_LFInst_0_n6 ,
         SubCellInst3_LFInst_2_LFInst_0_n5 ,
         SubCellInst3_LFInst_2_LFInst_0_n4 ,
         SubCellInst3_LFInst_2_LFInst_1_n18 ,
         SubCellInst3_LFInst_2_LFInst_1_n17 ,
         SubCellInst3_LFInst_2_LFInst_1_n16 ,
         SubCellInst3_LFInst_2_LFInst_1_n15 ,
         SubCellInst3_LFInst_2_LFInst_1_n14 ,
         SubCellInst3_LFInst_2_LFInst_1_n13 ,
         SubCellInst3_LFInst_2_LFInst_1_n12 ,
         SubCellInst3_LFInst_2_LFInst_1_n11 ,
         SubCellInst3_LFInst_2_LFInst_1_n10 ,
         SubCellInst3_LFInst_2_LFInst_2_n22 ,
         SubCellInst3_LFInst_2_LFInst_2_n21 ,
         SubCellInst3_LFInst_2_LFInst_2_n20 ,
         SubCellInst3_LFInst_2_LFInst_2_n19 ,
         SubCellInst3_LFInst_2_LFInst_2_n18 ,
         SubCellInst3_LFInst_2_LFInst_2_n17 ,
         SubCellInst3_LFInst_2_LFInst_2_n16 ,
         SubCellInst3_LFInst_2_LFInst_2_n15 ,
         SubCellInst3_LFInst_2_LFInst_3_n16 ,
         SubCellInst3_LFInst_2_LFInst_3_n15 ,
         SubCellInst3_LFInst_2_LFInst_3_n14 ,
         SubCellInst3_LFInst_2_LFInst_3_n13 ,
         SubCellInst3_LFInst_2_LFInst_3_n12 ,
         SubCellInst3_LFInst_2_LFInst_3_n11 ,
         SubCellInst3_LFInst_3_LFInst_0_n6 ,
         SubCellInst3_LFInst_3_LFInst_0_n5 ,
         SubCellInst3_LFInst_3_LFInst_0_n4 ,
         SubCellInst3_LFInst_3_LFInst_1_n18 ,
         SubCellInst3_LFInst_3_LFInst_1_n17 ,
         SubCellInst3_LFInst_3_LFInst_1_n16 ,
         SubCellInst3_LFInst_3_LFInst_1_n15 ,
         SubCellInst3_LFInst_3_LFInst_1_n14 ,
         SubCellInst3_LFInst_3_LFInst_1_n13 ,
         SubCellInst3_LFInst_3_LFInst_1_n12 ,
         SubCellInst3_LFInst_3_LFInst_1_n11 ,
         SubCellInst3_LFInst_3_LFInst_1_n10 ,
         SubCellInst3_LFInst_3_LFInst_2_n22 ,
         SubCellInst3_LFInst_3_LFInst_2_n21 ,
         SubCellInst3_LFInst_3_LFInst_2_n20 ,
         SubCellInst3_LFInst_3_LFInst_2_n19 ,
         SubCellInst3_LFInst_3_LFInst_2_n18 ,
         SubCellInst3_LFInst_3_LFInst_2_n17 ,
         SubCellInst3_LFInst_3_LFInst_2_n16 ,
         SubCellInst3_LFInst_3_LFInst_2_n15 ,
         SubCellInst3_LFInst_3_LFInst_3_n16 ,
         SubCellInst3_LFInst_3_LFInst_3_n15 ,
         SubCellInst3_LFInst_3_LFInst_3_n14 ,
         SubCellInst3_LFInst_3_LFInst_3_n13 ,
         SubCellInst3_LFInst_3_LFInst_3_n12 ,
         SubCellInst3_LFInst_3_LFInst_3_n11 ,
         SubCellInst3_LFInst_4_LFInst_0_n6 ,
         SubCellInst3_LFInst_4_LFInst_0_n5 ,
         SubCellInst3_LFInst_4_LFInst_0_n4 ,
         SubCellInst3_LFInst_4_LFInst_1_n18 ,
         SubCellInst3_LFInst_4_LFInst_1_n17 ,
         SubCellInst3_LFInst_4_LFInst_1_n16 ,
         SubCellInst3_LFInst_4_LFInst_1_n15 ,
         SubCellInst3_LFInst_4_LFInst_1_n14 ,
         SubCellInst3_LFInst_4_LFInst_1_n13 ,
         SubCellInst3_LFInst_4_LFInst_1_n12 ,
         SubCellInst3_LFInst_4_LFInst_1_n11 ,
         SubCellInst3_LFInst_4_LFInst_1_n10 ,
         SubCellInst3_LFInst_4_LFInst_2_n22 ,
         SubCellInst3_LFInst_4_LFInst_2_n21 ,
         SubCellInst3_LFInst_4_LFInst_2_n20 ,
         SubCellInst3_LFInst_4_LFInst_2_n19 ,
         SubCellInst3_LFInst_4_LFInst_2_n18 ,
         SubCellInst3_LFInst_4_LFInst_2_n17 ,
         SubCellInst3_LFInst_4_LFInst_2_n16 ,
         SubCellInst3_LFInst_4_LFInst_2_n15 ,
         SubCellInst3_LFInst_4_LFInst_3_n16 ,
         SubCellInst3_LFInst_4_LFInst_3_n15 ,
         SubCellInst3_LFInst_4_LFInst_3_n14 ,
         SubCellInst3_LFInst_4_LFInst_3_n13 ,
         SubCellInst3_LFInst_4_LFInst_3_n12 ,
         SubCellInst3_LFInst_4_LFInst_3_n11 ,
         SubCellInst3_LFInst_5_LFInst_0_n6 ,
         SubCellInst3_LFInst_5_LFInst_0_n5 ,
         SubCellInst3_LFInst_5_LFInst_0_n4 ,
         SubCellInst3_LFInst_5_LFInst_1_n18 ,
         SubCellInst3_LFInst_5_LFInst_1_n17 ,
         SubCellInst3_LFInst_5_LFInst_1_n16 ,
         SubCellInst3_LFInst_5_LFInst_1_n15 ,
         SubCellInst3_LFInst_5_LFInst_1_n14 ,
         SubCellInst3_LFInst_5_LFInst_1_n13 ,
         SubCellInst3_LFInst_5_LFInst_1_n12 ,
         SubCellInst3_LFInst_5_LFInst_1_n11 ,
         SubCellInst3_LFInst_5_LFInst_1_n10 ,
         SubCellInst3_LFInst_5_LFInst_2_n22 ,
         SubCellInst3_LFInst_5_LFInst_2_n21 ,
         SubCellInst3_LFInst_5_LFInst_2_n20 ,
         SubCellInst3_LFInst_5_LFInst_2_n19 ,
         SubCellInst3_LFInst_5_LFInst_2_n18 ,
         SubCellInst3_LFInst_5_LFInst_2_n17 ,
         SubCellInst3_LFInst_5_LFInst_2_n16 ,
         SubCellInst3_LFInst_5_LFInst_2_n15 ,
         SubCellInst3_LFInst_5_LFInst_3_n16 ,
         SubCellInst3_LFInst_5_LFInst_3_n15 ,
         SubCellInst3_LFInst_5_LFInst_3_n14 ,
         SubCellInst3_LFInst_5_LFInst_3_n13 ,
         SubCellInst3_LFInst_5_LFInst_3_n12 ,
         SubCellInst3_LFInst_5_LFInst_3_n11 ,
         SubCellInst3_LFInst_6_LFInst_0_n6 ,
         SubCellInst3_LFInst_6_LFInst_0_n5 ,
         SubCellInst3_LFInst_6_LFInst_0_n4 ,
         SubCellInst3_LFInst_6_LFInst_1_n18 ,
         SubCellInst3_LFInst_6_LFInst_1_n17 ,
         SubCellInst3_LFInst_6_LFInst_1_n16 ,
         SubCellInst3_LFInst_6_LFInst_1_n15 ,
         SubCellInst3_LFInst_6_LFInst_1_n14 ,
         SubCellInst3_LFInst_6_LFInst_1_n13 ,
         SubCellInst3_LFInst_6_LFInst_1_n12 ,
         SubCellInst3_LFInst_6_LFInst_1_n11 ,
         SubCellInst3_LFInst_6_LFInst_1_n10 ,
         SubCellInst3_LFInst_6_LFInst_2_n22 ,
         SubCellInst3_LFInst_6_LFInst_2_n21 ,
         SubCellInst3_LFInst_6_LFInst_2_n20 ,
         SubCellInst3_LFInst_6_LFInst_2_n19 ,
         SubCellInst3_LFInst_6_LFInst_2_n18 ,
         SubCellInst3_LFInst_6_LFInst_2_n17 ,
         SubCellInst3_LFInst_6_LFInst_2_n16 ,
         SubCellInst3_LFInst_6_LFInst_2_n15 ,
         SubCellInst3_LFInst_6_LFInst_3_n16 ,
         SubCellInst3_LFInst_6_LFInst_3_n15 ,
         SubCellInst3_LFInst_6_LFInst_3_n14 ,
         SubCellInst3_LFInst_6_LFInst_3_n13 ,
         SubCellInst3_LFInst_6_LFInst_3_n12 ,
         SubCellInst3_LFInst_6_LFInst_3_n11 ,
         SubCellInst3_LFInst_7_LFInst_0_n6 ,
         SubCellInst3_LFInst_7_LFInst_0_n5 ,
         SubCellInst3_LFInst_7_LFInst_0_n4 ,
         SubCellInst3_LFInst_7_LFInst_1_n18 ,
         SubCellInst3_LFInst_7_LFInst_1_n17 ,
         SubCellInst3_LFInst_7_LFInst_1_n16 ,
         SubCellInst3_LFInst_7_LFInst_1_n15 ,
         SubCellInst3_LFInst_7_LFInst_1_n14 ,
         SubCellInst3_LFInst_7_LFInst_1_n13 ,
         SubCellInst3_LFInst_7_LFInst_1_n12 ,
         SubCellInst3_LFInst_7_LFInst_1_n11 ,
         SubCellInst3_LFInst_7_LFInst_1_n10 ,
         SubCellInst3_LFInst_7_LFInst_2_n22 ,
         SubCellInst3_LFInst_7_LFInst_2_n21 ,
         SubCellInst3_LFInst_7_LFInst_2_n20 ,
         SubCellInst3_LFInst_7_LFInst_2_n19 ,
         SubCellInst3_LFInst_7_LFInst_2_n18 ,
         SubCellInst3_LFInst_7_LFInst_2_n17 ,
         SubCellInst3_LFInst_7_LFInst_2_n16 ,
         SubCellInst3_LFInst_7_LFInst_2_n15 ,
         SubCellInst3_LFInst_7_LFInst_3_n16 ,
         SubCellInst3_LFInst_7_LFInst_3_n15 ,
         SubCellInst3_LFInst_7_LFInst_3_n14 ,
         SubCellInst3_LFInst_7_LFInst_3_n13 ,
         SubCellInst3_LFInst_7_LFInst_3_n12 ,
         SubCellInst3_LFInst_7_LFInst_3_n11 ,
         SubCellInst3_LFInst_8_LFInst_0_n6 ,
         SubCellInst3_LFInst_8_LFInst_0_n5 ,
         SubCellInst3_LFInst_8_LFInst_0_n4 ,
         SubCellInst3_LFInst_8_LFInst_1_n18 ,
         SubCellInst3_LFInst_8_LFInst_1_n17 ,
         SubCellInst3_LFInst_8_LFInst_1_n16 ,
         SubCellInst3_LFInst_8_LFInst_1_n15 ,
         SubCellInst3_LFInst_8_LFInst_1_n14 ,
         SubCellInst3_LFInst_8_LFInst_1_n13 ,
         SubCellInst3_LFInst_8_LFInst_1_n12 ,
         SubCellInst3_LFInst_8_LFInst_1_n11 ,
         SubCellInst3_LFInst_8_LFInst_1_n10 ,
         SubCellInst3_LFInst_8_LFInst_2_n22 ,
         SubCellInst3_LFInst_8_LFInst_2_n21 ,
         SubCellInst3_LFInst_8_LFInst_2_n20 ,
         SubCellInst3_LFInst_8_LFInst_2_n19 ,
         SubCellInst3_LFInst_8_LFInst_2_n18 ,
         SubCellInst3_LFInst_8_LFInst_2_n17 ,
         SubCellInst3_LFInst_8_LFInst_2_n16 ,
         SubCellInst3_LFInst_8_LFInst_2_n15 ,
         SubCellInst3_LFInst_8_LFInst_3_n16 ,
         SubCellInst3_LFInst_8_LFInst_3_n15 ,
         SubCellInst3_LFInst_8_LFInst_3_n14 ,
         SubCellInst3_LFInst_8_LFInst_3_n13 ,
         SubCellInst3_LFInst_8_LFInst_3_n12 ,
         SubCellInst3_LFInst_8_LFInst_3_n11 ,
         SubCellInst3_LFInst_9_LFInst_0_n6 ,
         SubCellInst3_LFInst_9_LFInst_0_n5 ,
         SubCellInst3_LFInst_9_LFInst_0_n4 ,
         SubCellInst3_LFInst_9_LFInst_1_n18 ,
         SubCellInst3_LFInst_9_LFInst_1_n17 ,
         SubCellInst3_LFInst_9_LFInst_1_n16 ,
         SubCellInst3_LFInst_9_LFInst_1_n15 ,
         SubCellInst3_LFInst_9_LFInst_1_n14 ,
         SubCellInst3_LFInst_9_LFInst_1_n13 ,
         SubCellInst3_LFInst_9_LFInst_1_n12 ,
         SubCellInst3_LFInst_9_LFInst_1_n11 ,
         SubCellInst3_LFInst_9_LFInst_1_n10 ,
         SubCellInst3_LFInst_9_LFInst_2_n22 ,
         SubCellInst3_LFInst_9_LFInst_2_n21 ,
         SubCellInst3_LFInst_9_LFInst_2_n20 ,
         SubCellInst3_LFInst_9_LFInst_2_n19 ,
         SubCellInst3_LFInst_9_LFInst_2_n18 ,
         SubCellInst3_LFInst_9_LFInst_2_n17 ,
         SubCellInst3_LFInst_9_LFInst_2_n16 ,
         SubCellInst3_LFInst_9_LFInst_2_n15 ,
         SubCellInst3_LFInst_9_LFInst_3_n16 ,
         SubCellInst3_LFInst_9_LFInst_3_n15 ,
         SubCellInst3_LFInst_9_LFInst_3_n14 ,
         SubCellInst3_LFInst_9_LFInst_3_n13 ,
         SubCellInst3_LFInst_9_LFInst_3_n12 ,
         SubCellInst3_LFInst_9_LFInst_3_n11 ,
         SubCellInst3_LFInst_10_LFInst_0_n6 ,
         SubCellInst3_LFInst_10_LFInst_0_n5 ,
         SubCellInst3_LFInst_10_LFInst_0_n4 ,
         SubCellInst3_LFInst_10_LFInst_1_n18 ,
         SubCellInst3_LFInst_10_LFInst_1_n17 ,
         SubCellInst3_LFInst_10_LFInst_1_n16 ,
         SubCellInst3_LFInst_10_LFInst_1_n15 ,
         SubCellInst3_LFInst_10_LFInst_1_n14 ,
         SubCellInst3_LFInst_10_LFInst_1_n13 ,
         SubCellInst3_LFInst_10_LFInst_1_n12 ,
         SubCellInst3_LFInst_10_LFInst_1_n11 ,
         SubCellInst3_LFInst_10_LFInst_1_n10 ,
         SubCellInst3_LFInst_10_LFInst_2_n22 ,
         SubCellInst3_LFInst_10_LFInst_2_n21 ,
         SubCellInst3_LFInst_10_LFInst_2_n20 ,
         SubCellInst3_LFInst_10_LFInst_2_n19 ,
         SubCellInst3_LFInst_10_LFInst_2_n18 ,
         SubCellInst3_LFInst_10_LFInst_2_n17 ,
         SubCellInst3_LFInst_10_LFInst_2_n16 ,
         SubCellInst3_LFInst_10_LFInst_2_n15 ,
         SubCellInst3_LFInst_10_LFInst_3_n16 ,
         SubCellInst3_LFInst_10_LFInst_3_n15 ,
         SubCellInst3_LFInst_10_LFInst_3_n14 ,
         SubCellInst3_LFInst_10_LFInst_3_n13 ,
         SubCellInst3_LFInst_10_LFInst_3_n12 ,
         SubCellInst3_LFInst_10_LFInst_3_n11 ,
         SubCellInst3_LFInst_11_LFInst_0_n6 ,
         SubCellInst3_LFInst_11_LFInst_0_n5 ,
         SubCellInst3_LFInst_11_LFInst_0_n4 ,
         SubCellInst3_LFInst_11_LFInst_1_n18 ,
         SubCellInst3_LFInst_11_LFInst_1_n17 ,
         SubCellInst3_LFInst_11_LFInst_1_n16 ,
         SubCellInst3_LFInst_11_LFInst_1_n15 ,
         SubCellInst3_LFInst_11_LFInst_1_n14 ,
         SubCellInst3_LFInst_11_LFInst_1_n13 ,
         SubCellInst3_LFInst_11_LFInst_1_n12 ,
         SubCellInst3_LFInst_11_LFInst_1_n11 ,
         SubCellInst3_LFInst_11_LFInst_1_n10 ,
         SubCellInst3_LFInst_11_LFInst_2_n22 ,
         SubCellInst3_LFInst_11_LFInst_2_n21 ,
         SubCellInst3_LFInst_11_LFInst_2_n20 ,
         SubCellInst3_LFInst_11_LFInst_2_n19 ,
         SubCellInst3_LFInst_11_LFInst_2_n18 ,
         SubCellInst3_LFInst_11_LFInst_2_n17 ,
         SubCellInst3_LFInst_11_LFInst_2_n16 ,
         SubCellInst3_LFInst_11_LFInst_2_n15 ,
         SubCellInst3_LFInst_11_LFInst_3_n16 ,
         SubCellInst3_LFInst_11_LFInst_3_n15 ,
         SubCellInst3_LFInst_11_LFInst_3_n14 ,
         SubCellInst3_LFInst_11_LFInst_3_n13 ,
         SubCellInst3_LFInst_11_LFInst_3_n12 ,
         SubCellInst3_LFInst_11_LFInst_3_n11 ,
         SubCellInst3_LFInst_12_LFInst_0_n6 ,
         SubCellInst3_LFInst_12_LFInst_0_n5 ,
         SubCellInst3_LFInst_12_LFInst_0_n4 ,
         SubCellInst3_LFInst_12_LFInst_1_n18 ,
         SubCellInst3_LFInst_12_LFInst_1_n17 ,
         SubCellInst3_LFInst_12_LFInst_1_n16 ,
         SubCellInst3_LFInst_12_LFInst_1_n15 ,
         SubCellInst3_LFInst_12_LFInst_1_n14 ,
         SubCellInst3_LFInst_12_LFInst_1_n13 ,
         SubCellInst3_LFInst_12_LFInst_1_n12 ,
         SubCellInst3_LFInst_12_LFInst_1_n11 ,
         SubCellInst3_LFInst_12_LFInst_1_n10 ,
         SubCellInst3_LFInst_12_LFInst_2_n22 ,
         SubCellInst3_LFInst_12_LFInst_2_n21 ,
         SubCellInst3_LFInst_12_LFInst_2_n20 ,
         SubCellInst3_LFInst_12_LFInst_2_n19 ,
         SubCellInst3_LFInst_12_LFInst_2_n18 ,
         SubCellInst3_LFInst_12_LFInst_2_n17 ,
         SubCellInst3_LFInst_12_LFInst_2_n16 ,
         SubCellInst3_LFInst_12_LFInst_2_n15 ,
         SubCellInst3_LFInst_12_LFInst_3_n16 ,
         SubCellInst3_LFInst_12_LFInst_3_n15 ,
         SubCellInst3_LFInst_12_LFInst_3_n14 ,
         SubCellInst3_LFInst_12_LFInst_3_n13 ,
         SubCellInst3_LFInst_12_LFInst_3_n12 ,
         SubCellInst3_LFInst_12_LFInst_3_n11 ,
         SubCellInst3_LFInst_13_LFInst_0_n6 ,
         SubCellInst3_LFInst_13_LFInst_0_n5 ,
         SubCellInst3_LFInst_13_LFInst_0_n4 ,
         SubCellInst3_LFInst_13_LFInst_1_n18 ,
         SubCellInst3_LFInst_13_LFInst_1_n17 ,
         SubCellInst3_LFInst_13_LFInst_1_n16 ,
         SubCellInst3_LFInst_13_LFInst_1_n15 ,
         SubCellInst3_LFInst_13_LFInst_1_n14 ,
         SubCellInst3_LFInst_13_LFInst_1_n13 ,
         SubCellInst3_LFInst_13_LFInst_1_n12 ,
         SubCellInst3_LFInst_13_LFInst_1_n11 ,
         SubCellInst3_LFInst_13_LFInst_1_n10 ,
         SubCellInst3_LFInst_13_LFInst_2_n22 ,
         SubCellInst3_LFInst_13_LFInst_2_n21 ,
         SubCellInst3_LFInst_13_LFInst_2_n20 ,
         SubCellInst3_LFInst_13_LFInst_2_n19 ,
         SubCellInst3_LFInst_13_LFInst_2_n18 ,
         SubCellInst3_LFInst_13_LFInst_2_n17 ,
         SubCellInst3_LFInst_13_LFInst_2_n16 ,
         SubCellInst3_LFInst_13_LFInst_2_n15 ,
         SubCellInst3_LFInst_13_LFInst_3_n16 ,
         SubCellInst3_LFInst_13_LFInst_3_n15 ,
         SubCellInst3_LFInst_13_LFInst_3_n14 ,
         SubCellInst3_LFInst_13_LFInst_3_n13 ,
         SubCellInst3_LFInst_13_LFInst_3_n12 ,
         SubCellInst3_LFInst_13_LFInst_3_n11 ,
         SubCellInst3_LFInst_14_LFInst_0_n6 ,
         SubCellInst3_LFInst_14_LFInst_0_n5 ,
         SubCellInst3_LFInst_14_LFInst_0_n4 ,
         SubCellInst3_LFInst_14_LFInst_1_n18 ,
         SubCellInst3_LFInst_14_LFInst_1_n17 ,
         SubCellInst3_LFInst_14_LFInst_1_n16 ,
         SubCellInst3_LFInst_14_LFInst_1_n15 ,
         SubCellInst3_LFInst_14_LFInst_1_n14 ,
         SubCellInst3_LFInst_14_LFInst_1_n13 ,
         SubCellInst3_LFInst_14_LFInst_1_n12 ,
         SubCellInst3_LFInst_14_LFInst_1_n11 ,
         SubCellInst3_LFInst_14_LFInst_1_n10 ,
         SubCellInst3_LFInst_14_LFInst_2_n22 ,
         SubCellInst3_LFInst_14_LFInst_2_n21 ,
         SubCellInst3_LFInst_14_LFInst_2_n20 ,
         SubCellInst3_LFInst_14_LFInst_2_n19 ,
         SubCellInst3_LFInst_14_LFInst_2_n18 ,
         SubCellInst3_LFInst_14_LFInst_2_n17 ,
         SubCellInst3_LFInst_14_LFInst_2_n16 ,
         SubCellInst3_LFInst_14_LFInst_2_n15 ,
         SubCellInst3_LFInst_14_LFInst_3_n16 ,
         SubCellInst3_LFInst_14_LFInst_3_n15 ,
         SubCellInst3_LFInst_14_LFInst_3_n14 ,
         SubCellInst3_LFInst_14_LFInst_3_n13 ,
         SubCellInst3_LFInst_14_LFInst_3_n12 ,
         SubCellInst3_LFInst_14_LFInst_3_n11 ,
         SubCellInst3_LFInst_15_LFInst_0_n6 ,
         SubCellInst3_LFInst_15_LFInst_0_n5 ,
         SubCellInst3_LFInst_15_LFInst_0_n4 ,
         SubCellInst3_LFInst_15_LFInst_1_n18 ,
         SubCellInst3_LFInst_15_LFInst_1_n17 ,
         SubCellInst3_LFInst_15_LFInst_1_n16 ,
         SubCellInst3_LFInst_15_LFInst_1_n15 ,
         SubCellInst3_LFInst_15_LFInst_1_n14 ,
         SubCellInst3_LFInst_15_LFInst_1_n13 ,
         SubCellInst3_LFInst_15_LFInst_1_n12 ,
         SubCellInst3_LFInst_15_LFInst_1_n11 ,
         SubCellInst3_LFInst_15_LFInst_1_n10 ,
         SubCellInst3_LFInst_15_LFInst_2_n22 ,
         SubCellInst3_LFInst_15_LFInst_2_n21 ,
         SubCellInst3_LFInst_15_LFInst_2_n20 ,
         SubCellInst3_LFInst_15_LFInst_2_n19 ,
         SubCellInst3_LFInst_15_LFInst_2_n18 ,
         SubCellInst3_LFInst_15_LFInst_2_n17 ,
         SubCellInst3_LFInst_15_LFInst_2_n16 ,
         SubCellInst3_LFInst_15_LFInst_2_n15 ,
         SubCellInst3_LFInst_15_LFInst_3_n16 ,
         SubCellInst3_LFInst_15_LFInst_3_n15 ,
         SubCellInst3_LFInst_15_LFInst_3_n14 ,
         SubCellInst3_LFInst_15_LFInst_3_n13 ,
         SubCellInst3_LFInst_15_LFInst_3_n12 ,
         SubCellInst3_LFInst_15_LFInst_3_n11 , MCInst3_MC0_v0_2Inst_0_n2 ,
         MCInst3_MC0_v1_2Inst_0_n2 , MCInst3_MC0_v2_3Inst_0_n4 ,
         MCInst3_MC0_v2_3Inst_0_n3 , MCInst3_MC0_v3_3Inst_0_n2 ,
         MCInst3_MC0_v0_2Inst_1_n2 , MCInst3_MC0_v2_1Inst_1_n2 ,
         MCInst3_MC0_v2_2Inst_1_n4 , MCInst3_MC0_v2_2Inst_1_n3 ,
         MCInst3_MC0_v3_3Inst_1_n2 , MCInst3_MC0_v1_1Inst_2_n2 ,
         MCInst3_MC0_v1_2Inst_2_n2 , MCInst3_MC0_v2_1Inst_2_n2 ,
         MCInst3_MC0_v2_2Inst_2_n2 , MCInst3_MC0_v3_1Inst_2_n2 ,
         MCInst3_MC0_v1_2Inst_3_n4 , MCInst3_MC0_v1_2Inst_3_n3 ,
         MCInst3_MC0_v2_2Inst_3_n2 , MCInst3_MC0_v2_3Inst_3_n2 ,
         MCInst3_MC0_r0Inst_XORInst_0_0_n5 ,
         MCInst3_MC0_r0Inst_XORInst_0_0_n4 ,
         MCInst3_MC0_r0Inst_XORInst_0_1_n5 ,
         MCInst3_MC0_r0Inst_XORInst_0_1_n4 ,
         MCInst3_MC0_r0Inst_XORInst_0_2_n5 ,
         MCInst3_MC0_r0Inst_XORInst_0_2_n4 ,
         MCInst3_MC0_r0Inst_XORInst_0_3_n5 ,
         MCInst3_MC0_r0Inst_XORInst_0_3_n4 ,
         MCInst3_MC0_r1Inst_XORInst_0_0_n5 ,
         MCInst3_MC0_r1Inst_XORInst_0_0_n4 ,
         MCInst3_MC0_r1Inst_XORInst_0_1_n5 ,
         MCInst3_MC0_r1Inst_XORInst_0_1_n4 ,
         MCInst3_MC0_r1Inst_XORInst_0_2_n5 ,
         MCInst3_MC0_r1Inst_XORInst_0_2_n4 ,
         MCInst3_MC0_r1Inst_XORInst_0_3_n5 ,
         MCInst3_MC0_r1Inst_XORInst_0_3_n4 ,
         MCInst3_MC0_r2Inst_XORInst_0_0_n5 ,
         MCInst3_MC0_r2Inst_XORInst_0_0_n4 ,
         MCInst3_MC0_r2Inst_XORInst_0_1_n5 ,
         MCInst3_MC0_r2Inst_XORInst_0_1_n4 ,
         MCInst3_MC0_r2Inst_XORInst_0_2_n5 ,
         MCInst3_MC0_r2Inst_XORInst_0_2_n4 ,
         MCInst3_MC0_r2Inst_XORInst_0_3_n5 ,
         MCInst3_MC0_r2Inst_XORInst_0_3_n4 ,
         MCInst3_MC0_r3Inst_XORInst_0_0_n5 ,
         MCInst3_MC0_r3Inst_XORInst_0_0_n4 ,
         MCInst3_MC0_r3Inst_XORInst_0_1_n5 ,
         MCInst3_MC0_r3Inst_XORInst_0_1_n4 ,
         MCInst3_MC0_r3Inst_XORInst_0_2_n5 ,
         MCInst3_MC0_r3Inst_XORInst_0_2_n4 ,
         MCInst3_MC0_r3Inst_XORInst_0_3_n5 ,
         MCInst3_MC0_r3Inst_XORInst_0_3_n4 , MCInst3_MC1_v0_2Inst_0_n2 ,
         MCInst3_MC1_v1_2Inst_0_n2 , MCInst3_MC1_v2_3Inst_0_n4 ,
         MCInst3_MC1_v2_3Inst_0_n3 , MCInst3_MC1_v3_3Inst_0_n2 ,
         MCInst3_MC1_v0_2Inst_1_n2 , MCInst3_MC1_v2_1Inst_1_n2 ,
         MCInst3_MC1_v2_2Inst_1_n4 , MCInst3_MC1_v2_2Inst_1_n3 ,
         MCInst3_MC1_v3_3Inst_1_n2 , MCInst3_MC1_v1_1Inst_2_n2 ,
         MCInst3_MC1_v1_2Inst_2_n2 , MCInst3_MC1_v2_1Inst_2_n2 ,
         MCInst3_MC1_v2_2Inst_2_n2 , MCInst3_MC1_v3_1Inst_2_n2 ,
         MCInst3_MC1_v1_2Inst_3_n4 , MCInst3_MC1_v1_2Inst_3_n3 ,
         MCInst3_MC1_v2_2Inst_3_n2 , MCInst3_MC1_v2_3Inst_3_n2 ,
         MCInst3_MC1_r0Inst_XORInst_0_0_n5 ,
         MCInst3_MC1_r0Inst_XORInst_0_0_n4 ,
         MCInst3_MC1_r0Inst_XORInst_0_1_n5 ,
         MCInst3_MC1_r0Inst_XORInst_0_1_n4 ,
         MCInst3_MC1_r0Inst_XORInst_0_2_n5 ,
         MCInst3_MC1_r0Inst_XORInst_0_2_n4 ,
         MCInst3_MC1_r0Inst_XORInst_0_3_n5 ,
         MCInst3_MC1_r0Inst_XORInst_0_3_n4 ,
         MCInst3_MC1_r1Inst_XORInst_0_0_n5 ,
         MCInst3_MC1_r1Inst_XORInst_0_0_n4 ,
         MCInst3_MC1_r1Inst_XORInst_0_1_n5 ,
         MCInst3_MC1_r1Inst_XORInst_0_1_n4 ,
         MCInst3_MC1_r1Inst_XORInst_0_2_n5 ,
         MCInst3_MC1_r1Inst_XORInst_0_2_n4 ,
         MCInst3_MC1_r1Inst_XORInst_0_3_n5 ,
         MCInst3_MC1_r1Inst_XORInst_0_3_n4 ,
         MCInst3_MC1_r2Inst_XORInst_0_0_n5 ,
         MCInst3_MC1_r2Inst_XORInst_0_0_n4 ,
         MCInst3_MC1_r2Inst_XORInst_0_1_n5 ,
         MCInst3_MC1_r2Inst_XORInst_0_1_n4 ,
         MCInst3_MC1_r2Inst_XORInst_0_2_n5 ,
         MCInst3_MC1_r2Inst_XORInst_0_2_n4 ,
         MCInst3_MC1_r2Inst_XORInst_0_3_n5 ,
         MCInst3_MC1_r2Inst_XORInst_0_3_n4 ,
         MCInst3_MC1_r3Inst_XORInst_0_0_n5 ,
         MCInst3_MC1_r3Inst_XORInst_0_0_n4 ,
         MCInst3_MC1_r3Inst_XORInst_0_1_n5 ,
         MCInst3_MC1_r3Inst_XORInst_0_1_n4 ,
         MCInst3_MC1_r3Inst_XORInst_0_2_n5 ,
         MCInst3_MC1_r3Inst_XORInst_0_2_n4 ,
         MCInst3_MC1_r3Inst_XORInst_0_3_n5 ,
         MCInst3_MC1_r3Inst_XORInst_0_3_n4 , MCInst3_MC2_v0_2Inst_0_n2 ,
         MCInst3_MC2_v1_2Inst_0_n2 , MCInst3_MC2_v2_3Inst_0_n4 ,
         MCInst3_MC2_v2_3Inst_0_n3 , MCInst3_MC2_v3_3Inst_0_n2 ,
         MCInst3_MC2_v0_2Inst_1_n2 , MCInst3_MC2_v2_1Inst_1_n2 ,
         MCInst3_MC2_v2_2Inst_1_n4 , MCInst3_MC2_v2_2Inst_1_n3 ,
         MCInst3_MC2_v3_3Inst_1_n2 , MCInst3_MC2_v1_1Inst_2_n2 ,
         MCInst3_MC2_v1_2Inst_2_n2 , MCInst3_MC2_v2_1Inst_2_n2 ,
         MCInst3_MC2_v2_2Inst_2_n2 , MCInst3_MC2_v3_1Inst_2_n2 ,
         MCInst3_MC2_v1_2Inst_3_n4 , MCInst3_MC2_v1_2Inst_3_n3 ,
         MCInst3_MC2_v2_2Inst_3_n2 , MCInst3_MC2_v2_3Inst_3_n2 ,
         MCInst3_MC2_r0Inst_XORInst_0_0_n5 ,
         MCInst3_MC2_r0Inst_XORInst_0_0_n4 ,
         MCInst3_MC2_r0Inst_XORInst_0_1_n5 ,
         MCInst3_MC2_r0Inst_XORInst_0_1_n4 ,
         MCInst3_MC2_r0Inst_XORInst_0_2_n5 ,
         MCInst3_MC2_r0Inst_XORInst_0_2_n4 ,
         MCInst3_MC2_r0Inst_XORInst_0_3_n5 ,
         MCInst3_MC2_r0Inst_XORInst_0_3_n4 ,
         MCInst3_MC2_r1Inst_XORInst_0_0_n5 ,
         MCInst3_MC2_r1Inst_XORInst_0_0_n4 ,
         MCInst3_MC2_r1Inst_XORInst_0_1_n5 ,
         MCInst3_MC2_r1Inst_XORInst_0_1_n4 ,
         MCInst3_MC2_r1Inst_XORInst_0_2_n5 ,
         MCInst3_MC2_r1Inst_XORInst_0_2_n4 ,
         MCInst3_MC2_r1Inst_XORInst_0_3_n5 ,
         MCInst3_MC2_r1Inst_XORInst_0_3_n4 ,
         MCInst3_MC2_r2Inst_XORInst_0_0_n5 ,
         MCInst3_MC2_r2Inst_XORInst_0_0_n4 ,
         MCInst3_MC2_r2Inst_XORInst_0_1_n5 ,
         MCInst3_MC2_r2Inst_XORInst_0_1_n4 ,
         MCInst3_MC2_r2Inst_XORInst_0_2_n5 ,
         MCInst3_MC2_r2Inst_XORInst_0_2_n4 ,
         MCInst3_MC2_r2Inst_XORInst_0_3_n5 ,
         MCInst3_MC2_r2Inst_XORInst_0_3_n4 ,
         MCInst3_MC2_r3Inst_XORInst_0_0_n5 ,
         MCInst3_MC2_r3Inst_XORInst_0_0_n4 ,
         MCInst3_MC2_r3Inst_XORInst_0_1_n5 ,
         MCInst3_MC2_r3Inst_XORInst_0_1_n4 ,
         MCInst3_MC2_r3Inst_XORInst_0_2_n5 ,
         MCInst3_MC2_r3Inst_XORInst_0_2_n4 ,
         MCInst3_MC2_r3Inst_XORInst_0_3_n5 ,
         MCInst3_MC2_r3Inst_XORInst_0_3_n4 , MCInst3_MC3_v0_2Inst_0_n2 ,
         MCInst3_MC3_v1_2Inst_0_n2 , MCInst3_MC3_v2_3Inst_0_n4 ,
         MCInst3_MC3_v2_3Inst_0_n3 , MCInst3_MC3_v3_3Inst_0_n2 ,
         MCInst3_MC3_v0_2Inst_1_n2 , MCInst3_MC3_v2_1Inst_1_n2 ,
         MCInst3_MC3_v2_2Inst_1_n4 , MCInst3_MC3_v2_2Inst_1_n3 ,
         MCInst3_MC3_v3_3Inst_1_n2 , MCInst3_MC3_v1_1Inst_2_n2 ,
         MCInst3_MC3_v1_2Inst_2_n2 , MCInst3_MC3_v2_1Inst_2_n2 ,
         MCInst3_MC3_v2_2Inst_2_n2 , MCInst3_MC3_v3_1Inst_2_n2 ,
         MCInst3_MC3_v1_2Inst_3_n4 , MCInst3_MC3_v1_2Inst_3_n3 ,
         MCInst3_MC3_v2_2Inst_3_n2 , MCInst3_MC3_v2_3Inst_3_n2 ,
         MCInst3_MC3_r0Inst_XORInst_0_0_n5 ,
         MCInst3_MC3_r0Inst_XORInst_0_0_n4 ,
         MCInst3_MC3_r0Inst_XORInst_0_1_n5 ,
         MCInst3_MC3_r0Inst_XORInst_0_1_n4 ,
         MCInst3_MC3_r0Inst_XORInst_0_2_n5 ,
         MCInst3_MC3_r0Inst_XORInst_0_2_n4 ,
         MCInst3_MC3_r0Inst_XORInst_0_3_n5 ,
         MCInst3_MC3_r0Inst_XORInst_0_3_n4 ,
         MCInst3_MC3_r1Inst_XORInst_0_0_n5 ,
         MCInst3_MC3_r1Inst_XORInst_0_0_n4 ,
         MCInst3_MC3_r1Inst_XORInst_0_1_n5 ,
         MCInst3_MC3_r1Inst_XORInst_0_1_n4 ,
         MCInst3_MC3_r1Inst_XORInst_0_2_n5 ,
         MCInst3_MC3_r1Inst_XORInst_0_2_n4 ,
         MCInst3_MC3_r1Inst_XORInst_0_3_n5 ,
         MCInst3_MC3_r1Inst_XORInst_0_3_n4 ,
         MCInst3_MC3_r2Inst_XORInst_0_0_n5 ,
         MCInst3_MC3_r2Inst_XORInst_0_0_n4 ,
         MCInst3_MC3_r2Inst_XORInst_0_1_n5 ,
         MCInst3_MC3_r2Inst_XORInst_0_1_n4 ,
         MCInst3_MC3_r2Inst_XORInst_0_2_n5 ,
         MCInst3_MC3_r2Inst_XORInst_0_2_n4 ,
         MCInst3_MC3_r2Inst_XORInst_0_3_n5 ,
         MCInst3_MC3_r2Inst_XORInst_0_3_n4 ,
         MCInst3_MC3_r3Inst_XORInst_0_0_n5 ,
         MCInst3_MC3_r3Inst_XORInst_0_0_n4 ,
         MCInst3_MC3_r3Inst_XORInst_0_1_n5 ,
         MCInst3_MC3_r3Inst_XORInst_0_1_n4 ,
         MCInst3_MC3_r3Inst_XORInst_0_2_n5 ,
         MCInst3_MC3_r3Inst_XORInst_0_2_n4 ,
         MCInst3_MC3_r3Inst_XORInst_0_3_n5 ,
         MCInst3_MC3_r3Inst_XORInst_0_3_n4 ,
         Red_PlaintextInst_LFInst_0_LFInst_0_n4 ,
         Red_PlaintextInst_LFInst_0_LFInst_0_n3 ,
         Red_PlaintextInst_LFInst_1_LFInst_0_n4 ,
         Red_PlaintextInst_LFInst_1_LFInst_0_n3 ,
         Red_PlaintextInst_LFInst_2_LFInst_0_n4 ,
         Red_PlaintextInst_LFInst_2_LFInst_0_n3 ,
         Red_PlaintextInst_LFInst_3_LFInst_0_n4 ,
         Red_PlaintextInst_LFInst_3_LFInst_0_n3 ,
         Red_PlaintextInst_LFInst_4_LFInst_0_n4 ,
         Red_PlaintextInst_LFInst_4_LFInst_0_n3 ,
         Red_PlaintextInst_LFInst_5_LFInst_0_n4 ,
         Red_PlaintextInst_LFInst_5_LFInst_0_n3 ,
         Red_PlaintextInst_LFInst_6_LFInst_0_n4 ,
         Red_PlaintextInst_LFInst_6_LFInst_0_n3 ,
         Red_PlaintextInst_LFInst_7_LFInst_0_n4 ,
         Red_PlaintextInst_LFInst_7_LFInst_0_n3 ,
         Red_PlaintextInst_LFInst_8_LFInst_0_n4 ,
         Red_PlaintextInst_LFInst_8_LFInst_0_n3 ,
         Red_PlaintextInst_LFInst_9_LFInst_0_n4 ,
         Red_PlaintextInst_LFInst_9_LFInst_0_n3 ,
         Red_PlaintextInst_LFInst_10_LFInst_0_n4 ,
         Red_PlaintextInst_LFInst_10_LFInst_0_n3 ,
         Red_PlaintextInst_LFInst_11_LFInst_0_n4 ,
         Red_PlaintextInst_LFInst_11_LFInst_0_n3 ,
         Red_PlaintextInst_LFInst_12_LFInst_0_n4 ,
         Red_PlaintextInst_LFInst_12_LFInst_0_n3 ,
         Red_PlaintextInst_LFInst_13_LFInst_0_n4 ,
         Red_PlaintextInst_LFInst_13_LFInst_0_n3 ,
         Red_PlaintextInst_LFInst_14_LFInst_0_n4 ,
         Red_PlaintextInst_LFInst_14_LFInst_0_n3 ,
         Red_PlaintextInst_LFInst_15_LFInst_0_n4 ,
         Red_PlaintextInst_LFInst_15_LFInst_0_n3 ,
         Red_SubCellInst_LFInst_0_LFInst_0_n6 ,
         Red_SubCellInst_LFInst_0_LFInst_0_n5 ,
         Red_SubCellInst_LFInst_0_LFInst_0_n4 ,
         Red_SubCellInst_LFInst_1_LFInst_0_n6 ,
         Red_SubCellInst_LFInst_1_LFInst_0_n5 ,
         Red_SubCellInst_LFInst_1_LFInst_0_n4 ,
         Red_SubCellInst_LFInst_2_LFInst_0_n6 ,
         Red_SubCellInst_LFInst_2_LFInst_0_n5 ,
         Red_SubCellInst_LFInst_2_LFInst_0_n4 ,
         Red_SubCellInst_LFInst_3_LFInst_0_n6 ,
         Red_SubCellInst_LFInst_3_LFInst_0_n5 ,
         Red_SubCellInst_LFInst_3_LFInst_0_n4 ,
         Red_SubCellInst_LFInst_4_LFInst_0_n6 ,
         Red_SubCellInst_LFInst_4_LFInst_0_n5 ,
         Red_SubCellInst_LFInst_4_LFInst_0_n4 ,
         Red_SubCellInst_LFInst_5_LFInst_0_n6 ,
         Red_SubCellInst_LFInst_5_LFInst_0_n5 ,
         Red_SubCellInst_LFInst_5_LFInst_0_n4 ,
         Red_SubCellInst_LFInst_6_LFInst_0_n6 ,
         Red_SubCellInst_LFInst_6_LFInst_0_n5 ,
         Red_SubCellInst_LFInst_6_LFInst_0_n4 ,
         Red_SubCellInst_LFInst_7_LFInst_0_n6 ,
         Red_SubCellInst_LFInst_7_LFInst_0_n5 ,
         Red_SubCellInst_LFInst_7_LFInst_0_n4 ,
         Red_SubCellInst_LFInst_8_LFInst_0_n6 ,
         Red_SubCellInst_LFInst_8_LFInst_0_n5 ,
         Red_SubCellInst_LFInst_8_LFInst_0_n4 ,
         Red_SubCellInst_LFInst_9_LFInst_0_n6 ,
         Red_SubCellInst_LFInst_9_LFInst_0_n5 ,
         Red_SubCellInst_LFInst_9_LFInst_0_n4 ,
         Red_SubCellInst_LFInst_10_LFInst_0_n6 ,
         Red_SubCellInst_LFInst_10_LFInst_0_n5 ,
         Red_SubCellInst_LFInst_10_LFInst_0_n4 ,
         Red_SubCellInst_LFInst_11_LFInst_0_n6 ,
         Red_SubCellInst_LFInst_11_LFInst_0_n5 ,
         Red_SubCellInst_LFInst_11_LFInst_0_n4 ,
         Red_SubCellInst_LFInst_12_LFInst_0_n6 ,
         Red_SubCellInst_LFInst_12_LFInst_0_n5 ,
         Red_SubCellInst_LFInst_12_LFInst_0_n4 ,
         Red_SubCellInst_LFInst_13_LFInst_0_n6 ,
         Red_SubCellInst_LFInst_13_LFInst_0_n5 ,
         Red_SubCellInst_LFInst_13_LFInst_0_n4 ,
         Red_SubCellInst_LFInst_14_LFInst_0_n6 ,
         Red_SubCellInst_LFInst_14_LFInst_0_n5 ,
         Red_SubCellInst_LFInst_14_LFInst_0_n4 ,
         Red_SubCellInst_LFInst_15_LFInst_0_n6 ,
         Red_SubCellInst_LFInst_15_LFInst_0_n5 ,
         Red_SubCellInst_LFInst_15_LFInst_0_n4 , Red_MCInst_MC0_v3_3[0] ,
         Red_MCInst_MC0_v3_2[0] , Red_MCInst_MC0_v3_1[0] ,
         Red_MCInst_MC0_v3_0[0] , Red_MCInst_MC0_v2_3[0] ,
         Red_MCInst_MC0_v2_2[0] , Red_MCInst_MC0_v2_1[0] ,
         Red_MCInst_MC0_v2_0[0] , Red_MCInst_MC0_v1_3[0] ,
         Red_MCInst_MC0_v1_2[0] , Red_MCInst_MC0_v1_1[0] ,
         Red_MCInst_MC0_v1_0[0] , Red_MCInst_MC0_v0_3[0] ,
         Red_MCInst_MC0_v0_2[0] , Red_MCInst_MC0_v0_1[0] ,
         Red_MCInst_MC0_v0_0[0] , Red_MCInst_MC0_v0_3Inst_0_n2 ,
         Red_MCInst_MC0_v1_0Inst_0_n4 , Red_MCInst_MC0_v1_0Inst_0_n3 ,
         Red_MCInst_MC0_v1_3Inst_0_n2 , Red_MCInst_MC0_v2_0Inst_0_n2 ,
         Red_MCInst_MC0_v3_0Inst_0_n2 , Red_MCInst_MC0_v3_2Inst_0_n2 ,
         Red_MCInst_MC0_r0Inst_XORInst_0_0_n5 ,
         Red_MCInst_MC0_r0Inst_XORInst_0_0_n4 ,
         Red_MCInst_MC0_r1Inst_XORInst_0_0_n5 ,
         Red_MCInst_MC0_r1Inst_XORInst_0_0_n4 ,
         Red_MCInst_MC0_r2Inst_XORInst_0_0_n5 ,
         Red_MCInst_MC0_r2Inst_XORInst_0_0_n4 ,
         Red_MCInst_MC0_r3Inst_XORInst_0_0_n5 ,
         Red_MCInst_MC0_r3Inst_XORInst_0_0_n4 , Red_MCInst_MC1_v3_3[0] ,
         Red_MCInst_MC1_v3_2[0] , Red_MCInst_MC1_v3_1[0] ,
         Red_MCInst_MC1_v3_0[0] , Red_MCInst_MC1_v2_3[0] ,
         Red_MCInst_MC1_v2_2[0] , Red_MCInst_MC1_v2_1[0] ,
         Red_MCInst_MC1_v2_0[0] , Red_MCInst_MC1_v1_3[0] ,
         Red_MCInst_MC1_v1_2[0] , Red_MCInst_MC1_v1_1[0] ,
         Red_MCInst_MC1_v1_0[0] , Red_MCInst_MC1_v0_3[0] ,
         Red_MCInst_MC1_v0_2[0] , Red_MCInst_MC1_v0_1[0] ,
         Red_MCInst_MC1_v0_0[0] , Red_MCInst_MC1_v0_3Inst_0_n2 ,
         Red_MCInst_MC1_v1_0Inst_0_n4 , Red_MCInst_MC1_v1_0Inst_0_n3 ,
         Red_MCInst_MC1_v1_3Inst_0_n2 , Red_MCInst_MC1_v2_0Inst_0_n2 ,
         Red_MCInst_MC1_v3_0Inst_0_n2 , Red_MCInst_MC1_v3_2Inst_0_n2 ,
         Red_MCInst_MC1_r0Inst_XORInst_0_0_n5 ,
         Red_MCInst_MC1_r0Inst_XORInst_0_0_n4 ,
         Red_MCInst_MC1_r1Inst_XORInst_0_0_n5 ,
         Red_MCInst_MC1_r1Inst_XORInst_0_0_n4 ,
         Red_MCInst_MC1_r2Inst_XORInst_0_0_n5 ,
         Red_MCInst_MC1_r2Inst_XORInst_0_0_n4 ,
         Red_MCInst_MC1_r3Inst_XORInst_0_0_n5 ,
         Red_MCInst_MC1_r3Inst_XORInst_0_0_n4 , Red_MCInst_MC2_v3_3[0] ,
         Red_MCInst_MC2_v3_2[0] , Red_MCInst_MC2_v3_1[0] ,
         Red_MCInst_MC2_v3_0[0] , Red_MCInst_MC2_v2_3[0] ,
         Red_MCInst_MC2_v2_2[0] , Red_MCInst_MC2_v2_1[0] ,
         Red_MCInst_MC2_v2_0[0] , Red_MCInst_MC2_v1_3[0] ,
         Red_MCInst_MC2_v1_2[0] , Red_MCInst_MC2_v1_1[0] ,
         Red_MCInst_MC2_v1_0[0] , Red_MCInst_MC2_v0_3[0] ,
         Red_MCInst_MC2_v0_2[0] , Red_MCInst_MC2_v0_1[0] ,
         Red_MCInst_MC2_v0_0[0] , Red_MCInst_MC2_v0_3Inst_0_n2 ,
         Red_MCInst_MC2_v1_0Inst_0_n4 , Red_MCInst_MC2_v1_0Inst_0_n3 ,
         Red_MCInst_MC2_v1_3Inst_0_n2 , Red_MCInst_MC2_v2_0Inst_0_n2 ,
         Red_MCInst_MC2_v3_0Inst_0_n2 , Red_MCInst_MC2_v3_2Inst_0_n2 ,
         Red_MCInst_MC2_r0Inst_XORInst_0_0_n5 ,
         Red_MCInst_MC2_r0Inst_XORInst_0_0_n4 ,
         Red_MCInst_MC2_r1Inst_XORInst_0_0_n5 ,
         Red_MCInst_MC2_r1Inst_XORInst_0_0_n4 ,
         Red_MCInst_MC2_r2Inst_XORInst_0_0_n5 ,
         Red_MCInst_MC2_r2Inst_XORInst_0_0_n4 ,
         Red_MCInst_MC2_r3Inst_XORInst_0_0_n5 ,
         Red_MCInst_MC2_r3Inst_XORInst_0_0_n4 , Red_MCInst_MC3_v3_3[0] ,
         Red_MCInst_MC3_v3_2[0] , Red_MCInst_MC3_v3_1[0] ,
         Red_MCInst_MC3_v3_0[0] , Red_MCInst_MC3_v2_3[0] ,
         Red_MCInst_MC3_v2_2[0] , Red_MCInst_MC3_v2_1[0] ,
         Red_MCInst_MC3_v2_0[0] , Red_MCInst_MC3_v1_3[0] ,
         Red_MCInst_MC3_v1_2[0] , Red_MCInst_MC3_v1_1[0] ,
         Red_MCInst_MC3_v1_0[0] , Red_MCInst_MC3_v0_3[0] ,
         Red_MCInst_MC3_v0_2[0] , Red_MCInst_MC3_v0_1[0] ,
         Red_MCInst_MC3_v0_0[0] , Red_MCInst_MC3_v0_3Inst_0_n2 ,
         Red_MCInst_MC3_v1_0Inst_0_n4 , Red_MCInst_MC3_v1_0Inst_0_n3 ,
         Red_MCInst_MC3_v1_3Inst_0_n2 , Red_MCInst_MC3_v2_0Inst_0_n2 ,
         Red_MCInst_MC3_v3_0Inst_0_n2 , Red_MCInst_MC3_v3_2Inst_0_n2 ,
         Red_MCInst_MC3_r0Inst_XORInst_0_0_n5 ,
         Red_MCInst_MC3_r0Inst_XORInst_0_0_n4 ,
         Red_MCInst_MC3_r1Inst_XORInst_0_0_n5 ,
         Red_MCInst_MC3_r1Inst_XORInst_0_0_n4 ,
         Red_MCInst_MC3_r2Inst_XORInst_0_0_n5 ,
         Red_MCInst_MC3_r2Inst_XORInst_0_0_n4 ,
         Red_MCInst_MC3_r3Inst_XORInst_0_0_n5 ,
         Red_MCInst_MC3_r3Inst_XORInst_0_0_n4 ,
         Red_SubCellInst2_LFInst_0_LFInst_0_n6 ,
         Red_SubCellInst2_LFInst_0_LFInst_0_n5 ,
         Red_SubCellInst2_LFInst_0_LFInst_0_n4 ,
         Red_SubCellInst2_LFInst_1_LFInst_0_n6 ,
         Red_SubCellInst2_LFInst_1_LFInst_0_n5 ,
         Red_SubCellInst2_LFInst_1_LFInst_0_n4 ,
         Red_SubCellInst2_LFInst_2_LFInst_0_n6 ,
         Red_SubCellInst2_LFInst_2_LFInst_0_n5 ,
         Red_SubCellInst2_LFInst_2_LFInst_0_n4 ,
         Red_SubCellInst2_LFInst_3_LFInst_0_n6 ,
         Red_SubCellInst2_LFInst_3_LFInst_0_n5 ,
         Red_SubCellInst2_LFInst_3_LFInst_0_n4 ,
         Red_SubCellInst2_LFInst_4_LFInst_0_n6 ,
         Red_SubCellInst2_LFInst_4_LFInst_0_n5 ,
         Red_SubCellInst2_LFInst_4_LFInst_0_n4 ,
         Red_SubCellInst2_LFInst_5_LFInst_0_n6 ,
         Red_SubCellInst2_LFInst_5_LFInst_0_n5 ,
         Red_SubCellInst2_LFInst_5_LFInst_0_n4 ,
         Red_SubCellInst2_LFInst_6_LFInst_0_n6 ,
         Red_SubCellInst2_LFInst_6_LFInst_0_n5 ,
         Red_SubCellInst2_LFInst_6_LFInst_0_n4 ,
         Red_SubCellInst2_LFInst_7_LFInst_0_n6 ,
         Red_SubCellInst2_LFInst_7_LFInst_0_n5 ,
         Red_SubCellInst2_LFInst_7_LFInst_0_n4 ,
         Red_SubCellInst2_LFInst_8_LFInst_0_n6 ,
         Red_SubCellInst2_LFInst_8_LFInst_0_n5 ,
         Red_SubCellInst2_LFInst_8_LFInst_0_n4 ,
         Red_SubCellInst2_LFInst_9_LFInst_0_n6 ,
         Red_SubCellInst2_LFInst_9_LFInst_0_n5 ,
         Red_SubCellInst2_LFInst_9_LFInst_0_n4 ,
         Red_SubCellInst2_LFInst_10_LFInst_0_n6 ,
         Red_SubCellInst2_LFInst_10_LFInst_0_n5 ,
         Red_SubCellInst2_LFInst_10_LFInst_0_n4 ,
         Red_SubCellInst2_LFInst_11_LFInst_0_n6 ,
         Red_SubCellInst2_LFInst_11_LFInst_0_n5 ,
         Red_SubCellInst2_LFInst_11_LFInst_0_n4 ,
         Red_SubCellInst2_LFInst_12_LFInst_0_n6 ,
         Red_SubCellInst2_LFInst_12_LFInst_0_n5 ,
         Red_SubCellInst2_LFInst_12_LFInst_0_n4 ,
         Red_SubCellInst2_LFInst_13_LFInst_0_n6 ,
         Red_SubCellInst2_LFInst_13_LFInst_0_n5 ,
         Red_SubCellInst2_LFInst_13_LFInst_0_n4 ,
         Red_SubCellInst2_LFInst_14_LFInst_0_n6 ,
         Red_SubCellInst2_LFInst_14_LFInst_0_n5 ,
         Red_SubCellInst2_LFInst_14_LFInst_0_n4 ,
         Red_SubCellInst2_LFInst_15_LFInst_0_n6 ,
         Red_SubCellInst2_LFInst_15_LFInst_0_n5 ,
         Red_SubCellInst2_LFInst_15_LFInst_0_n4 , Red_MCInst2_MC0_v3_3[0] ,
         Red_MCInst2_MC0_v3_2[0] , Red_MCInst2_MC0_v3_1[0] ,
         Red_MCInst2_MC0_v3_0[0] , Red_MCInst2_MC0_v2_3[0] ,
         Red_MCInst2_MC0_v2_2[0] , Red_MCInst2_MC0_v2_1[0] ,
         Red_MCInst2_MC0_v2_0[0] , Red_MCInst2_MC0_v1_3[0] ,
         Red_MCInst2_MC0_v1_2[0] , Red_MCInst2_MC0_v1_1[0] ,
         Red_MCInst2_MC0_v1_0[0] , Red_MCInst2_MC0_v0_3[0] ,
         Red_MCInst2_MC0_v0_2[0] , Red_MCInst2_MC0_v0_1[0] ,
         Red_MCInst2_MC0_v0_0[0] , Red_MCInst2_MC0_v0_3Inst_0_n2 ,
         Red_MCInst2_MC0_v1_0Inst_0_n4 , Red_MCInst2_MC0_v1_0Inst_0_n3 ,
         Red_MCInst2_MC0_v1_3Inst_0_n2 , Red_MCInst2_MC0_v2_0Inst_0_n2 ,
         Red_MCInst2_MC0_v3_0Inst_0_n2 , Red_MCInst2_MC0_v3_2Inst_0_n2 ,
         Red_MCInst2_MC0_r0Inst_XORInst_0_0_n5 ,
         Red_MCInst2_MC0_r0Inst_XORInst_0_0_n4 ,
         Red_MCInst2_MC0_r1Inst_XORInst_0_0_n5 ,
         Red_MCInst2_MC0_r1Inst_XORInst_0_0_n4 ,
         Red_MCInst2_MC0_r2Inst_XORInst_0_0_n5 ,
         Red_MCInst2_MC0_r2Inst_XORInst_0_0_n4 ,
         Red_MCInst2_MC0_r3Inst_XORInst_0_0_n5 ,
         Red_MCInst2_MC0_r3Inst_XORInst_0_0_n4 , Red_MCInst2_MC1_v3_3[0] ,
         Red_MCInst2_MC1_v3_2[0] , Red_MCInst2_MC1_v3_1[0] ,
         Red_MCInst2_MC1_v3_0[0] , Red_MCInst2_MC1_v2_3[0] ,
         Red_MCInst2_MC1_v2_2[0] , Red_MCInst2_MC1_v2_1[0] ,
         Red_MCInst2_MC1_v2_0[0] , Red_MCInst2_MC1_v1_3[0] ,
         Red_MCInst2_MC1_v1_2[0] , Red_MCInst2_MC1_v1_1[0] ,
         Red_MCInst2_MC1_v1_0[0] , Red_MCInst2_MC1_v0_3[0] ,
         Red_MCInst2_MC1_v0_2[0] , Red_MCInst2_MC1_v0_1[0] ,
         Red_MCInst2_MC1_v0_0[0] , Red_MCInst2_MC1_v0_3Inst_0_n2 ,
         Red_MCInst2_MC1_v1_0Inst_0_n4 , Red_MCInst2_MC1_v1_0Inst_0_n3 ,
         Red_MCInst2_MC1_v1_3Inst_0_n2 , Red_MCInst2_MC1_v2_0Inst_0_n2 ,
         Red_MCInst2_MC1_v3_0Inst_0_n2 , Red_MCInst2_MC1_v3_2Inst_0_n2 ,
         Red_MCInst2_MC1_r0Inst_XORInst_0_0_n5 ,
         Red_MCInst2_MC1_r0Inst_XORInst_0_0_n4 ,
         Red_MCInst2_MC1_r1Inst_XORInst_0_0_n5 ,
         Red_MCInst2_MC1_r1Inst_XORInst_0_0_n4 ,
         Red_MCInst2_MC1_r2Inst_XORInst_0_0_n5 ,
         Red_MCInst2_MC1_r2Inst_XORInst_0_0_n4 ,
         Red_MCInst2_MC1_r3Inst_XORInst_0_0_n5 ,
         Red_MCInst2_MC1_r3Inst_XORInst_0_0_n4 , Red_MCInst2_MC2_v3_3[0] ,
         Red_MCInst2_MC2_v3_2[0] , Red_MCInst2_MC2_v3_1[0] ,
         Red_MCInst2_MC2_v3_0[0] , Red_MCInst2_MC2_v2_3[0] ,
         Red_MCInst2_MC2_v2_2[0] , Red_MCInst2_MC2_v2_1[0] ,
         Red_MCInst2_MC2_v2_0[0] , Red_MCInst2_MC2_v1_3[0] ,
         Red_MCInst2_MC2_v1_2[0] , Red_MCInst2_MC2_v1_1[0] ,
         Red_MCInst2_MC2_v1_0[0] , Red_MCInst2_MC2_v0_3[0] ,
         Red_MCInst2_MC2_v0_2[0] , Red_MCInst2_MC2_v0_1[0] ,
         Red_MCInst2_MC2_v0_0[0] , Red_MCInst2_MC2_v0_3Inst_0_n2 ,
         Red_MCInst2_MC2_v1_0Inst_0_n4 , Red_MCInst2_MC2_v1_0Inst_0_n3 ,
         Red_MCInst2_MC2_v1_3Inst_0_n2 , Red_MCInst2_MC2_v2_0Inst_0_n2 ,
         Red_MCInst2_MC2_v3_0Inst_0_n2 , Red_MCInst2_MC2_v3_2Inst_0_n2 ,
         Red_MCInst2_MC2_r0Inst_XORInst_0_0_n5 ,
         Red_MCInst2_MC2_r0Inst_XORInst_0_0_n4 ,
         Red_MCInst2_MC2_r1Inst_XORInst_0_0_n5 ,
         Red_MCInst2_MC2_r1Inst_XORInst_0_0_n4 ,
         Red_MCInst2_MC2_r2Inst_XORInst_0_0_n5 ,
         Red_MCInst2_MC2_r2Inst_XORInst_0_0_n4 ,
         Red_MCInst2_MC2_r3Inst_XORInst_0_0_n5 ,
         Red_MCInst2_MC2_r3Inst_XORInst_0_0_n4 , Red_MCInst2_MC3_v3_3[0] ,
         Red_MCInst2_MC3_v3_2[0] , Red_MCInst2_MC3_v3_1[0] ,
         Red_MCInst2_MC3_v3_0[0] , Red_MCInst2_MC3_v2_3[0] ,
         Red_MCInst2_MC3_v2_2[0] , Red_MCInst2_MC3_v2_1[0] ,
         Red_MCInst2_MC3_v2_0[0] , Red_MCInst2_MC3_v1_3[0] ,
         Red_MCInst2_MC3_v1_2[0] , Red_MCInst2_MC3_v1_1[0] ,
         Red_MCInst2_MC3_v1_0[0] , Red_MCInst2_MC3_v0_3[0] ,
         Red_MCInst2_MC3_v0_2[0] , Red_MCInst2_MC3_v0_1[0] ,
         Red_MCInst2_MC3_v0_0[0] , Red_MCInst2_MC3_v0_3Inst_0_n2 ,
         Red_MCInst2_MC3_v1_0Inst_0_n4 , Red_MCInst2_MC3_v1_0Inst_0_n3 ,
         Red_MCInst2_MC3_v1_3Inst_0_n2 , Red_MCInst2_MC3_v2_0Inst_0_n2 ,
         Red_MCInst2_MC3_v3_0Inst_0_n2 , Red_MCInst2_MC3_v3_2Inst_0_n2 ,
         Red_MCInst2_MC3_r0Inst_XORInst_0_0_n5 ,
         Red_MCInst2_MC3_r0Inst_XORInst_0_0_n4 ,
         Red_MCInst2_MC3_r1Inst_XORInst_0_0_n5 ,
         Red_MCInst2_MC3_r1Inst_XORInst_0_0_n4 ,
         Red_MCInst2_MC3_r2Inst_XORInst_0_0_n5 ,
         Red_MCInst2_MC3_r2Inst_XORInst_0_0_n4 ,
         Red_MCInst2_MC3_r3Inst_XORInst_0_0_n5 ,
         Red_MCInst2_MC3_r3Inst_XORInst_0_0_n4 ,
         Red_SubCellInst3_LFInst_0_LFInst_0_n6 ,
         Red_SubCellInst3_LFInst_0_LFInst_0_n5 ,
         Red_SubCellInst3_LFInst_0_LFInst_0_n4 ,
         Red_SubCellInst3_LFInst_1_LFInst_0_n6 ,
         Red_SubCellInst3_LFInst_1_LFInst_0_n5 ,
         Red_SubCellInst3_LFInst_1_LFInst_0_n4 ,
         Red_SubCellInst3_LFInst_2_LFInst_0_n6 ,
         Red_SubCellInst3_LFInst_2_LFInst_0_n5 ,
         Red_SubCellInst3_LFInst_2_LFInst_0_n4 ,
         Red_SubCellInst3_LFInst_3_LFInst_0_n6 ,
         Red_SubCellInst3_LFInst_3_LFInst_0_n5 ,
         Red_SubCellInst3_LFInst_3_LFInst_0_n4 ,
         Red_SubCellInst3_LFInst_4_LFInst_0_n6 ,
         Red_SubCellInst3_LFInst_4_LFInst_0_n5 ,
         Red_SubCellInst3_LFInst_4_LFInst_0_n4 ,
         Red_SubCellInst3_LFInst_5_LFInst_0_n6 ,
         Red_SubCellInst3_LFInst_5_LFInst_0_n5 ,
         Red_SubCellInst3_LFInst_5_LFInst_0_n4 ,
         Red_SubCellInst3_LFInst_6_LFInst_0_n6 ,
         Red_SubCellInst3_LFInst_6_LFInst_0_n5 ,
         Red_SubCellInst3_LFInst_6_LFInst_0_n4 ,
         Red_SubCellInst3_LFInst_7_LFInst_0_n6 ,
         Red_SubCellInst3_LFInst_7_LFInst_0_n5 ,
         Red_SubCellInst3_LFInst_7_LFInst_0_n4 ,
         Red_SubCellInst3_LFInst_8_LFInst_0_n6 ,
         Red_SubCellInst3_LFInst_8_LFInst_0_n5 ,
         Red_SubCellInst3_LFInst_8_LFInst_0_n4 ,
         Red_SubCellInst3_LFInst_9_LFInst_0_n6 ,
         Red_SubCellInst3_LFInst_9_LFInst_0_n5 ,
         Red_SubCellInst3_LFInst_9_LFInst_0_n4 ,
         Red_SubCellInst3_LFInst_10_LFInst_0_n6 ,
         Red_SubCellInst3_LFInst_10_LFInst_0_n5 ,
         Red_SubCellInst3_LFInst_10_LFInst_0_n4 ,
         Red_SubCellInst3_LFInst_11_LFInst_0_n6 ,
         Red_SubCellInst3_LFInst_11_LFInst_0_n5 ,
         Red_SubCellInst3_LFInst_11_LFInst_0_n4 ,
         Red_SubCellInst3_LFInst_12_LFInst_0_n6 ,
         Red_SubCellInst3_LFInst_12_LFInst_0_n5 ,
         Red_SubCellInst3_LFInst_12_LFInst_0_n4 ,
         Red_SubCellInst3_LFInst_13_LFInst_0_n6 ,
         Red_SubCellInst3_LFInst_13_LFInst_0_n5 ,
         Red_SubCellInst3_LFInst_13_LFInst_0_n4 ,
         Red_SubCellInst3_LFInst_14_LFInst_0_n6 ,
         Red_SubCellInst3_LFInst_14_LFInst_0_n5 ,
         Red_SubCellInst3_LFInst_14_LFInst_0_n4 ,
         Red_SubCellInst3_LFInst_15_LFInst_0_n6 ,
         Red_SubCellInst3_LFInst_15_LFInst_0_n5 ,
         Red_SubCellInst3_LFInst_15_LFInst_0_n4 , Red_MCInst3_MC0_v3_3[0] ,
         Red_MCInst3_MC0_v3_2[0] , Red_MCInst3_MC0_v3_1[0] ,
         Red_MCInst3_MC0_v3_0[0] , Red_MCInst3_MC0_v2_3[0] ,
         Red_MCInst3_MC0_v2_2[0] , Red_MCInst3_MC0_v2_1[0] ,
         Red_MCInst3_MC0_v2_0[0] , Red_MCInst3_MC0_v1_3[0] ,
         Red_MCInst3_MC0_v1_2[0] , Red_MCInst3_MC0_v1_1[0] ,
         Red_MCInst3_MC0_v1_0[0] , Red_MCInst3_MC0_v0_3[0] ,
         Red_MCInst3_MC0_v0_2[0] , Red_MCInst3_MC0_v0_1[0] ,
         Red_MCInst3_MC0_v0_0[0] , Red_MCInst3_MC0_v0_3Inst_0_n2 ,
         Red_MCInst3_MC0_v1_0Inst_0_n4 , Red_MCInst3_MC0_v1_0Inst_0_n3 ,
         Red_MCInst3_MC0_v1_3Inst_0_n2 , Red_MCInst3_MC0_v2_0Inst_0_n2 ,
         Red_MCInst3_MC0_v3_0Inst_0_n2 , Red_MCInst3_MC0_v3_2Inst_0_n2 ,
         Red_MCInst3_MC0_r0Inst_XORInst_0_0_n5 ,
         Red_MCInst3_MC0_r0Inst_XORInst_0_0_n4 ,
         Red_MCInst3_MC0_r1Inst_XORInst_0_0_n5 ,
         Red_MCInst3_MC0_r1Inst_XORInst_0_0_n4 ,
         Red_MCInst3_MC0_r2Inst_XORInst_0_0_n5 ,
         Red_MCInst3_MC0_r2Inst_XORInst_0_0_n4 ,
         Red_MCInst3_MC0_r3Inst_XORInst_0_0_n5 ,
         Red_MCInst3_MC0_r3Inst_XORInst_0_0_n4 , Red_MCInst3_MC1_v3_3[0] ,
         Red_MCInst3_MC1_v3_2[0] , Red_MCInst3_MC1_v3_1[0] ,
         Red_MCInst3_MC1_v3_0[0] , Red_MCInst3_MC1_v2_3[0] ,
         Red_MCInst3_MC1_v2_2[0] , Red_MCInst3_MC1_v2_1[0] ,
         Red_MCInst3_MC1_v2_0[0] , Red_MCInst3_MC1_v1_3[0] ,
         Red_MCInst3_MC1_v1_2[0] , Red_MCInst3_MC1_v1_1[0] ,
         Red_MCInst3_MC1_v1_0[0] , Red_MCInst3_MC1_v0_3[0] ,
         Red_MCInst3_MC1_v0_2[0] , Red_MCInst3_MC1_v0_1[0] ,
         Red_MCInst3_MC1_v0_0[0] , Red_MCInst3_MC1_v0_3Inst_0_n2 ,
         Red_MCInst3_MC1_v1_0Inst_0_n4 , Red_MCInst3_MC1_v1_0Inst_0_n3 ,
         Red_MCInst3_MC1_v1_3Inst_0_n2 , Red_MCInst3_MC1_v2_0Inst_0_n2 ,
         Red_MCInst3_MC1_v3_0Inst_0_n2 , Red_MCInst3_MC1_v3_2Inst_0_n2 ,
         Red_MCInst3_MC1_r0Inst_XORInst_0_0_n5 ,
         Red_MCInst3_MC1_r0Inst_XORInst_0_0_n4 ,
         Red_MCInst3_MC1_r1Inst_XORInst_0_0_n5 ,
         Red_MCInst3_MC1_r1Inst_XORInst_0_0_n4 ,
         Red_MCInst3_MC1_r2Inst_XORInst_0_0_n5 ,
         Red_MCInst3_MC1_r2Inst_XORInst_0_0_n4 ,
         Red_MCInst3_MC1_r3Inst_XORInst_0_0_n5 ,
         Red_MCInst3_MC1_r3Inst_XORInst_0_0_n4 , Red_MCInst3_MC2_v3_3[0] ,
         Red_MCInst3_MC2_v3_2[0] , Red_MCInst3_MC2_v3_1[0] ,
         Red_MCInst3_MC2_v3_0[0] , Red_MCInst3_MC2_v2_3[0] ,
         Red_MCInst3_MC2_v2_2[0] , Red_MCInst3_MC2_v2_1[0] ,
         Red_MCInst3_MC2_v2_0[0] , Red_MCInst3_MC2_v1_3[0] ,
         Red_MCInst3_MC2_v1_2[0] , Red_MCInst3_MC2_v1_1[0] ,
         Red_MCInst3_MC2_v1_0[0] , Red_MCInst3_MC2_v0_3[0] ,
         Red_MCInst3_MC2_v0_2[0] , Red_MCInst3_MC2_v0_1[0] ,
         Red_MCInst3_MC2_v0_0[0] , Red_MCInst3_MC2_v0_3Inst_0_n2 ,
         Red_MCInst3_MC2_v1_0Inst_0_n4 , Red_MCInst3_MC2_v1_0Inst_0_n3 ,
         Red_MCInst3_MC2_v1_3Inst_0_n2 , Red_MCInst3_MC2_v2_0Inst_0_n2 ,
         Red_MCInst3_MC2_v3_0Inst_0_n2 , Red_MCInst3_MC2_v3_2Inst_0_n2 ,
         Red_MCInst3_MC2_r0Inst_XORInst_0_0_n5 ,
         Red_MCInst3_MC2_r0Inst_XORInst_0_0_n4 ,
         Red_MCInst3_MC2_r1Inst_XORInst_0_0_n5 ,
         Red_MCInst3_MC2_r1Inst_XORInst_0_0_n4 ,
         Red_MCInst3_MC2_r2Inst_XORInst_0_0_n5 ,
         Red_MCInst3_MC2_r2Inst_XORInst_0_0_n4 ,
         Red_MCInst3_MC2_r3Inst_XORInst_0_0_n5 ,
         Red_MCInst3_MC2_r3Inst_XORInst_0_0_n4 , Red_MCInst3_MC3_v3_3[0] ,
         Red_MCInst3_MC3_v3_2[0] , Red_MCInst3_MC3_v3_1[0] ,
         Red_MCInst3_MC3_v3_0[0] , Red_MCInst3_MC3_v2_3[0] ,
         Red_MCInst3_MC3_v2_2[0] , Red_MCInst3_MC3_v2_1[0] ,
         Red_MCInst3_MC3_v2_0[0] , Red_MCInst3_MC3_v1_3[0] ,
         Red_MCInst3_MC3_v1_2[0] , Red_MCInst3_MC3_v1_1[0] ,
         Red_MCInst3_MC3_v1_0[0] , Red_MCInst3_MC3_v0_3[0] ,
         Red_MCInst3_MC3_v0_2[0] , Red_MCInst3_MC3_v0_1[0] ,
         Red_MCInst3_MC3_v0_0[0] , Red_MCInst3_MC3_v0_3Inst_0_n2 ,
         Red_MCInst3_MC3_v1_0Inst_0_n4 , Red_MCInst3_MC3_v1_0Inst_0_n3 ,
         Red_MCInst3_MC3_v1_3Inst_0_n2 , Red_MCInst3_MC3_v2_0Inst_0_n2 ,
         Red_MCInst3_MC3_v3_0Inst_0_n2 , Red_MCInst3_MC3_v3_2Inst_0_n2 ,
         Red_MCInst3_MC3_r0Inst_XORInst_0_0_n5 ,
         Red_MCInst3_MC3_r0Inst_XORInst_0_0_n4 ,
         Red_MCInst3_MC3_r1Inst_XORInst_0_0_n5 ,
         Red_MCInst3_MC3_r1Inst_XORInst_0_0_n4 ,
         Red_MCInst3_MC3_r2Inst_XORInst_0_0_n5 ,
         Red_MCInst3_MC3_r2Inst_XORInst_0_0_n4 ,
         Red_MCInst3_MC3_r3Inst_XORInst_0_0_n5 ,
         Red_MCInst3_MC3_r3Inst_XORInst_0_0_n4 ,
         Red_KeyInst_LFInst_0_LFInst_0_n4 ,
         Red_KeyInst_LFInst_0_LFInst_0_n3 ,
         Red_KeyInst_LFInst_1_LFInst_0_n4 ,
         Red_KeyInst_LFInst_1_LFInst_0_n3 ,
         Red_KeyInst_LFInst_2_LFInst_0_n4 ,
         Red_KeyInst_LFInst_2_LFInst_0_n3 ,
         Red_KeyInst_LFInst_3_LFInst_0_n4 ,
         Red_KeyInst_LFInst_3_LFInst_0_n3 ,
         Red_KeyInst_LFInst_4_LFInst_0_n4 ,
         Red_KeyInst_LFInst_4_LFInst_0_n3 ,
         Red_KeyInst_LFInst_5_LFInst_0_n4 ,
         Red_KeyInst_LFInst_5_LFInst_0_n3 ,
         Red_KeyInst_LFInst_6_LFInst_0_n4 ,
         Red_KeyInst_LFInst_6_LFInst_0_n3 ,
         Red_KeyInst_LFInst_7_LFInst_0_n4 ,
         Red_KeyInst_LFInst_7_LFInst_0_n3 ,
         Red_KeyInst_LFInst_8_LFInst_0_n4 ,
         Red_KeyInst_LFInst_8_LFInst_0_n3 ,
         Red_KeyInst_LFInst_9_LFInst_0_n4 ,
         Red_KeyInst_LFInst_9_LFInst_0_n3 ,
         Red_KeyInst_LFInst_10_LFInst_0_n4 ,
         Red_KeyInst_LFInst_10_LFInst_0_n3 ,
         Red_KeyInst_LFInst_11_LFInst_0_n4 ,
         Red_KeyInst_LFInst_11_LFInst_0_n3 ,
         Red_KeyInst_LFInst_12_LFInst_0_n4 ,
         Red_KeyInst_LFInst_12_LFInst_0_n3 ,
         Red_KeyInst_LFInst_13_LFInst_0_n4 ,
         Red_KeyInst_LFInst_13_LFInst_0_n3 ,
         Red_KeyInst_LFInst_14_LFInst_0_n4 ,
         Red_KeyInst_LFInst_14_LFInst_0_n3 ,
         Red_KeyInst_LFInst_15_LFInst_0_n4 ,
         Red_KeyInst_LFInst_15_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_0_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_0_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_1_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_1_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_2_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_2_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_3_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_3_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_4_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_4_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_5_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_5_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_6_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_6_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_7_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_7_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_8_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_8_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_9_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_9_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_10_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_10_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_11_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_11_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_12_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_12_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_13_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_13_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_14_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_14_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_15_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_15_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_16_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_16_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_17_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_17_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_18_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_18_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_19_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_19_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_20_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_20_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_21_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_21_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_22_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_22_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_23_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_23_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_24_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_24_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_25_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_25_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_26_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_26_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_27_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_27_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_28_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_28_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_29_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_29_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_30_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_30_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_31_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_31_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_32_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_32_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_33_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_33_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_34_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_34_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_35_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_35_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_36_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_36_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_37_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_37_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_38_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_38_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_39_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_39_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_40_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_40_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_41_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_41_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_42_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_42_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_43_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_43_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_44_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_44_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_45_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_45_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_46_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_46_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_47_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_47_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_48_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_48_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_49_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_49_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_50_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_50_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_51_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_51_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_52_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_52_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_53_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_53_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_54_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_54_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_55_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_55_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_56_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_56_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_57_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_57_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_58_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_58_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_59_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_59_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_60_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_60_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_61_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_61_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_62_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_62_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_63_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_63_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_64_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_64_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_65_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_65_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_66_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_66_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_67_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_67_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_68_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_68_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_69_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_69_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_70_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_70_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_71_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_71_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_72_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_72_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_73_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_73_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_74_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_74_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_75_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_75_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_76_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_76_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_77_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_77_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_78_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_78_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_79_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_79_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_80_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_80_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_81_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_81_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_82_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_82_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_83_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_83_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_84_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_84_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_85_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_85_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_86_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_86_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_87_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_87_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_88_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_88_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_89_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_89_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_90_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_90_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_91_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_91_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_92_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_92_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_93_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_93_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_94_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_94_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_95_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_95_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_96_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_96_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_97_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_97_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_98_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_98_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_99_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_99_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_100_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_100_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_101_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_101_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_102_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_102_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_103_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_103_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_104_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_104_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_105_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_105_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_106_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_106_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_107_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_107_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_108_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_108_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_109_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_109_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_110_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_110_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_111_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_111_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_112_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_112_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_113_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_113_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_114_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_114_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_115_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_115_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_116_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_116_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_117_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_117_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_118_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_118_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_119_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_119_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_120_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_120_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_121_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_121_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_122_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_122_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_123_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_123_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_124_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_124_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_125_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_125_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_126_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_126_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_127_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_127_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_128_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_128_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_129_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_129_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_130_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_130_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_131_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_131_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_132_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_132_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_133_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_133_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_134_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_134_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_135_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_135_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_136_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_136_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_137_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_137_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_138_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_138_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_139_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_139_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_140_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_140_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_141_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_141_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_142_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_142_LFInst_0_n3 ,
         Red_ToCheckInst_LFInst_143_LFInst_0_n4 ,
         Red_ToCheckInst_LFInst_143_LFInst_0_n3 , Check1_CheckInst_0_n286 ,
         Check1_CheckInst_0_n285 , Check1_CheckInst_0_n284 ,
         Check1_CheckInst_0_n283 , Check1_CheckInst_0_n282 ,
         Check1_CheckInst_0_n281 , Check1_CheckInst_0_n280 ,
         Check1_CheckInst_0_n279 , Check1_CheckInst_0_n278 ,
         Check1_CheckInst_0_n277 , Check1_CheckInst_0_n276 ,
         Check1_CheckInst_0_n275 , Check1_CheckInst_0_n274 ,
         Check1_CheckInst_0_n273 , Check1_CheckInst_0_n272 ,
         Check1_CheckInst_0_n271 , Check1_CheckInst_0_n270 ,
         Check1_CheckInst_0_n269 , Check1_CheckInst_0_n268 ,
         Check1_CheckInst_0_n267 , Check1_CheckInst_0_n266 ,
         Check1_CheckInst_0_n265 , Check1_CheckInst_0_n264 ,
         Check1_CheckInst_0_n263 , Check1_CheckInst_0_n262 ,
         Check1_CheckInst_0_n261 , Check1_CheckInst_0_n260 ,
         Check1_CheckInst_0_n259 , Check1_CheckInst_0_n258 ,
         Check1_CheckInst_0_n257 , Check1_CheckInst_0_n256 ,
         Check1_CheckInst_0_n255 , Check1_CheckInst_0_n254 ,
         Check1_CheckInst_0_n253 , Check1_CheckInst_0_n252 ,
         Check1_CheckInst_0_n251 , Check1_CheckInst_0_n250 ,
         Check1_CheckInst_0_n249 , Check1_CheckInst_0_n248 ,
         Check1_CheckInst_0_n247 , Check1_CheckInst_0_n246 ,
         Check1_CheckInst_0_n245 , Check1_CheckInst_0_n244 ,
         Check1_CheckInst_0_n243 , Check1_CheckInst_0_n242 ,
         Check1_CheckInst_0_n241 , Check1_CheckInst_0_n240 ,
         Check1_CheckInst_0_n239 , Check1_CheckInst_0_n238 ,
         Check1_CheckInst_0_n237 , Check1_CheckInst_0_n236 ,
         Check1_CheckInst_0_n235 , Check1_CheckInst_0_n234 ,
         Check1_CheckInst_0_n233 , Check1_CheckInst_0_n232 ,
         Check1_CheckInst_0_n231 , Check1_CheckInst_0_n230 ,
         Check1_CheckInst_0_n229 , Check1_CheckInst_0_n228 ,
         Check1_CheckInst_0_n227 , Check1_CheckInst_0_n226 ,
         Check1_CheckInst_0_n225 , Check1_CheckInst_0_n224 ,
         Check1_CheckInst_0_n223 , Check1_CheckInst_0_n222 ,
         Check1_CheckInst_0_n221 , Check1_CheckInst_0_n220 ,
         Check1_CheckInst_0_n219 , Check1_CheckInst_0_n218 ,
         Check1_CheckInst_0_n217 , Check1_CheckInst_0_n216 ,
         Check1_CheckInst_0_n215 , Check1_CheckInst_0_n214 ,
         Check1_CheckInst_0_n213 , Check1_CheckInst_0_n212 ,
         Check1_CheckInst_0_n211 , Check1_CheckInst_0_n210 ,
         Check1_CheckInst_0_n209 , Check1_CheckInst_0_n208 ,
         Check1_CheckInst_0_n207 , Check1_CheckInst_0_n206 ,
         Check1_CheckInst_0_n205 , Check1_CheckInst_0_n204 ,
         Check1_CheckInst_0_n203 , Check1_CheckInst_0_n202 ,
         Check1_CheckInst_0_n201 , Check1_CheckInst_0_n200 ,
         Check1_CheckInst_0_n199 , Check1_CheckInst_0_n198 ,
         Check1_CheckInst_0_n197 , Check1_CheckInst_0_n196 ,
         Check1_CheckInst_0_n195 , Check1_CheckInst_0_n194 ,
         Check1_CheckInst_0_n193 , Check1_CheckInst_0_n192 ,
         Check1_CheckInst_0_n191 , Check1_CheckInst_0_n190 ,
         Check1_CheckInst_0_n189 , Check1_CheckInst_0_n188 ,
         Check1_CheckInst_0_n187 , Check1_CheckInst_0_n186 ,
         Check1_CheckInst_0_n185 , Check1_CheckInst_0_n184 ,
         Check1_CheckInst_0_n183 , Check1_CheckInst_0_n182 ,
         Check1_CheckInst_0_n181 , Check1_CheckInst_0_n180 ,
         Check1_CheckInst_0_n179 , Check1_CheckInst_0_n178 ,
         Check1_CheckInst_0_n177 , Check1_CheckInst_0_n176 ,
         Check1_CheckInst_0_n175 , Check1_CheckInst_0_n174 ,
         Check1_CheckInst_0_n173 , Check1_CheckInst_0_n172 ,
         Check1_CheckInst_0_n171 , Check1_CheckInst_0_n170 ,
         Check1_CheckInst_0_n169 , Check1_CheckInst_0_n168 ,
         Check1_CheckInst_0_n167 , Check1_CheckInst_0_n166 ,
         Check1_CheckInst_0_n165 , Check1_CheckInst_0_n164 ,
         Check1_CheckInst_0_n163 , Check1_CheckInst_0_n162 ,
         Check1_CheckInst_0_n161 , Check1_CheckInst_0_n160 ,
         Check1_CheckInst_0_n159 , Check1_CheckInst_0_n158 ,
         Check1_CheckInst_0_n157 , Check1_CheckInst_0_n156 ,
         Check1_CheckInst_0_n155 , Check1_CheckInst_0_n154 ,
         Check1_CheckInst_0_n153 , Check1_CheckInst_0_n152 ,
         Check1_CheckInst_0_n151 , Check1_CheckInst_0_n150 ,
         Check1_CheckInst_0_n149 , Check1_CheckInst_0_n148 ,
         Check1_CheckInst_0_n147 , Check1_CheckInst_0_n146 ,
         Check1_CheckInst_0_n145 , Check1_CheckInst_0_n144 ,
         Check1_CheckInst_0_n143 , Check1_CheckInst_0_n142 ,
         Check1_CheckInst_0_n141 , Check1_CheckInst_0_n140 ,
         Check1_CheckInst_0_n139 , Check1_CheckInst_0_n138 ,
         Check1_CheckInst_0_n137 , Check1_CheckInst_0_n136 ,
         Check1_CheckInst_0_n135 , Check1_CheckInst_0_n134 ,
         Check1_CheckInst_0_n133 , Check1_CheckInst_0_n132 ,
         Check1_CheckInst_0_n131 , Check1_CheckInst_0_n130 ,
         Check1_CheckInst_0_n129 , Check1_CheckInst_0_n128 ,
         Check1_CheckInst_0_n127 , Check1_CheckInst_0_n126 ,
         Check1_CheckInst_0_n125 , Check1_CheckInst_0_n124 ,
         Check1_CheckInst_0_n123 , Check1_CheckInst_0_n122 ,
         Check1_CheckInst_0_n121 , Check1_CheckInst_0_n120 ,
         Check1_CheckInst_0_n119 , Check1_CheckInst_0_n118 ,
         Check1_CheckInst_0_n117 , Check1_CheckInst_0_n116 ,
         Check1_CheckInst_0_n115 , Check1_CheckInst_0_n114 ,
         Check1_CheckInst_0_n113 , Check1_CheckInst_0_n112 ,
         Check1_CheckInst_0_n111 , Check1_CheckInst_0_n110 ,
         Check1_CheckInst_0_n109 , Check1_CheckInst_0_n108 ,
         Check1_CheckInst_0_n107 , Check1_CheckInst_0_n106 ,
         Check1_CheckInst_0_n105 , Check1_CheckInst_0_n104 ,
         Check1_CheckInst_0_n103 , Check1_CheckInst_0_n102 ,
         Check1_CheckInst_0_n101 , Check1_CheckInst_0_n100 ,
         Check1_CheckInst_0_n99 , Check1_CheckInst_0_n98 ,
         Check1_CheckInst_0_n97 , Check1_CheckInst_0_n96 ,
         Check1_CheckInst_0_n95 , Check1_CheckInst_0_n94 ,
         Check1_CheckInst_0_n93 , Check1_CheckInst_0_n92 ,
         Check1_CheckInst_0_n91 , Check1_CheckInst_0_n90 ,
         Check1_CheckInst_0_n89 , Check1_CheckInst_0_n88 ,
         Check1_CheckInst_0_n87 , Check1_CheckInst_0_n86 ,
         Check1_CheckInst_0_n85 , Check1_CheckInst_0_n84 ,
         Check1_CheckInst_0_n83 , Check1_CheckInst_0_n82 ,
         Check1_CheckInst_0_n81 , Check1_CheckInst_0_n80 ,
         Check1_CheckInst_0_n79 , Check1_CheckInst_0_n78 ,
         Check1_CheckInst_0_n77 , Check1_CheckInst_0_n76 ,
         Check1_CheckInst_0_n75 , Check1_CheckInst_0_n74 ,
         Check1_CheckInst_0_n73 , Check1_CheckInst_0_n72 ,
         Check1_CheckInst_0_n71 , Check1_CheckInst_0_n70 ,
         Check1_CheckInst_0_n69 , Check1_CheckInst_0_n68 ,
         Check1_CheckInst_0_n67 , Check1_CheckInst_0_n66 ,
         Check1_CheckInst_0_n65 , Check1_CheckInst_0_n64 ,
         Check1_CheckInst_0_n63 , Check1_CheckInst_0_n62 ,
         Check1_CheckInst_0_n61 , Check1_CheckInst_0_n60 ,
         Check1_CheckInst_0_n59 , Check1_CheckInst_0_n58 ,
         Check1_CheckInst_0_n57 , Check1_CheckInst_0_n56 ,
         Check1_CheckInst_0_n55 , Check1_CheckInst_0_n54 ,
         Check1_CheckInst_0_n53 , Check1_CheckInst_0_n52 ,
         Check1_CheckInst_0_n51 , Check1_CheckInst_0_n50 ,
         Check1_CheckInst_0_n49 , Check1_CheckInst_0_n48 ,
         Check1_CheckInst_0_n47 , Check1_CheckInst_0_n46 ,
         Check1_CheckInst_0_n45 , Check1_CheckInst_0_n44 ,
         Check1_CheckInst_0_n43 , Check1_CheckInst_0_n42 ,
         Check1_CheckInst_0_n41 , Check1_CheckInst_0_n40 ,
         Check1_CheckInst_0_n39 , Check1_CheckInst_0_n38 ,
         Check1_CheckInst_0_n37 , Check1_CheckInst_0_n36 ,
         Check1_CheckInst_0_n35 , Check1_CheckInst_0_n34 ,
         Check1_CheckInst_0_n33 , Check1_CheckInst_0_n32 ,
         Check1_CheckInst_0_n31 , Check1_CheckInst_0_n30 ,
         Check1_CheckInst_0_n29 , Check1_CheckInst_0_n28 ,
         Check1_CheckInst_0_n27 , Check1_CheckInst_0_n26 ,
         Check1_CheckInst_0_n25 , Check1_CheckInst_0_n24 ,
         Check1_CheckInst_0_n23 , Check1_CheckInst_0_n22 ,
         Check1_CheckInst_0_n21 , Check1_CheckInst_0_n20 ,
         Check1_CheckInst_0_n19 , Check1_CheckInst_0_n18 ,
         Check1_CheckInst_0_n17 , Check1_CheckInst_0_n16 ,
         Check1_CheckInst_0_n15 , Check1_CheckInst_0_n14 ,
         Check1_CheckInst_0_n13 , Check1_CheckInst_0_n12 ,
         Check1_CheckInst_0_n11 , Check1_CheckInst_0_n10 ,
         Check1_CheckInst_0_n9 , Check1_CheckInst_0_n8 ,
         Check1_CheckInst_0_n7 , Check1_CheckInst_0_n6 ,
         Check1_CheckInst_0_n5 , Check1_CheckInst_0_n4 ,
         Check1_CheckInst_0_n3 , Check1_CheckInst_0_n2 ,
         Check1_CheckInst_0_n1 ;
  wire   [63:0] AddRoundKeyOutput;
  wire   [63:0] Feedback;
  wire   [63:0] SubCellInput;
  wire   [63:0] Feedback2;
  wire   [63:0] SubCellInput2;
  wire   [15:0] Red_Plaintext;
  wire   [15:0] Red_RoundKey;
  wire   [15:0] Red_AddRoundKeyOutput;
  wire   [15:0] Red_ShiftRowsOutput;
  wire   [15:0] Red_Feedback;
  wire   [15:0] Red_SubCellInput;
  wire   [15:0] Red_ShiftRowsOutput2;
  wire   [15:0] Red_Feedback2;
  wire   [15:0] Red_SubCellInput2;
  wire   [15:0] Red_ShiftRowsOutput3;
  wire   [15:0] Red_Feedback3;
  wire   [143:0] Red_SignaltoCheck;
  wire   [3:0] MCInst_MC0_v3_3 ;
  wire   [3:0] MCInst_MC0_v3_2 ;
  wire   [3:0] MCInst_MC0_v3_1 ;
  wire   [3:0] MCInst_MC0_v3_0 ;
  wire   [3:0] MCInst_MC0_v2_3 ;
  wire   [3:0] MCInst_MC0_v2_2 ;
  wire   [3:0] MCInst_MC0_v2_1 ;
  wire   [3:0] MCInst_MC0_v2_0 ;
  wire   [3:0] MCInst_MC0_v1_3 ;
  wire   [3:0] MCInst_MC0_v1_2 ;
  wire   [3:0] MCInst_MC0_v1_1 ;
  wire   [3:0] MCInst_MC0_v1_0 ;
  wire   [3:0] MCInst_MC0_v0_3 ;
  wire   [3:0] MCInst_MC0_v0_2 ;
  wire   [3:0] MCInst_MC0_v0_1 ;
  wire   [3:0] MCInst_MC0_v0_0 ;
  wire   [3:0] MCInst_MC1_v3_3 ;
  wire   [3:0] MCInst_MC1_v3_2 ;
  wire   [3:0] MCInst_MC1_v3_1 ;
  wire   [3:0] MCInst_MC1_v3_0 ;
  wire   [3:0] MCInst_MC1_v2_3 ;
  wire   [3:0] MCInst_MC1_v2_2 ;
  wire   [3:0] MCInst_MC1_v2_1 ;
  wire   [3:0] MCInst_MC1_v2_0 ;
  wire   [3:0] MCInst_MC1_v1_3 ;
  wire   [3:0] MCInst_MC1_v1_2 ;
  wire   [3:0] MCInst_MC1_v1_1 ;
  wire   [3:0] MCInst_MC1_v1_0 ;
  wire   [3:0] MCInst_MC1_v0_3 ;
  wire   [3:0] MCInst_MC1_v0_2 ;
  wire   [3:0] MCInst_MC1_v0_1 ;
  wire   [3:0] MCInst_MC1_v0_0 ;
  wire   [3:0] MCInst_MC2_v3_3 ;
  wire   [3:0] MCInst_MC2_v3_2 ;
  wire   [3:0] MCInst_MC2_v3_1 ;
  wire   [3:0] MCInst_MC2_v3_0 ;
  wire   [3:0] MCInst_MC2_v2_3 ;
  wire   [3:0] MCInst_MC2_v2_2 ;
  wire   [3:0] MCInst_MC2_v2_1 ;
  wire   [3:0] MCInst_MC2_v2_0 ;
  wire   [3:0] MCInst_MC2_v1_3 ;
  wire   [3:0] MCInst_MC2_v1_2 ;
  wire   [3:0] MCInst_MC2_v1_1 ;
  wire   [3:0] MCInst_MC2_v1_0 ;
  wire   [3:0] MCInst_MC2_v0_3 ;
  wire   [3:0] MCInst_MC2_v0_2 ;
  wire   [3:0] MCInst_MC2_v0_1 ;
  wire   [3:0] MCInst_MC2_v0_0 ;
  wire   [3:0] MCInst_MC3_v3_3 ;
  wire   [3:0] MCInst_MC3_v3_2 ;
  wire   [3:0] MCInst_MC3_v3_1 ;
  wire   [3:0] MCInst_MC3_v3_0 ;
  wire   [3:0] MCInst_MC3_v2_3 ;
  wire   [3:0] MCInst_MC3_v2_2 ;
  wire   [3:0] MCInst_MC3_v2_1 ;
  wire   [3:0] MCInst_MC3_v2_0 ;
  wire   [3:0] MCInst_MC3_v1_3 ;
  wire   [3:0] MCInst_MC3_v1_2 ;
  wire   [3:0] MCInst_MC3_v1_1 ;
  wire   [3:0] MCInst_MC3_v1_0 ;
  wire   [3:0] MCInst_MC3_v0_3 ;
  wire   [3:0] MCInst_MC3_v0_2 ;
  wire   [3:0] MCInst_MC3_v0_1 ;
  wire   [3:0] MCInst_MC3_v0_0 ;
  wire   [3:0] MCInst2_MC0_v3_3 ;
  wire   [3:0] MCInst2_MC0_v3_2 ;
  wire   [3:0] MCInst2_MC0_v3_1 ;
  wire   [3:0] MCInst2_MC0_v3_0 ;
  wire   [3:0] MCInst2_MC0_v2_3 ;
  wire   [3:0] MCInst2_MC0_v2_2 ;
  wire   [3:0] MCInst2_MC0_v2_1 ;
  wire   [3:0] MCInst2_MC0_v2_0 ;
  wire   [3:0] MCInst2_MC0_v1_3 ;
  wire   [3:0] MCInst2_MC0_v1_2 ;
  wire   [3:0] MCInst2_MC0_v1_1 ;
  wire   [3:0] MCInst2_MC0_v1_0 ;
  wire   [3:0] MCInst2_MC0_v0_3 ;
  wire   [3:0] MCInst2_MC0_v0_2 ;
  wire   [3:0] MCInst2_MC0_v0_1 ;
  wire   [3:0] MCInst2_MC0_v0_0 ;
  wire   [3:0] MCInst2_MC1_v3_3 ;
  wire   [3:0] MCInst2_MC1_v3_2 ;
  wire   [3:0] MCInst2_MC1_v3_1 ;
  wire   [3:0] MCInst2_MC1_v3_0 ;
  wire   [3:0] MCInst2_MC1_v2_3 ;
  wire   [3:0] MCInst2_MC1_v2_2 ;
  wire   [3:0] MCInst2_MC1_v2_1 ;
  wire   [3:0] MCInst2_MC1_v2_0 ;
  wire   [3:0] MCInst2_MC1_v1_3 ;
  wire   [3:0] MCInst2_MC1_v1_2 ;
  wire   [3:0] MCInst2_MC1_v1_1 ;
  wire   [3:0] MCInst2_MC1_v1_0 ;
  wire   [3:0] MCInst2_MC1_v0_3 ;
  wire   [3:0] MCInst2_MC1_v0_2 ;
  wire   [3:0] MCInst2_MC1_v0_1 ;
  wire   [3:0] MCInst2_MC1_v0_0 ;
  wire   [3:0] MCInst2_MC2_v3_3 ;
  wire   [3:0] MCInst2_MC2_v3_2 ;
  wire   [3:0] MCInst2_MC2_v3_1 ;
  wire   [3:0] MCInst2_MC2_v3_0 ;
  wire   [3:0] MCInst2_MC2_v2_3 ;
  wire   [3:0] MCInst2_MC2_v2_2 ;
  wire   [3:0] MCInst2_MC2_v2_1 ;
  wire   [3:0] MCInst2_MC2_v2_0 ;
  wire   [3:0] MCInst2_MC2_v1_3 ;
  wire   [3:0] MCInst2_MC2_v1_2 ;
  wire   [3:0] MCInst2_MC2_v1_1 ;
  wire   [3:0] MCInst2_MC2_v1_0 ;
  wire   [3:0] MCInst2_MC2_v0_3 ;
  wire   [3:0] MCInst2_MC2_v0_2 ;
  wire   [3:0] MCInst2_MC2_v0_1 ;
  wire   [3:0] MCInst2_MC2_v0_0 ;
  wire   [3:0] MCInst2_MC3_v3_3 ;
  wire   [3:0] MCInst2_MC3_v3_2 ;
  wire   [3:0] MCInst2_MC3_v3_1 ;
  wire   [3:0] MCInst2_MC3_v3_0 ;
  wire   [3:0] MCInst2_MC3_v2_3 ;
  wire   [3:0] MCInst2_MC3_v2_2 ;
  wire   [3:0] MCInst2_MC3_v2_1 ;
  wire   [3:0] MCInst2_MC3_v2_0 ;
  wire   [3:0] MCInst2_MC3_v1_3 ;
  wire   [3:0] MCInst2_MC3_v1_2 ;
  wire   [3:0] MCInst2_MC3_v1_1 ;
  wire   [3:0] MCInst2_MC3_v1_0 ;
  wire   [3:0] MCInst2_MC3_v0_3 ;
  wire   [3:0] MCInst2_MC3_v0_2 ;
  wire   [3:0] MCInst2_MC3_v0_1 ;
  wire   [3:0] MCInst2_MC3_v0_0 ;
  wire   [3:0] MCInst3_MC0_v3_3 ;
  wire   [3:0] MCInst3_MC0_v3_2 ;
  wire   [3:0] MCInst3_MC0_v3_1 ;
  wire   [3:0] MCInst3_MC0_v3_0 ;
  wire   [3:0] MCInst3_MC0_v2_3 ;
  wire   [3:0] MCInst3_MC0_v2_2 ;
  wire   [3:0] MCInst3_MC0_v2_1 ;
  wire   [3:0] MCInst3_MC0_v2_0 ;
  wire   [3:0] MCInst3_MC0_v1_3 ;
  wire   [3:0] MCInst3_MC0_v1_2 ;
  wire   [3:0] MCInst3_MC0_v1_1 ;
  wire   [3:0] MCInst3_MC0_v1_0 ;
  wire   [3:0] MCInst3_MC0_v0_3 ;
  wire   [3:0] MCInst3_MC0_v0_2 ;
  wire   [3:0] MCInst3_MC0_v0_1 ;
  wire   [3:0] MCInst3_MC0_v0_0 ;
  wire   [3:0] MCInst3_MC1_v3_3 ;
  wire   [3:0] MCInst3_MC1_v3_2 ;
  wire   [3:0] MCInst3_MC1_v3_1 ;
  wire   [3:0] MCInst3_MC1_v3_0 ;
  wire   [3:0] MCInst3_MC1_v2_3 ;
  wire   [3:0] MCInst3_MC1_v2_2 ;
  wire   [3:0] MCInst3_MC1_v2_1 ;
  wire   [3:0] MCInst3_MC1_v2_0 ;
  wire   [3:0] MCInst3_MC1_v1_3 ;
  wire   [3:0] MCInst3_MC1_v1_2 ;
  wire   [3:0] MCInst3_MC1_v1_1 ;
  wire   [3:0] MCInst3_MC1_v1_0 ;
  wire   [3:0] MCInst3_MC1_v0_3 ;
  wire   [3:0] MCInst3_MC1_v0_2 ;
  wire   [3:0] MCInst3_MC1_v0_1 ;
  wire   [3:0] MCInst3_MC1_v0_0 ;
  wire   [3:0] MCInst3_MC2_v3_3 ;
  wire   [3:0] MCInst3_MC2_v3_2 ;
  wire   [3:0] MCInst3_MC2_v3_1 ;
  wire   [3:0] MCInst3_MC2_v3_0 ;
  wire   [3:0] MCInst3_MC2_v2_3 ;
  wire   [3:0] MCInst3_MC2_v2_2 ;
  wire   [3:0] MCInst3_MC2_v2_1 ;
  wire   [3:0] MCInst3_MC2_v2_0 ;
  wire   [3:0] MCInst3_MC2_v1_3 ;
  wire   [3:0] MCInst3_MC2_v1_2 ;
  wire   [3:0] MCInst3_MC2_v1_1 ;
  wire   [3:0] MCInst3_MC2_v1_0 ;
  wire   [3:0] MCInst3_MC2_v0_3 ;
  wire   [3:0] MCInst3_MC2_v0_2 ;
  wire   [3:0] MCInst3_MC2_v0_1 ;
  wire   [3:0] MCInst3_MC2_v0_0 ;
  wire   [3:0] MCInst3_MC3_v3_3 ;
  wire   [3:0] MCInst3_MC3_v3_2 ;
  wire   [3:0] MCInst3_MC3_v3_1 ;
  wire   [3:0] MCInst3_MC3_v3_0 ;
  wire   [3:0] MCInst3_MC3_v2_3 ;
  wire   [3:0] MCInst3_MC3_v2_2 ;
  wire   [3:0] MCInst3_MC3_v2_1 ;
  wire   [3:0] MCInst3_MC3_v2_0 ;
  wire   [3:0] MCInst3_MC3_v1_3 ;
  wire   [3:0] MCInst3_MC3_v1_2 ;
  wire   [3:0] MCInst3_MC3_v1_1 ;
  wire   [3:0] MCInst3_MC3_v1_0 ;
  wire   [3:0] MCInst3_MC3_v0_3 ;
  wire   [3:0] MCInst3_MC3_v0_2 ;
  wire   [3:0] MCInst3_MC3_v0_1 ;
  wire   [3:0] MCInst3_MC3_v0_0 ;

  INV_X1 U3 ( .A(Error[0] ), .ZN(ErrorFlag) );
  INV_X1 AddKeyXOR_XORInst_0_0_U2  ( .A(AddKeyXOR_XORInst_0_0_n2 ), .ZN(
        AddRoundKeyOutput[0]) );
  XNOR2_X1 AddKeyXOR_XORInst_0_0_U1  ( .A(Plaintext[0]), .B(Key[0]), .ZN(
        AddKeyXOR_XORInst_0_0_n2 ) );
  XOR2_X1 AddKeyXOR_XORInst_0_1_U1  ( .A(Plaintext[1]), .B(Key[1]), .Z(
        AddRoundKeyOutput[1]) );
  INV_X1 AddKeyXOR_XORInst_0_2_U2  ( .A(AddKeyXOR_XORInst_0_2_n2 ), .ZN(
        AddRoundKeyOutput[2]) );
  XNOR2_X1 AddKeyXOR_XORInst_0_2_U1  ( .A(Plaintext[2]), .B(Key[2]), .ZN(
        AddKeyXOR_XORInst_0_2_n2 ) );
  XOR2_X1 AddKeyXOR_XORInst_0_3_U1  ( .A(Plaintext[3]), .B(Key[3]), .Z(
        AddRoundKeyOutput[3]) );
  INV_X1 AddKeyXOR_XORInst_1_0_U2  ( .A(AddKeyXOR_XORInst_1_0_n2 ), .ZN(
        AddRoundKeyOutput[4]) );
  XNOR2_X1 AddKeyXOR_XORInst_1_0_U1  ( .A(Plaintext[4]), .B(Key[4]), .ZN(
        AddKeyXOR_XORInst_1_0_n2 ) );
  XOR2_X1 AddKeyXOR_XORInst_1_1_U1  ( .A(Plaintext[5]), .B(Key[5]), .Z(
        AddRoundKeyOutput[5]) );
  INV_X1 AddKeyXOR_XORInst_1_2_U2  ( .A(AddKeyXOR_XORInst_1_2_n2 ), .ZN(
        AddRoundKeyOutput[6]) );
  XNOR2_X1 AddKeyXOR_XORInst_1_2_U1  ( .A(Plaintext[6]), .B(Key[6]), .ZN(
        AddKeyXOR_XORInst_1_2_n2 ) );
  XOR2_X1 AddKeyXOR_XORInst_1_3_U1  ( .A(Plaintext[7]), .B(Key[7]), .Z(
        AddRoundKeyOutput[7]) );
  INV_X1 AddKeyXOR_XORInst_2_0_U2  ( .A(AddKeyXOR_XORInst_2_0_n2 ), .ZN(
        AddRoundKeyOutput[8]) );
  XNOR2_X1 AddKeyXOR_XORInst_2_0_U1  ( .A(Plaintext[8]), .B(Key[8]), .ZN(
        AddKeyXOR_XORInst_2_0_n2 ) );
  XOR2_X1 AddKeyXOR_XORInst_2_1_U1  ( .A(Plaintext[9]), .B(Key[9]), .Z(
        AddRoundKeyOutput[9]) );
  INV_X1 AddKeyXOR_XORInst_2_2_U2  ( .A(AddKeyXOR_XORInst_2_2_n2 ), .ZN(
        AddRoundKeyOutput[10]) );
  XNOR2_X1 AddKeyXOR_XORInst_2_2_U1  ( .A(Plaintext[10]), .B(Key[10]), .ZN(
        AddKeyXOR_XORInst_2_2_n2 ) );
  XOR2_X1 AddKeyXOR_XORInst_2_3_U1  ( .A(Plaintext[11]), .B(Key[11]), .Z(
        AddRoundKeyOutput[11]) );
  INV_X1 AddKeyXOR_XORInst_3_0_U2  ( .A(AddKeyXOR_XORInst_3_0_n2 ), .ZN(
        AddRoundKeyOutput[12]) );
  XNOR2_X1 AddKeyXOR_XORInst_3_0_U1  ( .A(Plaintext[12]), .B(Key[12]), .ZN(
        AddKeyXOR_XORInst_3_0_n2 ) );
  XOR2_X1 AddKeyXOR_XORInst_3_1_U1  ( .A(Plaintext[13]), .B(Key[13]), .Z(
        AddRoundKeyOutput[13]) );
  INV_X1 AddKeyXOR_XORInst_3_2_U2  ( .A(AddKeyXOR_XORInst_3_2_n2 ), .ZN(
        AddRoundKeyOutput[14]) );
  XNOR2_X1 AddKeyXOR_XORInst_3_2_U1  ( .A(Plaintext[14]), .B(Key[14]), .ZN(
        AddKeyXOR_XORInst_3_2_n2 ) );
  XOR2_X1 AddKeyXOR_XORInst_3_3_U1  ( .A(Plaintext[15]), .B(Key[15]), .Z(
        AddRoundKeyOutput[15]) );
  INV_X1 AddKeyXOR_XORInst_4_0_U2  ( .A(AddKeyXOR_XORInst_4_0_n2 ), .ZN(
        AddRoundKeyOutput[16]) );
  XNOR2_X1 AddKeyXOR_XORInst_4_0_U1  ( .A(Plaintext[16]), .B(Key[16]), .ZN(
        AddKeyXOR_XORInst_4_0_n2 ) );
  XOR2_X1 AddKeyXOR_XORInst_4_1_U1  ( .A(Plaintext[17]), .B(Key[17]), .Z(
        AddRoundKeyOutput[17]) );
  INV_X1 AddKeyXOR_XORInst_4_2_U2  ( .A(AddKeyXOR_XORInst_4_2_n2 ), .ZN(
        AddRoundKeyOutput[18]) );
  XNOR2_X1 AddKeyXOR_XORInst_4_2_U1  ( .A(Plaintext[18]), .B(Key[18]), .ZN(
        AddKeyXOR_XORInst_4_2_n2 ) );
  XOR2_X1 AddKeyXOR_XORInst_4_3_U1  ( .A(Plaintext[19]), .B(Key[19]), .Z(
        AddRoundKeyOutput[19]) );
  INV_X1 AddKeyXOR_XORInst_5_0_U2  ( .A(AddKeyXOR_XORInst_5_0_n2 ), .ZN(
        AddRoundKeyOutput[20]) );
  XNOR2_X1 AddKeyXOR_XORInst_5_0_U1  ( .A(Plaintext[20]), .B(Key[20]), .ZN(
        AddKeyXOR_XORInst_5_0_n2 ) );
  XOR2_X1 AddKeyXOR_XORInst_5_1_U1  ( .A(Plaintext[21]), .B(Key[21]), .Z(
        AddRoundKeyOutput[21]) );
  INV_X1 AddKeyXOR_XORInst_5_2_U2  ( .A(AddKeyXOR_XORInst_5_2_n2 ), .ZN(
        AddRoundKeyOutput[22]) );
  XNOR2_X1 AddKeyXOR_XORInst_5_2_U1  ( .A(Plaintext[22]), .B(Key[22]), .ZN(
        AddKeyXOR_XORInst_5_2_n2 ) );
  XOR2_X1 AddKeyXOR_XORInst_5_3_U1  ( .A(Plaintext[23]), .B(Key[23]), .Z(
        AddRoundKeyOutput[23]) );
  INV_X1 AddKeyXOR_XORInst_6_0_U2  ( .A(AddKeyXOR_XORInst_6_0_n2 ), .ZN(
        AddRoundKeyOutput[24]) );
  XNOR2_X1 AddKeyXOR_XORInst_6_0_U1  ( .A(Plaintext[24]), .B(Key[24]), .ZN(
        AddKeyXOR_XORInst_6_0_n2 ) );
  XOR2_X1 AddKeyXOR_XORInst_6_1_U1  ( .A(Plaintext[25]), .B(Key[25]), .Z(
        AddRoundKeyOutput[25]) );
  INV_X1 AddKeyXOR_XORInst_6_2_U2  ( .A(AddKeyXOR_XORInst_6_2_n2 ), .ZN(
        AddRoundKeyOutput[26]) );
  XNOR2_X1 AddKeyXOR_XORInst_6_2_U1  ( .A(Plaintext[26]), .B(Key[26]), .ZN(
        AddKeyXOR_XORInst_6_2_n2 ) );
  XOR2_X1 AddKeyXOR_XORInst_6_3_U1  ( .A(Plaintext[27]), .B(Key[27]), .Z(
        AddRoundKeyOutput[27]) );
  INV_X1 AddKeyXOR_XORInst_7_0_U2  ( .A(AddKeyXOR_XORInst_7_0_n2 ), .ZN(
        AddRoundKeyOutput[28]) );
  XNOR2_X1 AddKeyXOR_XORInst_7_0_U1  ( .A(Plaintext[28]), .B(Key[28]), .ZN(
        AddKeyXOR_XORInst_7_0_n2 ) );
  XOR2_X1 AddKeyXOR_XORInst_7_1_U1  ( .A(Plaintext[29]), .B(Key[29]), .Z(
        AddRoundKeyOutput[29]) );
  INV_X1 AddKeyXOR_XORInst_7_2_U2  ( .A(AddKeyXOR_XORInst_7_2_n2 ), .ZN(
        AddRoundKeyOutput[30]) );
  XNOR2_X1 AddKeyXOR_XORInst_7_2_U1  ( .A(Plaintext[30]), .B(Key[30]), .ZN(
        AddKeyXOR_XORInst_7_2_n2 ) );
  XOR2_X1 AddKeyXOR_XORInst_7_3_U1  ( .A(Plaintext[31]), .B(Key[31]), .Z(
        AddRoundKeyOutput[31]) );
  INV_X1 AddKeyXOR_XORInst_8_0_U2  ( .A(AddKeyXOR_XORInst_8_0_n2 ), .ZN(
        AddRoundKeyOutput[32]) );
  XNOR2_X1 AddKeyXOR_XORInst_8_0_U1  ( .A(Plaintext[32]), .B(Key[32]), .ZN(
        AddKeyXOR_XORInst_8_0_n2 ) );
  XOR2_X1 AddKeyXOR_XORInst_8_1_U1  ( .A(Plaintext[33]), .B(Key[33]), .Z(
        AddRoundKeyOutput[33]) );
  INV_X1 AddKeyXOR_XORInst_8_2_U2  ( .A(AddKeyXOR_XORInst_8_2_n2 ), .ZN(
        AddRoundKeyOutput[34]) );
  XNOR2_X1 AddKeyXOR_XORInst_8_2_U1  ( .A(Plaintext[34]), .B(Key[34]), .ZN(
        AddKeyXOR_XORInst_8_2_n2 ) );
  XOR2_X1 AddKeyXOR_XORInst_8_3_U1  ( .A(Plaintext[35]), .B(Key[35]), .Z(
        AddRoundKeyOutput[35]) );
  INV_X1 AddKeyXOR_XORInst_9_0_U2  ( .A(AddKeyXOR_XORInst_9_0_n2 ), .ZN(
        AddRoundKeyOutput[36]) );
  XNOR2_X1 AddKeyXOR_XORInst_9_0_U1  ( .A(Plaintext[36]), .B(Key[36]), .ZN(
        AddKeyXOR_XORInst_9_0_n2 ) );
  XOR2_X1 AddKeyXOR_XORInst_9_1_U1  ( .A(Plaintext[37]), .B(Key[37]), .Z(
        AddRoundKeyOutput[37]) );
  INV_X1 AddKeyXOR_XORInst_9_2_U2  ( .A(AddKeyXOR_XORInst_9_2_n2 ), .ZN(
        AddRoundKeyOutput[38]) );
  XNOR2_X1 AddKeyXOR_XORInst_9_2_U1  ( .A(Plaintext[38]), .B(Key[38]), .ZN(
        AddKeyXOR_XORInst_9_2_n2 ) );
  XOR2_X1 AddKeyXOR_XORInst_9_3_U1  ( .A(Plaintext[39]), .B(Key[39]), .Z(
        AddRoundKeyOutput[39]) );
  INV_X1 AddKeyXOR_XORInst_10_0_U2  ( .A(AddKeyXOR_XORInst_10_0_n2 ), .ZN(
        AddRoundKeyOutput[40]) );
  XNOR2_X1 AddKeyXOR_XORInst_10_0_U1  ( .A(Plaintext[40]), .B(Key[40]), .ZN(
        AddKeyXOR_XORInst_10_0_n2 ) );
  XOR2_X1 AddKeyXOR_XORInst_10_1_U1  ( .A(Plaintext[41]), .B(Key[41]), .Z(
        AddRoundKeyOutput[41]) );
  INV_X1 AddKeyXOR_XORInst_10_2_U2  ( .A(AddKeyXOR_XORInst_10_2_n2 ), .ZN(
        AddRoundKeyOutput[42]) );
  XNOR2_X1 AddKeyXOR_XORInst_10_2_U1  ( .A(Plaintext[42]), .B(Key[42]), .ZN(
        AddKeyXOR_XORInst_10_2_n2 ) );
  XOR2_X1 AddKeyXOR_XORInst_10_3_U1  ( .A(Plaintext[43]), .B(Key[43]), .Z(
        AddRoundKeyOutput[43]) );
  INV_X1 AddKeyXOR_XORInst_11_0_U2  ( .A(AddKeyXOR_XORInst_11_0_n2 ), .ZN(
        AddRoundKeyOutput[44]) );
  XNOR2_X1 AddKeyXOR_XORInst_11_0_U1  ( .A(Plaintext[44]), .B(Key[44]), .ZN(
        AddKeyXOR_XORInst_11_0_n2 ) );
  XOR2_X1 AddKeyXOR_XORInst_11_1_U1  ( .A(Plaintext[45]), .B(Key[45]), .Z(
        AddRoundKeyOutput[45]) );
  INV_X1 AddKeyXOR_XORInst_11_2_U2  ( .A(AddKeyXOR_XORInst_11_2_n2 ), .ZN(
        AddRoundKeyOutput[46]) );
  XNOR2_X1 AddKeyXOR_XORInst_11_2_U1  ( .A(Plaintext[46]), .B(Key[46]), .ZN(
        AddKeyXOR_XORInst_11_2_n2 ) );
  XOR2_X1 AddKeyXOR_XORInst_11_3_U1  ( .A(Plaintext[47]), .B(Key[47]), .Z(
        AddRoundKeyOutput[47]) );
  INV_X1 AddKeyXOR_XORInst_12_0_U2  ( .A(AddKeyXOR_XORInst_12_0_n2 ), .ZN(
        AddRoundKeyOutput[48]) );
  XNOR2_X1 AddKeyXOR_XORInst_12_0_U1  ( .A(Plaintext[48]), .B(Key[48]), .ZN(
        AddKeyXOR_XORInst_12_0_n2 ) );
  XOR2_X1 AddKeyXOR_XORInst_12_1_U1  ( .A(Plaintext[49]), .B(Key[49]), .Z(
        AddRoundKeyOutput[49]) );
  INV_X1 AddKeyXOR_XORInst_12_2_U2  ( .A(AddKeyXOR_XORInst_12_2_n2 ), .ZN(
        AddRoundKeyOutput[50]) );
  XNOR2_X1 AddKeyXOR_XORInst_12_2_U1  ( .A(Plaintext[50]), .B(Key[50]), .ZN(
        AddKeyXOR_XORInst_12_2_n2 ) );
  XOR2_X1 AddKeyXOR_XORInst_12_3_U1  ( .A(Plaintext[51]), .B(Key[51]), .Z(
        AddRoundKeyOutput[51]) );
  INV_X1 AddKeyXOR_XORInst_13_0_U2  ( .A(AddKeyXOR_XORInst_13_0_n2 ), .ZN(
        AddRoundKeyOutput[52]) );
  XNOR2_X1 AddKeyXOR_XORInst_13_0_U1  ( .A(Plaintext[52]), .B(Key[52]), .ZN(
        AddKeyXOR_XORInst_13_0_n2 ) );
  XOR2_X1 AddKeyXOR_XORInst_13_1_U1  ( .A(Plaintext[53]), .B(Key[53]), .Z(
        AddRoundKeyOutput[53]) );
  INV_X1 AddKeyXOR_XORInst_13_2_U2  ( .A(AddKeyXOR_XORInst_13_2_n2 ), .ZN(
        AddRoundKeyOutput[54]) );
  XNOR2_X1 AddKeyXOR_XORInst_13_2_U1  ( .A(Plaintext[54]), .B(Key[54]), .ZN(
        AddKeyXOR_XORInst_13_2_n2 ) );
  XOR2_X1 AddKeyXOR_XORInst_13_3_U1  ( .A(Plaintext[55]), .B(Key[55]), .Z(
        AddRoundKeyOutput[55]) );
  INV_X1 AddKeyXOR_XORInst_14_0_U2  ( .A(AddKeyXOR_XORInst_14_0_n2 ), .ZN(
        AddRoundKeyOutput[56]) );
  XNOR2_X1 AddKeyXOR_XORInst_14_0_U1  ( .A(Plaintext[56]), .B(Key[56]), .ZN(
        AddKeyXOR_XORInst_14_0_n2 ) );
  XOR2_X1 AddKeyXOR_XORInst_14_1_U1  ( .A(Plaintext[57]), .B(Key[57]), .Z(
        AddRoundKeyOutput[57]) );
  INV_X1 AddKeyXOR_XORInst_14_2_U2  ( .A(AddKeyXOR_XORInst_14_2_n2 ), .ZN(
        AddRoundKeyOutput[58]) );
  XNOR2_X1 AddKeyXOR_XORInst_14_2_U1  ( .A(Plaintext[58]), .B(Key[58]), .ZN(
        AddKeyXOR_XORInst_14_2_n2 ) );
  XOR2_X1 AddKeyXOR_XORInst_14_3_U1  ( .A(Plaintext[59]), .B(Key[59]), .Z(
        AddRoundKeyOutput[59]) );
  INV_X1 AddKeyXOR_XORInst_15_0_U2  ( .A(AddKeyXOR_XORInst_15_0_n2 ), .ZN(
        AddRoundKeyOutput[60]) );
  XNOR2_X1 AddKeyXOR_XORInst_15_0_U1  ( .A(Plaintext[60]), .B(Key[60]), .ZN(
        AddKeyXOR_XORInst_15_0_n2 ) );
  XOR2_X1 AddKeyXOR_XORInst_15_1_U1  ( .A(Plaintext[61]), .B(Key[61]), .Z(
        AddRoundKeyOutput[61]) );
  INV_X1 AddKeyXOR_XORInst_15_2_U2  ( .A(AddKeyXOR_XORInst_15_2_n2 ), .ZN(
        AddRoundKeyOutput[62]) );
  XNOR2_X1 AddKeyXOR_XORInst_15_2_U1  ( .A(Plaintext[62]), .B(Key[62]), .ZN(
        AddKeyXOR_XORInst_15_2_n2 ) );
  XOR2_X1 AddKeyXOR_XORInst_15_3_U1  ( .A(Plaintext[63]), .B(Key[63]), .Z(
        AddRoundKeyOutput[63]) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_0_U6  ( .A1(AddRoundKeyOutput[2]), 
        .A2(SubCellInst_LFInst_0_LFInst_0_n4 ), .ZN(
        SubCellInst_LFInst_0_LFInst_0_n5 ) );
  INV_X1 SubCellInst_LFInst_0_LFInst_0_U5  ( .A(AddRoundKeyOutput[1]), .ZN(
        SubCellInst_LFInst_0_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst_LFInst_0_LFInst_0_U4  ( .A(AddRoundKeyOutput[0]), .B(
        AddRoundKeyOutput[3]), .Z(SubCellInst_LFInst_0_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst_LFInst_0_LFInst_0_U3  ( .A(
        SubCellInst_LFInst_0_LFInst_0_n6 ), .B(
        SubCellInst_LFInst_0_LFInst_0_n5 ), .ZN(MCInst_MC0_v3_2 [3]) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_1_U12  ( .A1(
        SubCellInst_LFInst_0_LFInst_1_n18 ), .A2(
        SubCellInst_LFInst_0_LFInst_1_n17 ), .ZN(MCInst_MC0_v3_0 [2]) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_1_U11  ( .A1(AddRoundKeyOutput[1]), 
        .A2(SubCellInst_LFInst_0_LFInst_1_n16 ), .ZN(
        SubCellInst_LFInst_0_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst_LFInst_0_LFInst_1_U10  ( .A1(AddRoundKeyOutput[3]), 
        .A2(SubCellInst_LFInst_0_LFInst_1_n15 ), .ZN(
        SubCellInst_LFInst_0_LFInst_1_n16 ) );
  AND2_X1 SubCellInst_LFInst_0_LFInst_1_U9  ( .A1(AddRoundKeyOutput[0]), .A2(
        AddRoundKeyOutput[2]), .ZN(SubCellInst_LFInst_0_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_1_U8  ( .A1(AddRoundKeyOutput[3]), 
        .A2(SubCellInst_LFInst_0_LFInst_1_n14 ), .ZN(
        SubCellInst_LFInst_0_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_1_U7  ( .A1(
        SubCellInst_LFInst_0_LFInst_1_n13 ), .A2(
        SubCellInst_LFInst_0_LFInst_1_n12 ), .ZN(
        SubCellInst_LFInst_0_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_1_U6  ( .A1(AddRoundKeyOutput[0]), 
        .A2(AddRoundKeyOutput[2]), .ZN(SubCellInst_LFInst_0_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_1_U5  ( .A1(
        SubCellInst_LFInst_0_LFInst_1_n11 ), .A2(
        SubCellInst_LFInst_0_LFInst_1_n10 ), .ZN(
        SubCellInst_LFInst_0_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_1_U4  ( .A1(AddRoundKeyOutput[0]), 
        .A2(AddRoundKeyOutput[1]), .ZN(SubCellInst_LFInst_0_LFInst_1_n10 ) );
  INV_X1 SubCellInst_LFInst_0_LFInst_1_U3  ( .A(AddRoundKeyOutput[2]), .ZN(
        SubCellInst_LFInst_0_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_2_U11  ( .A1(
        SubCellInst_LFInst_0_LFInst_2_n22 ), .A2(
        SubCellInst_LFInst_0_LFInst_2_n21 ), .ZN(Red_MCInst_MC0_v3_1[0] ) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_2_U10  ( .A1(AddRoundKeyOutput[2]), 
        .A2(SubCellInst_LFInst_0_LFInst_2_n20 ), .ZN(
        SubCellInst_LFInst_0_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst_LFInst_0_LFInst_2_U9  ( .A1(AddRoundKeyOutput[1]), .A2(
        SubCellInst_LFInst_0_LFInst_2_n19 ), .ZN(
        SubCellInst_LFInst_0_LFInst_2_n20 ) );
  INV_X1 SubCellInst_LFInst_0_LFInst_2_U8  ( .A(AddRoundKeyOutput[3]), .ZN(
        SubCellInst_LFInst_0_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_2_U7  ( .A1(
        SubCellInst_LFInst_0_LFInst_2_n18 ), .A2(
        SubCellInst_LFInst_0_LFInst_2_n17 ), .ZN(
        SubCellInst_LFInst_0_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst_LFInst_0_LFInst_2_U6  ( .A(
        SubCellInst_LFInst_0_LFInst_2_n16 ), .B(AddRoundKeyOutput[2]), .Z(
        SubCellInst_LFInst_0_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_2_U5  ( .A1(AddRoundKeyOutput[0]), 
        .A2(AddRoundKeyOutput[1]), .ZN(SubCellInst_LFInst_0_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_2_U4  ( .A1(
        SubCellInst_LFInst_0_LFInst_2_n15 ), .A2(AddRoundKeyOutput[3]), .ZN(
        SubCellInst_LFInst_0_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst_LFInst_0_LFInst_2_U3  ( .A(AddRoundKeyOutput[0]), .B(
        AddRoundKeyOutput[1]), .ZN(SubCellInst_LFInst_0_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_3_U9  ( .A1(
        SubCellInst_LFInst_0_LFInst_3_n16 ), .A2(
        SubCellInst_LFInst_0_LFInst_3_n15 ), .ZN(MCInst_MC0_v3_2 [2]) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_3_U8  ( .A1(AddRoundKeyOutput[1]), 
        .A2(SubCellInst_LFInst_0_LFInst_3_n14 ), .ZN(
        SubCellInst_LFInst_0_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst_LFInst_0_LFInst_3_U7  ( .A(AddRoundKeyOutput[3]), .B(
        AddRoundKeyOutput[2]), .Z(SubCellInst_LFInst_0_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_3_U6  ( .A1(
        SubCellInst_LFInst_0_LFInst_3_n13 ), .A2(
        SubCellInst_LFInst_0_LFInst_3_n12 ), .ZN(
        SubCellInst_LFInst_0_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_3_U5  ( .A1(AddRoundKeyOutput[0]), 
        .A2(AddRoundKeyOutput[2]), .ZN(SubCellInst_LFInst_0_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst_LFInst_0_LFInst_3_U4  ( .A(AddRoundKeyOutput[0]), .B(
        SubCellInst_LFInst_0_LFInst_3_n11 ), .ZN(
        SubCellInst_LFInst_0_LFInst_3_n13 ) );
  OR2_X1 SubCellInst_LFInst_0_LFInst_3_U3  ( .A1(AddRoundKeyOutput[3]), .A2(
        AddRoundKeyOutput[1]), .ZN(SubCellInst_LFInst_0_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_0_U6  ( .A1(AddRoundKeyOutput[6]), 
        .A2(SubCellInst_LFInst_1_LFInst_0_n4 ), .ZN(
        SubCellInst_LFInst_1_LFInst_0_n5 ) );
  INV_X1 SubCellInst_LFInst_1_LFInst_0_U5  ( .A(AddRoundKeyOutput[5]), .ZN(
        SubCellInst_LFInst_1_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst_LFInst_1_LFInst_0_U4  ( .A(AddRoundKeyOutput[4]), .B(
        AddRoundKeyOutput[7]), .Z(SubCellInst_LFInst_1_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst_LFInst_1_LFInst_0_U3  ( .A(
        SubCellInst_LFInst_1_LFInst_0_n6 ), .B(
        SubCellInst_LFInst_1_LFInst_0_n5 ), .ZN(MCInst_MC3_v3_2 [3]) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_1_U12  ( .A1(
        SubCellInst_LFInst_1_LFInst_1_n18 ), .A2(
        SubCellInst_LFInst_1_LFInst_1_n17 ), .ZN(MCInst_MC3_v3_0 [2]) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_1_U11  ( .A1(AddRoundKeyOutput[5]), 
        .A2(SubCellInst_LFInst_1_LFInst_1_n16 ), .ZN(
        SubCellInst_LFInst_1_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst_LFInst_1_LFInst_1_U10  ( .A1(AddRoundKeyOutput[7]), 
        .A2(SubCellInst_LFInst_1_LFInst_1_n15 ), .ZN(
        SubCellInst_LFInst_1_LFInst_1_n16 ) );
  AND2_X1 SubCellInst_LFInst_1_LFInst_1_U9  ( .A1(AddRoundKeyOutput[4]), .A2(
        AddRoundKeyOutput[6]), .ZN(SubCellInst_LFInst_1_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_1_U8  ( .A1(AddRoundKeyOutput[7]), 
        .A2(SubCellInst_LFInst_1_LFInst_1_n14 ), .ZN(
        SubCellInst_LFInst_1_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_1_U7  ( .A1(
        SubCellInst_LFInst_1_LFInst_1_n13 ), .A2(
        SubCellInst_LFInst_1_LFInst_1_n12 ), .ZN(
        SubCellInst_LFInst_1_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_1_U6  ( .A1(AddRoundKeyOutput[4]), 
        .A2(AddRoundKeyOutput[6]), .ZN(SubCellInst_LFInst_1_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_1_U5  ( .A1(
        SubCellInst_LFInst_1_LFInst_1_n11 ), .A2(
        SubCellInst_LFInst_1_LFInst_1_n10 ), .ZN(
        SubCellInst_LFInst_1_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_1_U4  ( .A1(AddRoundKeyOutput[4]), 
        .A2(AddRoundKeyOutput[5]), .ZN(SubCellInst_LFInst_1_LFInst_1_n10 ) );
  INV_X1 SubCellInst_LFInst_1_LFInst_1_U3  ( .A(AddRoundKeyOutput[6]), .ZN(
        SubCellInst_LFInst_1_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_2_U11  ( .A1(
        SubCellInst_LFInst_1_LFInst_2_n22 ), .A2(
        SubCellInst_LFInst_1_LFInst_2_n21 ), .ZN(Red_MCInst_MC3_v3_1[0] ) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_2_U10  ( .A1(AddRoundKeyOutput[6]), 
        .A2(SubCellInst_LFInst_1_LFInst_2_n20 ), .ZN(
        SubCellInst_LFInst_1_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst_LFInst_1_LFInst_2_U9  ( .A1(AddRoundKeyOutput[5]), .A2(
        SubCellInst_LFInst_1_LFInst_2_n19 ), .ZN(
        SubCellInst_LFInst_1_LFInst_2_n20 ) );
  INV_X1 SubCellInst_LFInst_1_LFInst_2_U8  ( .A(AddRoundKeyOutput[7]), .ZN(
        SubCellInst_LFInst_1_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_2_U7  ( .A1(
        SubCellInst_LFInst_1_LFInst_2_n18 ), .A2(
        SubCellInst_LFInst_1_LFInst_2_n17 ), .ZN(
        SubCellInst_LFInst_1_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst_LFInst_1_LFInst_2_U6  ( .A(
        SubCellInst_LFInst_1_LFInst_2_n16 ), .B(AddRoundKeyOutput[6]), .Z(
        SubCellInst_LFInst_1_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_2_U5  ( .A1(AddRoundKeyOutput[4]), 
        .A2(AddRoundKeyOutput[5]), .ZN(SubCellInst_LFInst_1_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_2_U4  ( .A1(
        SubCellInst_LFInst_1_LFInst_2_n15 ), .A2(AddRoundKeyOutput[7]), .ZN(
        SubCellInst_LFInst_1_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst_LFInst_1_LFInst_2_U3  ( .A(AddRoundKeyOutput[4]), .B(
        AddRoundKeyOutput[5]), .ZN(SubCellInst_LFInst_1_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_3_U9  ( .A1(
        SubCellInst_LFInst_1_LFInst_3_n16 ), .A2(
        SubCellInst_LFInst_1_LFInst_3_n15 ), .ZN(MCInst_MC3_v3_2 [2]) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_3_U8  ( .A1(AddRoundKeyOutput[5]), 
        .A2(SubCellInst_LFInst_1_LFInst_3_n14 ), .ZN(
        SubCellInst_LFInst_1_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst_LFInst_1_LFInst_3_U7  ( .A(AddRoundKeyOutput[7]), .B(
        AddRoundKeyOutput[6]), .Z(SubCellInst_LFInst_1_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_3_U6  ( .A1(
        SubCellInst_LFInst_1_LFInst_3_n13 ), .A2(
        SubCellInst_LFInst_1_LFInst_3_n12 ), .ZN(
        SubCellInst_LFInst_1_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_3_U5  ( .A1(AddRoundKeyOutput[4]), 
        .A2(AddRoundKeyOutput[6]), .ZN(SubCellInst_LFInst_1_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst_LFInst_1_LFInst_3_U4  ( .A(AddRoundKeyOutput[4]), .B(
        SubCellInst_LFInst_1_LFInst_3_n11 ), .ZN(
        SubCellInst_LFInst_1_LFInst_3_n13 ) );
  OR2_X1 SubCellInst_LFInst_1_LFInst_3_U3  ( .A1(AddRoundKeyOutput[7]), .A2(
        AddRoundKeyOutput[5]), .ZN(SubCellInst_LFInst_1_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_0_U6  ( .A1(AddRoundKeyOutput[10]), 
        .A2(SubCellInst_LFInst_2_LFInst_0_n4 ), .ZN(
        SubCellInst_LFInst_2_LFInst_0_n5 ) );
  INV_X1 SubCellInst_LFInst_2_LFInst_0_U5  ( .A(AddRoundKeyOutput[9]), .ZN(
        SubCellInst_LFInst_2_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst_LFInst_2_LFInst_0_U4  ( .A(AddRoundKeyOutput[8]), .B(
        AddRoundKeyOutput[11]), .Z(SubCellInst_LFInst_2_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst_LFInst_2_LFInst_0_U3  ( .A(
        SubCellInst_LFInst_2_LFInst_0_n6 ), .B(
        SubCellInst_LFInst_2_LFInst_0_n5 ), .ZN(MCInst_MC2_v3_2 [3]) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_1_U12  ( .A1(
        SubCellInst_LFInst_2_LFInst_1_n18 ), .A2(
        SubCellInst_LFInst_2_LFInst_1_n17 ), .ZN(MCInst_MC2_v3_0 [2]) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_1_U11  ( .A1(AddRoundKeyOutput[9]), 
        .A2(SubCellInst_LFInst_2_LFInst_1_n16 ), .ZN(
        SubCellInst_LFInst_2_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst_LFInst_2_LFInst_1_U10  ( .A1(AddRoundKeyOutput[11]), 
        .A2(SubCellInst_LFInst_2_LFInst_1_n15 ), .ZN(
        SubCellInst_LFInst_2_LFInst_1_n16 ) );
  AND2_X1 SubCellInst_LFInst_2_LFInst_1_U9  ( .A1(AddRoundKeyOutput[8]), .A2(
        AddRoundKeyOutput[10]), .ZN(SubCellInst_LFInst_2_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_1_U8  ( .A1(AddRoundKeyOutput[11]), 
        .A2(SubCellInst_LFInst_2_LFInst_1_n14 ), .ZN(
        SubCellInst_LFInst_2_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_1_U7  ( .A1(
        SubCellInst_LFInst_2_LFInst_1_n13 ), .A2(
        SubCellInst_LFInst_2_LFInst_1_n12 ), .ZN(
        SubCellInst_LFInst_2_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_1_U6  ( .A1(AddRoundKeyOutput[8]), 
        .A2(AddRoundKeyOutput[10]), .ZN(SubCellInst_LFInst_2_LFInst_1_n12 )
         );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_1_U5  ( .A1(
        SubCellInst_LFInst_2_LFInst_1_n11 ), .A2(
        SubCellInst_LFInst_2_LFInst_1_n10 ), .ZN(
        SubCellInst_LFInst_2_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_1_U4  ( .A1(AddRoundKeyOutput[8]), 
        .A2(AddRoundKeyOutput[9]), .ZN(SubCellInst_LFInst_2_LFInst_1_n10 ) );
  INV_X1 SubCellInst_LFInst_2_LFInst_1_U3  ( .A(AddRoundKeyOutput[10]), .ZN(
        SubCellInst_LFInst_2_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_2_U11  ( .A1(
        SubCellInst_LFInst_2_LFInst_2_n22 ), .A2(
        SubCellInst_LFInst_2_LFInst_2_n21 ), .ZN(Red_MCInst_MC2_v3_1[0] ) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_2_U10  ( .A1(AddRoundKeyOutput[10]), 
        .A2(SubCellInst_LFInst_2_LFInst_2_n20 ), .ZN(
        SubCellInst_LFInst_2_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst_LFInst_2_LFInst_2_U9  ( .A1(AddRoundKeyOutput[9]), .A2(
        SubCellInst_LFInst_2_LFInst_2_n19 ), .ZN(
        SubCellInst_LFInst_2_LFInst_2_n20 ) );
  INV_X1 SubCellInst_LFInst_2_LFInst_2_U8  ( .A(AddRoundKeyOutput[11]), .ZN(
        SubCellInst_LFInst_2_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_2_U7  ( .A1(
        SubCellInst_LFInst_2_LFInst_2_n18 ), .A2(
        SubCellInst_LFInst_2_LFInst_2_n17 ), .ZN(
        SubCellInst_LFInst_2_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst_LFInst_2_LFInst_2_U6  ( .A(
        SubCellInst_LFInst_2_LFInst_2_n16 ), .B(AddRoundKeyOutput[10]), .Z(
        SubCellInst_LFInst_2_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_2_U5  ( .A1(AddRoundKeyOutput[8]), 
        .A2(AddRoundKeyOutput[9]), .ZN(SubCellInst_LFInst_2_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_2_U4  ( .A1(
        SubCellInst_LFInst_2_LFInst_2_n15 ), .A2(AddRoundKeyOutput[11]), .ZN(
        SubCellInst_LFInst_2_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst_LFInst_2_LFInst_2_U3  ( .A(AddRoundKeyOutput[8]), .B(
        AddRoundKeyOutput[9]), .ZN(SubCellInst_LFInst_2_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_3_U9  ( .A1(
        SubCellInst_LFInst_2_LFInst_3_n16 ), .A2(
        SubCellInst_LFInst_2_LFInst_3_n15 ), .ZN(MCInst_MC2_v3_2 [2]) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_3_U8  ( .A1(AddRoundKeyOutput[9]), 
        .A2(SubCellInst_LFInst_2_LFInst_3_n14 ), .ZN(
        SubCellInst_LFInst_2_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst_LFInst_2_LFInst_3_U7  ( .A(AddRoundKeyOutput[11]), .B(
        AddRoundKeyOutput[10]), .Z(SubCellInst_LFInst_2_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_3_U6  ( .A1(
        SubCellInst_LFInst_2_LFInst_3_n13 ), .A2(
        SubCellInst_LFInst_2_LFInst_3_n12 ), .ZN(
        SubCellInst_LFInst_2_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_3_U5  ( .A1(AddRoundKeyOutput[8]), 
        .A2(AddRoundKeyOutput[10]), .ZN(SubCellInst_LFInst_2_LFInst_3_n12 )
         );
  XNOR2_X1 SubCellInst_LFInst_2_LFInst_3_U4  ( .A(AddRoundKeyOutput[8]), .B(
        SubCellInst_LFInst_2_LFInst_3_n11 ), .ZN(
        SubCellInst_LFInst_2_LFInst_3_n13 ) );
  OR2_X1 SubCellInst_LFInst_2_LFInst_3_U3  ( .A1(AddRoundKeyOutput[11]), .A2(
        AddRoundKeyOutput[9]), .ZN(SubCellInst_LFInst_2_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_0_U6  ( .A1(AddRoundKeyOutput[14]), 
        .A2(SubCellInst_LFInst_3_LFInst_0_n4 ), .ZN(
        SubCellInst_LFInst_3_LFInst_0_n5 ) );
  INV_X1 SubCellInst_LFInst_3_LFInst_0_U5  ( .A(AddRoundKeyOutput[13]), .ZN(
        SubCellInst_LFInst_3_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst_LFInst_3_LFInst_0_U4  ( .A(AddRoundKeyOutput[12]), .B(
        AddRoundKeyOutput[15]), .Z(SubCellInst_LFInst_3_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst_LFInst_3_LFInst_0_U3  ( .A(
        SubCellInst_LFInst_3_LFInst_0_n6 ), .B(
        SubCellInst_LFInst_3_LFInst_0_n5 ), .ZN(MCInst_MC1_v3_2 [3]) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_1_U12  ( .A1(
        SubCellInst_LFInst_3_LFInst_1_n18 ), .A2(
        SubCellInst_LFInst_3_LFInst_1_n17 ), .ZN(MCInst_MC1_v3_0 [2]) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_1_U11  ( .A1(AddRoundKeyOutput[13]), 
        .A2(SubCellInst_LFInst_3_LFInst_1_n16 ), .ZN(
        SubCellInst_LFInst_3_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst_LFInst_3_LFInst_1_U10  ( .A1(AddRoundKeyOutput[15]), 
        .A2(SubCellInst_LFInst_3_LFInst_1_n15 ), .ZN(
        SubCellInst_LFInst_3_LFInst_1_n16 ) );
  AND2_X1 SubCellInst_LFInst_3_LFInst_1_U9  ( .A1(AddRoundKeyOutput[12]), 
        .A2(AddRoundKeyOutput[14]), .ZN(SubCellInst_LFInst_3_LFInst_1_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_1_U8  ( .A1(AddRoundKeyOutput[15]), 
        .A2(SubCellInst_LFInst_3_LFInst_1_n14 ), .ZN(
        SubCellInst_LFInst_3_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_1_U7  ( .A1(
        SubCellInst_LFInst_3_LFInst_1_n13 ), .A2(
        SubCellInst_LFInst_3_LFInst_1_n12 ), .ZN(
        SubCellInst_LFInst_3_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_1_U6  ( .A1(AddRoundKeyOutput[12]), 
        .A2(AddRoundKeyOutput[14]), .ZN(SubCellInst_LFInst_3_LFInst_1_n12 )
         );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_1_U5  ( .A1(
        SubCellInst_LFInst_3_LFInst_1_n11 ), .A2(
        SubCellInst_LFInst_3_LFInst_1_n10 ), .ZN(
        SubCellInst_LFInst_3_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_1_U4  ( .A1(AddRoundKeyOutput[12]), 
        .A2(AddRoundKeyOutput[13]), .ZN(SubCellInst_LFInst_3_LFInst_1_n10 )
         );
  INV_X1 SubCellInst_LFInst_3_LFInst_1_U3  ( .A(AddRoundKeyOutput[14]), .ZN(
        SubCellInst_LFInst_3_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_2_U11  ( .A1(
        SubCellInst_LFInst_3_LFInst_2_n22 ), .A2(
        SubCellInst_LFInst_3_LFInst_2_n21 ), .ZN(Red_MCInst_MC1_v3_1[0] ) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_2_U10  ( .A1(AddRoundKeyOutput[14]), 
        .A2(SubCellInst_LFInst_3_LFInst_2_n20 ), .ZN(
        SubCellInst_LFInst_3_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst_LFInst_3_LFInst_2_U9  ( .A1(AddRoundKeyOutput[13]), 
        .A2(SubCellInst_LFInst_3_LFInst_2_n19 ), .ZN(
        SubCellInst_LFInst_3_LFInst_2_n20 ) );
  INV_X1 SubCellInst_LFInst_3_LFInst_2_U8  ( .A(AddRoundKeyOutput[15]), .ZN(
        SubCellInst_LFInst_3_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_2_U7  ( .A1(
        SubCellInst_LFInst_3_LFInst_2_n18 ), .A2(
        SubCellInst_LFInst_3_LFInst_2_n17 ), .ZN(
        SubCellInst_LFInst_3_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst_LFInst_3_LFInst_2_U6  ( .A(
        SubCellInst_LFInst_3_LFInst_2_n16 ), .B(AddRoundKeyOutput[14]), .Z(
        SubCellInst_LFInst_3_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_2_U5  ( .A1(AddRoundKeyOutput[12]), 
        .A2(AddRoundKeyOutput[13]), .ZN(SubCellInst_LFInst_3_LFInst_2_n16 )
         );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_2_U4  ( .A1(
        SubCellInst_LFInst_3_LFInst_2_n15 ), .A2(AddRoundKeyOutput[15]), .ZN(
        SubCellInst_LFInst_3_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst_LFInst_3_LFInst_2_U3  ( .A(AddRoundKeyOutput[12]), .B(
        AddRoundKeyOutput[13]), .ZN(SubCellInst_LFInst_3_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_3_U9  ( .A1(
        SubCellInst_LFInst_3_LFInst_3_n16 ), .A2(
        SubCellInst_LFInst_3_LFInst_3_n15 ), .ZN(MCInst_MC1_v3_2 [2]) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_3_U8  ( .A1(AddRoundKeyOutput[13]), 
        .A2(SubCellInst_LFInst_3_LFInst_3_n14 ), .ZN(
        SubCellInst_LFInst_3_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst_LFInst_3_LFInst_3_U7  ( .A(AddRoundKeyOutput[15]), .B(
        AddRoundKeyOutput[14]), .Z(SubCellInst_LFInst_3_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_3_U6  ( .A1(
        SubCellInst_LFInst_3_LFInst_3_n13 ), .A2(
        SubCellInst_LFInst_3_LFInst_3_n12 ), .ZN(
        SubCellInst_LFInst_3_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_3_U5  ( .A1(AddRoundKeyOutput[12]), 
        .A2(AddRoundKeyOutput[14]), .ZN(SubCellInst_LFInst_3_LFInst_3_n12 )
         );
  XNOR2_X1 SubCellInst_LFInst_3_LFInst_3_U4  ( .A(AddRoundKeyOutput[12]), .B(
        SubCellInst_LFInst_3_LFInst_3_n11 ), .ZN(
        SubCellInst_LFInst_3_LFInst_3_n13 ) );
  OR2_X1 SubCellInst_LFInst_3_LFInst_3_U3  ( .A1(AddRoundKeyOutput[15]), .A2(
        AddRoundKeyOutput[13]), .ZN(SubCellInst_LFInst_3_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_0_U6  ( .A1(AddRoundKeyOutput[18]), 
        .A2(SubCellInst_LFInst_4_LFInst_0_n4 ), .ZN(
        SubCellInst_LFInst_4_LFInst_0_n5 ) );
  INV_X1 SubCellInst_LFInst_4_LFInst_0_U5  ( .A(AddRoundKeyOutput[17]), .ZN(
        SubCellInst_LFInst_4_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst_LFInst_4_LFInst_0_U4  ( .A(AddRoundKeyOutput[16]), .B(
        AddRoundKeyOutput[19]), .Z(SubCellInst_LFInst_4_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst_LFInst_4_LFInst_0_U3  ( .A(
        SubCellInst_LFInst_4_LFInst_0_n6 ), .B(
        SubCellInst_LFInst_4_LFInst_0_n5 ), .ZN(MCInst_MC1_v2_3 [1]) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_1_U12  ( .A1(
        SubCellInst_LFInst_4_LFInst_1_n18 ), .A2(
        SubCellInst_LFInst_4_LFInst_1_n17 ), .ZN(MCInst_MC1_v2_0 [2]) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_1_U11  ( .A1(AddRoundKeyOutput[17]), 
        .A2(SubCellInst_LFInst_4_LFInst_1_n16 ), .ZN(
        SubCellInst_LFInst_4_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst_LFInst_4_LFInst_1_U10  ( .A1(AddRoundKeyOutput[19]), 
        .A2(SubCellInst_LFInst_4_LFInst_1_n15 ), .ZN(
        SubCellInst_LFInst_4_LFInst_1_n16 ) );
  AND2_X1 SubCellInst_LFInst_4_LFInst_1_U9  ( .A1(AddRoundKeyOutput[16]), 
        .A2(AddRoundKeyOutput[18]), .ZN(SubCellInst_LFInst_4_LFInst_1_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_1_U8  ( .A1(AddRoundKeyOutput[19]), 
        .A2(SubCellInst_LFInst_4_LFInst_1_n14 ), .ZN(
        SubCellInst_LFInst_4_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_1_U7  ( .A1(
        SubCellInst_LFInst_4_LFInst_1_n13 ), .A2(
        SubCellInst_LFInst_4_LFInst_1_n12 ), .ZN(
        SubCellInst_LFInst_4_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_1_U6  ( .A1(AddRoundKeyOutput[16]), 
        .A2(AddRoundKeyOutput[18]), .ZN(SubCellInst_LFInst_4_LFInst_1_n12 )
         );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_1_U5  ( .A1(
        SubCellInst_LFInst_4_LFInst_1_n11 ), .A2(
        SubCellInst_LFInst_4_LFInst_1_n10 ), .ZN(
        SubCellInst_LFInst_4_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_1_U4  ( .A1(AddRoundKeyOutput[16]), 
        .A2(AddRoundKeyOutput[17]), .ZN(SubCellInst_LFInst_4_LFInst_1_n10 )
         );
  INV_X1 SubCellInst_LFInst_4_LFInst_1_U3  ( .A(AddRoundKeyOutput[18]), .ZN(
        SubCellInst_LFInst_4_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_2_U11  ( .A1(
        SubCellInst_LFInst_4_LFInst_2_n22 ), .A2(
        SubCellInst_LFInst_4_LFInst_2_n21 ), .ZN(MCInst_MC1_v2_0 [3]) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_2_U10  ( .A1(AddRoundKeyOutput[18]), 
        .A2(SubCellInst_LFInst_4_LFInst_2_n20 ), .ZN(
        SubCellInst_LFInst_4_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst_LFInst_4_LFInst_2_U9  ( .A1(AddRoundKeyOutput[17]), 
        .A2(SubCellInst_LFInst_4_LFInst_2_n19 ), .ZN(
        SubCellInst_LFInst_4_LFInst_2_n20 ) );
  INV_X1 SubCellInst_LFInst_4_LFInst_2_U8  ( .A(AddRoundKeyOutput[19]), .ZN(
        SubCellInst_LFInst_4_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_2_U7  ( .A1(
        SubCellInst_LFInst_4_LFInst_2_n18 ), .A2(
        SubCellInst_LFInst_4_LFInst_2_n17 ), .ZN(
        SubCellInst_LFInst_4_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst_LFInst_4_LFInst_2_U6  ( .A(
        SubCellInst_LFInst_4_LFInst_2_n16 ), .B(AddRoundKeyOutput[18]), .Z(
        SubCellInst_LFInst_4_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_2_U5  ( .A1(AddRoundKeyOutput[16]), 
        .A2(AddRoundKeyOutput[17]), .ZN(SubCellInst_LFInst_4_LFInst_2_n16 )
         );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_2_U4  ( .A1(
        SubCellInst_LFInst_4_LFInst_2_n15 ), .A2(AddRoundKeyOutput[19]), .ZN(
        SubCellInst_LFInst_4_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst_LFInst_4_LFInst_2_U3  ( .A(AddRoundKeyOutput[16]), .B(
        AddRoundKeyOutput[17]), .ZN(SubCellInst_LFInst_4_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_3_U9  ( .A1(
        SubCellInst_LFInst_4_LFInst_3_n16 ), .A2(
        SubCellInst_LFInst_4_LFInst_3_n15 ), .ZN(MCInst_MC1_v2_0 [0]) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_3_U8  ( .A1(AddRoundKeyOutput[17]), 
        .A2(SubCellInst_LFInst_4_LFInst_3_n14 ), .ZN(
        SubCellInst_LFInst_4_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst_LFInst_4_LFInst_3_U7  ( .A(AddRoundKeyOutput[19]), .B(
        AddRoundKeyOutput[18]), .Z(SubCellInst_LFInst_4_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_3_U6  ( .A1(
        SubCellInst_LFInst_4_LFInst_3_n13 ), .A2(
        SubCellInst_LFInst_4_LFInst_3_n12 ), .ZN(
        SubCellInst_LFInst_4_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_3_U5  ( .A1(AddRoundKeyOutput[16]), 
        .A2(AddRoundKeyOutput[18]), .ZN(SubCellInst_LFInst_4_LFInst_3_n12 )
         );
  XNOR2_X1 SubCellInst_LFInst_4_LFInst_3_U4  ( .A(AddRoundKeyOutput[16]), .B(
        SubCellInst_LFInst_4_LFInst_3_n11 ), .ZN(
        SubCellInst_LFInst_4_LFInst_3_n13 ) );
  OR2_X1 SubCellInst_LFInst_4_LFInst_3_U3  ( .A1(AddRoundKeyOutput[19]), .A2(
        AddRoundKeyOutput[17]), .ZN(SubCellInst_LFInst_4_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_0_U6  ( .A1(AddRoundKeyOutput[22]), 
        .A2(SubCellInst_LFInst_5_LFInst_0_n4 ), .ZN(
        SubCellInst_LFInst_5_LFInst_0_n5 ) );
  INV_X1 SubCellInst_LFInst_5_LFInst_0_U5  ( .A(AddRoundKeyOutput[21]), .ZN(
        SubCellInst_LFInst_5_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst_LFInst_5_LFInst_0_U4  ( .A(AddRoundKeyOutput[20]), .B(
        AddRoundKeyOutput[23]), .Z(SubCellInst_LFInst_5_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst_LFInst_5_LFInst_0_U3  ( .A(
        SubCellInst_LFInst_5_LFInst_0_n6 ), .B(
        SubCellInst_LFInst_5_LFInst_0_n5 ), .ZN(MCInst_MC0_v2_3 [1]) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_1_U12  ( .A1(
        SubCellInst_LFInst_5_LFInst_1_n18 ), .A2(
        SubCellInst_LFInst_5_LFInst_1_n17 ), .ZN(MCInst_MC0_v2_0 [2]) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_1_U11  ( .A1(AddRoundKeyOutput[21]), 
        .A2(SubCellInst_LFInst_5_LFInst_1_n16 ), .ZN(
        SubCellInst_LFInst_5_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst_LFInst_5_LFInst_1_U10  ( .A1(AddRoundKeyOutput[23]), 
        .A2(SubCellInst_LFInst_5_LFInst_1_n15 ), .ZN(
        SubCellInst_LFInst_5_LFInst_1_n16 ) );
  AND2_X1 SubCellInst_LFInst_5_LFInst_1_U9  ( .A1(AddRoundKeyOutput[20]), 
        .A2(AddRoundKeyOutput[22]), .ZN(SubCellInst_LFInst_5_LFInst_1_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_1_U8  ( .A1(AddRoundKeyOutput[23]), 
        .A2(SubCellInst_LFInst_5_LFInst_1_n14 ), .ZN(
        SubCellInst_LFInst_5_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_1_U7  ( .A1(
        SubCellInst_LFInst_5_LFInst_1_n13 ), .A2(
        SubCellInst_LFInst_5_LFInst_1_n12 ), .ZN(
        SubCellInst_LFInst_5_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_1_U6  ( .A1(AddRoundKeyOutput[20]), 
        .A2(AddRoundKeyOutput[22]), .ZN(SubCellInst_LFInst_5_LFInst_1_n12 )
         );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_1_U5  ( .A1(
        SubCellInst_LFInst_5_LFInst_1_n11 ), .A2(
        SubCellInst_LFInst_5_LFInst_1_n10 ), .ZN(
        SubCellInst_LFInst_5_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_1_U4  ( .A1(AddRoundKeyOutput[20]), 
        .A2(AddRoundKeyOutput[21]), .ZN(SubCellInst_LFInst_5_LFInst_1_n10 )
         );
  INV_X1 SubCellInst_LFInst_5_LFInst_1_U3  ( .A(AddRoundKeyOutput[22]), .ZN(
        SubCellInst_LFInst_5_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_2_U11  ( .A1(
        SubCellInst_LFInst_5_LFInst_2_n22 ), .A2(
        SubCellInst_LFInst_5_LFInst_2_n21 ), .ZN(MCInst_MC0_v2_0 [3]) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_2_U10  ( .A1(AddRoundKeyOutput[22]), 
        .A2(SubCellInst_LFInst_5_LFInst_2_n20 ), .ZN(
        SubCellInst_LFInst_5_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst_LFInst_5_LFInst_2_U9  ( .A1(AddRoundKeyOutput[21]), 
        .A2(SubCellInst_LFInst_5_LFInst_2_n19 ), .ZN(
        SubCellInst_LFInst_5_LFInst_2_n20 ) );
  INV_X1 SubCellInst_LFInst_5_LFInst_2_U8  ( .A(AddRoundKeyOutput[23]), .ZN(
        SubCellInst_LFInst_5_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_2_U7  ( .A1(
        SubCellInst_LFInst_5_LFInst_2_n18 ), .A2(
        SubCellInst_LFInst_5_LFInst_2_n17 ), .ZN(
        SubCellInst_LFInst_5_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst_LFInst_5_LFInst_2_U6  ( .A(
        SubCellInst_LFInst_5_LFInst_2_n16 ), .B(AddRoundKeyOutput[22]), .Z(
        SubCellInst_LFInst_5_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_2_U5  ( .A1(AddRoundKeyOutput[20]), 
        .A2(AddRoundKeyOutput[21]), .ZN(SubCellInst_LFInst_5_LFInst_2_n16 )
         );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_2_U4  ( .A1(
        SubCellInst_LFInst_5_LFInst_2_n15 ), .A2(AddRoundKeyOutput[23]), .ZN(
        SubCellInst_LFInst_5_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst_LFInst_5_LFInst_2_U3  ( .A(AddRoundKeyOutput[20]), .B(
        AddRoundKeyOutput[21]), .ZN(SubCellInst_LFInst_5_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_3_U9  ( .A1(
        SubCellInst_LFInst_5_LFInst_3_n16 ), .A2(
        SubCellInst_LFInst_5_LFInst_3_n15 ), .ZN(MCInst_MC0_v2_0 [0]) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_3_U8  ( .A1(AddRoundKeyOutput[21]), 
        .A2(SubCellInst_LFInst_5_LFInst_3_n14 ), .ZN(
        SubCellInst_LFInst_5_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst_LFInst_5_LFInst_3_U7  ( .A(AddRoundKeyOutput[23]), .B(
        AddRoundKeyOutput[22]), .Z(SubCellInst_LFInst_5_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_3_U6  ( .A1(
        SubCellInst_LFInst_5_LFInst_3_n13 ), .A2(
        SubCellInst_LFInst_5_LFInst_3_n12 ), .ZN(
        SubCellInst_LFInst_5_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_3_U5  ( .A1(AddRoundKeyOutput[20]), 
        .A2(AddRoundKeyOutput[22]), .ZN(SubCellInst_LFInst_5_LFInst_3_n12 )
         );
  XNOR2_X1 SubCellInst_LFInst_5_LFInst_3_U4  ( .A(AddRoundKeyOutput[20]), .B(
        SubCellInst_LFInst_5_LFInst_3_n11 ), .ZN(
        SubCellInst_LFInst_5_LFInst_3_n13 ) );
  OR2_X1 SubCellInst_LFInst_5_LFInst_3_U3  ( .A1(AddRoundKeyOutput[23]), .A2(
        AddRoundKeyOutput[21]), .ZN(SubCellInst_LFInst_5_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_0_U6  ( .A1(AddRoundKeyOutput[26]), 
        .A2(SubCellInst_LFInst_6_LFInst_0_n4 ), .ZN(
        SubCellInst_LFInst_6_LFInst_0_n5 ) );
  INV_X1 SubCellInst_LFInst_6_LFInst_0_U5  ( .A(AddRoundKeyOutput[25]), .ZN(
        SubCellInst_LFInst_6_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst_LFInst_6_LFInst_0_U4  ( .A(AddRoundKeyOutput[24]), .B(
        AddRoundKeyOutput[27]), .Z(SubCellInst_LFInst_6_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst_LFInst_6_LFInst_0_U3  ( .A(
        SubCellInst_LFInst_6_LFInst_0_n6 ), .B(
        SubCellInst_LFInst_6_LFInst_0_n5 ), .ZN(MCInst_MC3_v2_3 [1]) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_1_U12  ( .A1(
        SubCellInst_LFInst_6_LFInst_1_n18 ), .A2(
        SubCellInst_LFInst_6_LFInst_1_n17 ), .ZN(MCInst_MC3_v2_0 [2]) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_1_U11  ( .A1(AddRoundKeyOutput[25]), 
        .A2(SubCellInst_LFInst_6_LFInst_1_n16 ), .ZN(
        SubCellInst_LFInst_6_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst_LFInst_6_LFInst_1_U10  ( .A1(AddRoundKeyOutput[27]), 
        .A2(SubCellInst_LFInst_6_LFInst_1_n15 ), .ZN(
        SubCellInst_LFInst_6_LFInst_1_n16 ) );
  AND2_X1 SubCellInst_LFInst_6_LFInst_1_U9  ( .A1(AddRoundKeyOutput[24]), 
        .A2(AddRoundKeyOutput[26]), .ZN(SubCellInst_LFInst_6_LFInst_1_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_1_U8  ( .A1(AddRoundKeyOutput[27]), 
        .A2(SubCellInst_LFInst_6_LFInst_1_n14 ), .ZN(
        SubCellInst_LFInst_6_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_1_U7  ( .A1(
        SubCellInst_LFInst_6_LFInst_1_n13 ), .A2(
        SubCellInst_LFInst_6_LFInst_1_n12 ), .ZN(
        SubCellInst_LFInst_6_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_1_U6  ( .A1(AddRoundKeyOutput[24]), 
        .A2(AddRoundKeyOutput[26]), .ZN(SubCellInst_LFInst_6_LFInst_1_n12 )
         );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_1_U5  ( .A1(
        SubCellInst_LFInst_6_LFInst_1_n11 ), .A2(
        SubCellInst_LFInst_6_LFInst_1_n10 ), .ZN(
        SubCellInst_LFInst_6_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_1_U4  ( .A1(AddRoundKeyOutput[24]), 
        .A2(AddRoundKeyOutput[25]), .ZN(SubCellInst_LFInst_6_LFInst_1_n10 )
         );
  INV_X1 SubCellInst_LFInst_6_LFInst_1_U3  ( .A(AddRoundKeyOutput[26]), .ZN(
        SubCellInst_LFInst_6_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_2_U11  ( .A1(
        SubCellInst_LFInst_6_LFInst_2_n22 ), .A2(
        SubCellInst_LFInst_6_LFInst_2_n21 ), .ZN(MCInst_MC3_v2_0 [3]) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_2_U10  ( .A1(AddRoundKeyOutput[26]), 
        .A2(SubCellInst_LFInst_6_LFInst_2_n20 ), .ZN(
        SubCellInst_LFInst_6_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst_LFInst_6_LFInst_2_U9  ( .A1(AddRoundKeyOutput[25]), 
        .A2(SubCellInst_LFInst_6_LFInst_2_n19 ), .ZN(
        SubCellInst_LFInst_6_LFInst_2_n20 ) );
  INV_X1 SubCellInst_LFInst_6_LFInst_2_U8  ( .A(AddRoundKeyOutput[27]), .ZN(
        SubCellInst_LFInst_6_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_2_U7  ( .A1(
        SubCellInst_LFInst_6_LFInst_2_n18 ), .A2(
        SubCellInst_LFInst_6_LFInst_2_n17 ), .ZN(
        SubCellInst_LFInst_6_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst_LFInst_6_LFInst_2_U6  ( .A(
        SubCellInst_LFInst_6_LFInst_2_n16 ), .B(AddRoundKeyOutput[26]), .Z(
        SubCellInst_LFInst_6_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_2_U5  ( .A1(AddRoundKeyOutput[24]), 
        .A2(AddRoundKeyOutput[25]), .ZN(SubCellInst_LFInst_6_LFInst_2_n16 )
         );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_2_U4  ( .A1(
        SubCellInst_LFInst_6_LFInst_2_n15 ), .A2(AddRoundKeyOutput[27]), .ZN(
        SubCellInst_LFInst_6_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst_LFInst_6_LFInst_2_U3  ( .A(AddRoundKeyOutput[24]), .B(
        AddRoundKeyOutput[25]), .ZN(SubCellInst_LFInst_6_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_3_U9  ( .A1(
        SubCellInst_LFInst_6_LFInst_3_n16 ), .A2(
        SubCellInst_LFInst_6_LFInst_3_n15 ), .ZN(MCInst_MC3_v2_0 [0]) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_3_U8  ( .A1(AddRoundKeyOutput[25]), 
        .A2(SubCellInst_LFInst_6_LFInst_3_n14 ), .ZN(
        SubCellInst_LFInst_6_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst_LFInst_6_LFInst_3_U7  ( .A(AddRoundKeyOutput[27]), .B(
        AddRoundKeyOutput[26]), .Z(SubCellInst_LFInst_6_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_3_U6  ( .A1(
        SubCellInst_LFInst_6_LFInst_3_n13 ), .A2(
        SubCellInst_LFInst_6_LFInst_3_n12 ), .ZN(
        SubCellInst_LFInst_6_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_3_U5  ( .A1(AddRoundKeyOutput[24]), 
        .A2(AddRoundKeyOutput[26]), .ZN(SubCellInst_LFInst_6_LFInst_3_n12 )
         );
  XNOR2_X1 SubCellInst_LFInst_6_LFInst_3_U4  ( .A(AddRoundKeyOutput[24]), .B(
        SubCellInst_LFInst_6_LFInst_3_n11 ), .ZN(
        SubCellInst_LFInst_6_LFInst_3_n13 ) );
  OR2_X1 SubCellInst_LFInst_6_LFInst_3_U3  ( .A1(AddRoundKeyOutput[27]), .A2(
        AddRoundKeyOutput[25]), .ZN(SubCellInst_LFInst_6_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_0_U6  ( .A1(AddRoundKeyOutput[30]), 
        .A2(SubCellInst_LFInst_7_LFInst_0_n4 ), .ZN(
        SubCellInst_LFInst_7_LFInst_0_n5 ) );
  INV_X1 SubCellInst_LFInst_7_LFInst_0_U5  ( .A(AddRoundKeyOutput[29]), .ZN(
        SubCellInst_LFInst_7_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst_LFInst_7_LFInst_0_U4  ( .A(AddRoundKeyOutput[28]), .B(
        AddRoundKeyOutput[31]), .Z(SubCellInst_LFInst_7_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst_LFInst_7_LFInst_0_U3  ( .A(
        SubCellInst_LFInst_7_LFInst_0_n6 ), .B(
        SubCellInst_LFInst_7_LFInst_0_n5 ), .ZN(MCInst_MC2_v2_3 [1]) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_1_U12  ( .A1(
        SubCellInst_LFInst_7_LFInst_1_n18 ), .A2(
        SubCellInst_LFInst_7_LFInst_1_n17 ), .ZN(MCInst_MC2_v2_0 [2]) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_1_U11  ( .A1(AddRoundKeyOutput[29]), 
        .A2(SubCellInst_LFInst_7_LFInst_1_n16 ), .ZN(
        SubCellInst_LFInst_7_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst_LFInst_7_LFInst_1_U10  ( .A1(AddRoundKeyOutput[31]), 
        .A2(SubCellInst_LFInst_7_LFInst_1_n15 ), .ZN(
        SubCellInst_LFInst_7_LFInst_1_n16 ) );
  AND2_X1 SubCellInst_LFInst_7_LFInst_1_U9  ( .A1(AddRoundKeyOutput[28]), 
        .A2(AddRoundKeyOutput[30]), .ZN(SubCellInst_LFInst_7_LFInst_1_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_1_U8  ( .A1(AddRoundKeyOutput[31]), 
        .A2(SubCellInst_LFInst_7_LFInst_1_n14 ), .ZN(
        SubCellInst_LFInst_7_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_1_U7  ( .A1(
        SubCellInst_LFInst_7_LFInst_1_n13 ), .A2(
        SubCellInst_LFInst_7_LFInst_1_n12 ), .ZN(
        SubCellInst_LFInst_7_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_1_U6  ( .A1(AddRoundKeyOutput[28]), 
        .A2(AddRoundKeyOutput[30]), .ZN(SubCellInst_LFInst_7_LFInst_1_n12 )
         );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_1_U5  ( .A1(
        SubCellInst_LFInst_7_LFInst_1_n11 ), .A2(
        SubCellInst_LFInst_7_LFInst_1_n10 ), .ZN(
        SubCellInst_LFInst_7_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_1_U4  ( .A1(AddRoundKeyOutput[28]), 
        .A2(AddRoundKeyOutput[29]), .ZN(SubCellInst_LFInst_7_LFInst_1_n10 )
         );
  INV_X1 SubCellInst_LFInst_7_LFInst_1_U3  ( .A(AddRoundKeyOutput[30]), .ZN(
        SubCellInst_LFInst_7_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_2_U11  ( .A1(
        SubCellInst_LFInst_7_LFInst_2_n22 ), .A2(
        SubCellInst_LFInst_7_LFInst_2_n21 ), .ZN(MCInst_MC2_v2_0 [3]) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_2_U10  ( .A1(AddRoundKeyOutput[30]), 
        .A2(SubCellInst_LFInst_7_LFInst_2_n20 ), .ZN(
        SubCellInst_LFInst_7_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst_LFInst_7_LFInst_2_U9  ( .A1(AddRoundKeyOutput[29]), 
        .A2(SubCellInst_LFInst_7_LFInst_2_n19 ), .ZN(
        SubCellInst_LFInst_7_LFInst_2_n20 ) );
  INV_X1 SubCellInst_LFInst_7_LFInst_2_U8  ( .A(AddRoundKeyOutput[31]), .ZN(
        SubCellInst_LFInst_7_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_2_U7  ( .A1(
        SubCellInst_LFInst_7_LFInst_2_n18 ), .A2(
        SubCellInst_LFInst_7_LFInst_2_n17 ), .ZN(
        SubCellInst_LFInst_7_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst_LFInst_7_LFInst_2_U6  ( .A(
        SubCellInst_LFInst_7_LFInst_2_n16 ), .B(AddRoundKeyOutput[30]), .Z(
        SubCellInst_LFInst_7_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_2_U5  ( .A1(AddRoundKeyOutput[28]), 
        .A2(AddRoundKeyOutput[29]), .ZN(SubCellInst_LFInst_7_LFInst_2_n16 )
         );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_2_U4  ( .A1(
        SubCellInst_LFInst_7_LFInst_2_n15 ), .A2(AddRoundKeyOutput[31]), .ZN(
        SubCellInst_LFInst_7_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst_LFInst_7_LFInst_2_U3  ( .A(AddRoundKeyOutput[28]), .B(
        AddRoundKeyOutput[29]), .ZN(SubCellInst_LFInst_7_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_3_U9  ( .A1(
        SubCellInst_LFInst_7_LFInst_3_n16 ), .A2(
        SubCellInst_LFInst_7_LFInst_3_n15 ), .ZN(MCInst_MC2_v2_0 [0]) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_3_U8  ( .A1(AddRoundKeyOutput[29]), 
        .A2(SubCellInst_LFInst_7_LFInst_3_n14 ), .ZN(
        SubCellInst_LFInst_7_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst_LFInst_7_LFInst_3_U7  ( .A(AddRoundKeyOutput[31]), .B(
        AddRoundKeyOutput[30]), .Z(SubCellInst_LFInst_7_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_3_U6  ( .A1(
        SubCellInst_LFInst_7_LFInst_3_n13 ), .A2(
        SubCellInst_LFInst_7_LFInst_3_n12 ), .ZN(
        SubCellInst_LFInst_7_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_3_U5  ( .A1(AddRoundKeyOutput[28]), 
        .A2(AddRoundKeyOutput[30]), .ZN(SubCellInst_LFInst_7_LFInst_3_n12 )
         );
  XNOR2_X1 SubCellInst_LFInst_7_LFInst_3_U4  ( .A(AddRoundKeyOutput[28]), .B(
        SubCellInst_LFInst_7_LFInst_3_n11 ), .ZN(
        SubCellInst_LFInst_7_LFInst_3_n13 ) );
  OR2_X1 SubCellInst_LFInst_7_LFInst_3_U3  ( .A1(AddRoundKeyOutput[31]), .A2(
        AddRoundKeyOutput[29]), .ZN(SubCellInst_LFInst_7_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_0_U6  ( .A1(AddRoundKeyOutput[34]), 
        .A2(SubCellInst_LFInst_8_LFInst_0_n4 ), .ZN(
        SubCellInst_LFInst_8_LFInst_0_n5 ) );
  INV_X1 SubCellInst_LFInst_8_LFInst_0_U5  ( .A(AddRoundKeyOutput[33]), .ZN(
        SubCellInst_LFInst_8_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst_LFInst_8_LFInst_0_U4  ( .A(AddRoundKeyOutput[32]), .B(
        AddRoundKeyOutput[35]), .Z(SubCellInst_LFInst_8_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst_LFInst_8_LFInst_0_U3  ( .A(
        SubCellInst_LFInst_8_LFInst_0_n6 ), .B(
        SubCellInst_LFInst_8_LFInst_0_n5 ), .ZN(MCInst_MC2_v1_0 [0]) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_1_U12  ( .A1(
        SubCellInst_LFInst_8_LFInst_1_n18 ), .A2(
        SubCellInst_LFInst_8_LFInst_1_n17 ), .ZN(MCInst_MC2_v1_3 [2]) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_1_U11  ( .A1(AddRoundKeyOutput[33]), 
        .A2(SubCellInst_LFInst_8_LFInst_1_n16 ), .ZN(
        SubCellInst_LFInst_8_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst_LFInst_8_LFInst_1_U10  ( .A1(AddRoundKeyOutput[35]), 
        .A2(SubCellInst_LFInst_8_LFInst_1_n15 ), .ZN(
        SubCellInst_LFInst_8_LFInst_1_n16 ) );
  AND2_X1 SubCellInst_LFInst_8_LFInst_1_U9  ( .A1(AddRoundKeyOutput[32]), 
        .A2(AddRoundKeyOutput[34]), .ZN(SubCellInst_LFInst_8_LFInst_1_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_1_U8  ( .A1(AddRoundKeyOutput[35]), 
        .A2(SubCellInst_LFInst_8_LFInst_1_n14 ), .ZN(
        SubCellInst_LFInst_8_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_1_U7  ( .A1(
        SubCellInst_LFInst_8_LFInst_1_n13 ), .A2(
        SubCellInst_LFInst_8_LFInst_1_n12 ), .ZN(
        SubCellInst_LFInst_8_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_1_U6  ( .A1(AddRoundKeyOutput[32]), 
        .A2(AddRoundKeyOutput[34]), .ZN(SubCellInst_LFInst_8_LFInst_1_n12 )
         );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_1_U5  ( .A1(
        SubCellInst_LFInst_8_LFInst_1_n11 ), .A2(
        SubCellInst_LFInst_8_LFInst_1_n10 ), .ZN(
        SubCellInst_LFInst_8_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_1_U4  ( .A1(AddRoundKeyOutput[32]), 
        .A2(AddRoundKeyOutput[33]), .ZN(SubCellInst_LFInst_8_LFInst_1_n10 )
         );
  INV_X1 SubCellInst_LFInst_8_LFInst_1_U3  ( .A(AddRoundKeyOutput[34]), .ZN(
        SubCellInst_LFInst_8_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_2_U11  ( .A1(
        SubCellInst_LFInst_8_LFInst_2_n22 ), .A2(
        SubCellInst_LFInst_8_LFInst_2_n21 ), .ZN(Red_MCInst_MC2_v1_1[0] ) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_2_U10  ( .A1(AddRoundKeyOutput[34]), 
        .A2(SubCellInst_LFInst_8_LFInst_2_n20 ), .ZN(
        SubCellInst_LFInst_8_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst_LFInst_8_LFInst_2_U9  ( .A1(AddRoundKeyOutput[33]), 
        .A2(SubCellInst_LFInst_8_LFInst_2_n19 ), .ZN(
        SubCellInst_LFInst_8_LFInst_2_n20 ) );
  INV_X1 SubCellInst_LFInst_8_LFInst_2_U8  ( .A(AddRoundKeyOutput[35]), .ZN(
        SubCellInst_LFInst_8_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_2_U7  ( .A1(
        SubCellInst_LFInst_8_LFInst_2_n18 ), .A2(
        SubCellInst_LFInst_8_LFInst_2_n17 ), .ZN(
        SubCellInst_LFInst_8_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst_LFInst_8_LFInst_2_U6  ( .A(
        SubCellInst_LFInst_8_LFInst_2_n16 ), .B(AddRoundKeyOutput[34]), .Z(
        SubCellInst_LFInst_8_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_2_U5  ( .A1(AddRoundKeyOutput[32]), 
        .A2(AddRoundKeyOutput[33]), .ZN(SubCellInst_LFInst_8_LFInst_2_n16 )
         );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_2_U4  ( .A1(
        SubCellInst_LFInst_8_LFInst_2_n15 ), .A2(AddRoundKeyOutput[35]), .ZN(
        SubCellInst_LFInst_8_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst_LFInst_8_LFInst_2_U3  ( .A(AddRoundKeyOutput[32]), .B(
        AddRoundKeyOutput[33]), .ZN(SubCellInst_LFInst_8_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_3_U9  ( .A1(
        SubCellInst_LFInst_8_LFInst_3_n16 ), .A2(
        SubCellInst_LFInst_8_LFInst_3_n15 ), .ZN(MCInst_MC2_v1_0 [3]) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_3_U8  ( .A1(AddRoundKeyOutput[33]), 
        .A2(SubCellInst_LFInst_8_LFInst_3_n14 ), .ZN(
        SubCellInst_LFInst_8_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst_LFInst_8_LFInst_3_U7  ( .A(AddRoundKeyOutput[35]), .B(
        AddRoundKeyOutput[34]), .Z(SubCellInst_LFInst_8_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_3_U6  ( .A1(
        SubCellInst_LFInst_8_LFInst_3_n13 ), .A2(
        SubCellInst_LFInst_8_LFInst_3_n12 ), .ZN(
        SubCellInst_LFInst_8_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_3_U5  ( .A1(AddRoundKeyOutput[32]), 
        .A2(AddRoundKeyOutput[34]), .ZN(SubCellInst_LFInst_8_LFInst_3_n12 )
         );
  XNOR2_X1 SubCellInst_LFInst_8_LFInst_3_U4  ( .A(AddRoundKeyOutput[32]), .B(
        SubCellInst_LFInst_8_LFInst_3_n11 ), .ZN(
        SubCellInst_LFInst_8_LFInst_3_n13 ) );
  OR2_X1 SubCellInst_LFInst_8_LFInst_3_U3  ( .A1(AddRoundKeyOutput[35]), .A2(
        AddRoundKeyOutput[33]), .ZN(SubCellInst_LFInst_8_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_0_U6  ( .A1(AddRoundKeyOutput[38]), 
        .A2(SubCellInst_LFInst_9_LFInst_0_n4 ), .ZN(
        SubCellInst_LFInst_9_LFInst_0_n5 ) );
  INV_X1 SubCellInst_LFInst_9_LFInst_0_U5  ( .A(AddRoundKeyOutput[37]), .ZN(
        SubCellInst_LFInst_9_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst_LFInst_9_LFInst_0_U4  ( .A(AddRoundKeyOutput[36]), .B(
        AddRoundKeyOutput[39]), .Z(SubCellInst_LFInst_9_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst_LFInst_9_LFInst_0_U3  ( .A(
        SubCellInst_LFInst_9_LFInst_0_n6 ), .B(
        SubCellInst_LFInst_9_LFInst_0_n5 ), .ZN(MCInst_MC1_v1_0 [0]) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_1_U12  ( .A1(
        SubCellInst_LFInst_9_LFInst_1_n18 ), .A2(
        SubCellInst_LFInst_9_LFInst_1_n17 ), .ZN(MCInst_MC1_v1_3 [2]) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_1_U11  ( .A1(AddRoundKeyOutput[37]), 
        .A2(SubCellInst_LFInst_9_LFInst_1_n16 ), .ZN(
        SubCellInst_LFInst_9_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst_LFInst_9_LFInst_1_U10  ( .A1(AddRoundKeyOutput[39]), 
        .A2(SubCellInst_LFInst_9_LFInst_1_n15 ), .ZN(
        SubCellInst_LFInst_9_LFInst_1_n16 ) );
  AND2_X1 SubCellInst_LFInst_9_LFInst_1_U9  ( .A1(AddRoundKeyOutput[36]), 
        .A2(AddRoundKeyOutput[38]), .ZN(SubCellInst_LFInst_9_LFInst_1_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_1_U8  ( .A1(AddRoundKeyOutput[39]), 
        .A2(SubCellInst_LFInst_9_LFInst_1_n14 ), .ZN(
        SubCellInst_LFInst_9_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_1_U7  ( .A1(
        SubCellInst_LFInst_9_LFInst_1_n13 ), .A2(
        SubCellInst_LFInst_9_LFInst_1_n12 ), .ZN(
        SubCellInst_LFInst_9_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_1_U6  ( .A1(AddRoundKeyOutput[36]), 
        .A2(AddRoundKeyOutput[38]), .ZN(SubCellInst_LFInst_9_LFInst_1_n12 )
         );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_1_U5  ( .A1(
        SubCellInst_LFInst_9_LFInst_1_n11 ), .A2(
        SubCellInst_LFInst_9_LFInst_1_n10 ), .ZN(
        SubCellInst_LFInst_9_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_1_U4  ( .A1(AddRoundKeyOutput[36]), 
        .A2(AddRoundKeyOutput[37]), .ZN(SubCellInst_LFInst_9_LFInst_1_n10 )
         );
  INV_X1 SubCellInst_LFInst_9_LFInst_1_U3  ( .A(AddRoundKeyOutput[38]), .ZN(
        SubCellInst_LFInst_9_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_2_U11  ( .A1(
        SubCellInst_LFInst_9_LFInst_2_n22 ), .A2(
        SubCellInst_LFInst_9_LFInst_2_n21 ), .ZN(Red_MCInst_MC1_v1_1[0] ) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_2_U10  ( .A1(AddRoundKeyOutput[38]), 
        .A2(SubCellInst_LFInst_9_LFInst_2_n20 ), .ZN(
        SubCellInst_LFInst_9_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst_LFInst_9_LFInst_2_U9  ( .A1(AddRoundKeyOutput[37]), 
        .A2(SubCellInst_LFInst_9_LFInst_2_n19 ), .ZN(
        SubCellInst_LFInst_9_LFInst_2_n20 ) );
  INV_X1 SubCellInst_LFInst_9_LFInst_2_U8  ( .A(AddRoundKeyOutput[39]), .ZN(
        SubCellInst_LFInst_9_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_2_U7  ( .A1(
        SubCellInst_LFInst_9_LFInst_2_n18 ), .A2(
        SubCellInst_LFInst_9_LFInst_2_n17 ), .ZN(
        SubCellInst_LFInst_9_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst_LFInst_9_LFInst_2_U6  ( .A(
        SubCellInst_LFInst_9_LFInst_2_n16 ), .B(AddRoundKeyOutput[38]), .Z(
        SubCellInst_LFInst_9_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_2_U5  ( .A1(AddRoundKeyOutput[36]), 
        .A2(AddRoundKeyOutput[37]), .ZN(SubCellInst_LFInst_9_LFInst_2_n16 )
         );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_2_U4  ( .A1(
        SubCellInst_LFInst_9_LFInst_2_n15 ), .A2(AddRoundKeyOutput[39]), .ZN(
        SubCellInst_LFInst_9_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst_LFInst_9_LFInst_2_U3  ( .A(AddRoundKeyOutput[36]), .B(
        AddRoundKeyOutput[37]), .ZN(SubCellInst_LFInst_9_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_3_U9  ( .A1(
        SubCellInst_LFInst_9_LFInst_3_n16 ), .A2(
        SubCellInst_LFInst_9_LFInst_3_n15 ), .ZN(MCInst_MC1_v1_0 [3]) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_3_U8  ( .A1(AddRoundKeyOutput[37]), 
        .A2(SubCellInst_LFInst_9_LFInst_3_n14 ), .ZN(
        SubCellInst_LFInst_9_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst_LFInst_9_LFInst_3_U7  ( .A(AddRoundKeyOutput[39]), .B(
        AddRoundKeyOutput[38]), .Z(SubCellInst_LFInst_9_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_3_U6  ( .A1(
        SubCellInst_LFInst_9_LFInst_3_n13 ), .A2(
        SubCellInst_LFInst_9_LFInst_3_n12 ), .ZN(
        SubCellInst_LFInst_9_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_3_U5  ( .A1(AddRoundKeyOutput[36]), 
        .A2(AddRoundKeyOutput[38]), .ZN(SubCellInst_LFInst_9_LFInst_3_n12 )
         );
  XNOR2_X1 SubCellInst_LFInst_9_LFInst_3_U4  ( .A(AddRoundKeyOutput[36]), .B(
        SubCellInst_LFInst_9_LFInst_3_n11 ), .ZN(
        SubCellInst_LFInst_9_LFInst_3_n13 ) );
  OR2_X1 SubCellInst_LFInst_9_LFInst_3_U3  ( .A1(AddRoundKeyOutput[39]), .A2(
        AddRoundKeyOutput[37]), .ZN(SubCellInst_LFInst_9_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_0_U6  ( .A1(AddRoundKeyOutput[42]), 
        .A2(SubCellInst_LFInst_10_LFInst_0_n4 ), .ZN(
        SubCellInst_LFInst_10_LFInst_0_n5 ) );
  INV_X1 SubCellInst_LFInst_10_LFInst_0_U5  ( .A(AddRoundKeyOutput[41]), .ZN(
        SubCellInst_LFInst_10_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst_LFInst_10_LFInst_0_U4  ( .A(AddRoundKeyOutput[40]), .B(
        AddRoundKeyOutput[43]), .Z(SubCellInst_LFInst_10_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst_LFInst_10_LFInst_0_U3  ( .A(
        SubCellInst_LFInst_10_LFInst_0_n6 ), .B(
        SubCellInst_LFInst_10_LFInst_0_n5 ), .ZN(MCInst_MC0_v1_0 [0]) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_1_U12  ( .A1(
        SubCellInst_LFInst_10_LFInst_1_n18 ), .A2(
        SubCellInst_LFInst_10_LFInst_1_n17 ), .ZN(MCInst_MC0_v1_3 [2]) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_1_U11  ( .A1(AddRoundKeyOutput[41]), 
        .A2(SubCellInst_LFInst_10_LFInst_1_n16 ), .ZN(
        SubCellInst_LFInst_10_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst_LFInst_10_LFInst_1_U10  ( .A1(AddRoundKeyOutput[43]), 
        .A2(SubCellInst_LFInst_10_LFInst_1_n15 ), .ZN(
        SubCellInst_LFInst_10_LFInst_1_n16 ) );
  AND2_X1 SubCellInst_LFInst_10_LFInst_1_U9  ( .A1(AddRoundKeyOutput[40]), 
        .A2(AddRoundKeyOutput[42]), .ZN(SubCellInst_LFInst_10_LFInst_1_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_1_U8  ( .A1(AddRoundKeyOutput[43]), 
        .A2(SubCellInst_LFInst_10_LFInst_1_n14 ), .ZN(
        SubCellInst_LFInst_10_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_1_U7  ( .A1(
        SubCellInst_LFInst_10_LFInst_1_n13 ), .A2(
        SubCellInst_LFInst_10_LFInst_1_n12 ), .ZN(
        SubCellInst_LFInst_10_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_1_U6  ( .A1(AddRoundKeyOutput[40]), 
        .A2(AddRoundKeyOutput[42]), .ZN(SubCellInst_LFInst_10_LFInst_1_n12 )
         );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_1_U5  ( .A1(
        SubCellInst_LFInst_10_LFInst_1_n11 ), .A2(
        SubCellInst_LFInst_10_LFInst_1_n10 ), .ZN(
        SubCellInst_LFInst_10_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_1_U4  ( .A1(AddRoundKeyOutput[40]), 
        .A2(AddRoundKeyOutput[41]), .ZN(SubCellInst_LFInst_10_LFInst_1_n10 )
         );
  INV_X1 SubCellInst_LFInst_10_LFInst_1_U3  ( .A(AddRoundKeyOutput[42]), .ZN(
        SubCellInst_LFInst_10_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_2_U11  ( .A1(
        SubCellInst_LFInst_10_LFInst_2_n22 ), .A2(
        SubCellInst_LFInst_10_LFInst_2_n21 ), .ZN(Red_MCInst_MC0_v1_1[0] )
         );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_2_U10  ( .A1(AddRoundKeyOutput[42]), 
        .A2(SubCellInst_LFInst_10_LFInst_2_n20 ), .ZN(
        SubCellInst_LFInst_10_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst_LFInst_10_LFInst_2_U9  ( .A1(AddRoundKeyOutput[41]), 
        .A2(SubCellInst_LFInst_10_LFInst_2_n19 ), .ZN(
        SubCellInst_LFInst_10_LFInst_2_n20 ) );
  INV_X1 SubCellInst_LFInst_10_LFInst_2_U8  ( .A(AddRoundKeyOutput[43]), .ZN(
        SubCellInst_LFInst_10_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_2_U7  ( .A1(
        SubCellInst_LFInst_10_LFInst_2_n18 ), .A2(
        SubCellInst_LFInst_10_LFInst_2_n17 ), .ZN(
        SubCellInst_LFInst_10_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst_LFInst_10_LFInst_2_U6  ( .A(
        SubCellInst_LFInst_10_LFInst_2_n16 ), .B(AddRoundKeyOutput[42]), .Z(
        SubCellInst_LFInst_10_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_2_U5  ( .A1(AddRoundKeyOutput[40]), 
        .A2(AddRoundKeyOutput[41]), .ZN(SubCellInst_LFInst_10_LFInst_2_n16 )
         );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_2_U4  ( .A1(
        SubCellInst_LFInst_10_LFInst_2_n15 ), .A2(AddRoundKeyOutput[43]), 
        .ZN(SubCellInst_LFInst_10_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst_LFInst_10_LFInst_2_U3  ( .A(AddRoundKeyOutput[40]), 
        .B(AddRoundKeyOutput[41]), .ZN(SubCellInst_LFInst_10_LFInst_2_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_3_U9  ( .A1(
        SubCellInst_LFInst_10_LFInst_3_n16 ), .A2(
        SubCellInst_LFInst_10_LFInst_3_n15 ), .ZN(MCInst_MC0_v1_0 [3]) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_3_U8  ( .A1(AddRoundKeyOutput[41]), 
        .A2(SubCellInst_LFInst_10_LFInst_3_n14 ), .ZN(
        SubCellInst_LFInst_10_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst_LFInst_10_LFInst_3_U7  ( .A(AddRoundKeyOutput[43]), .B(
        AddRoundKeyOutput[42]), .Z(SubCellInst_LFInst_10_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_3_U6  ( .A1(
        SubCellInst_LFInst_10_LFInst_3_n13 ), .A2(
        SubCellInst_LFInst_10_LFInst_3_n12 ), .ZN(
        SubCellInst_LFInst_10_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_3_U5  ( .A1(AddRoundKeyOutput[40]), 
        .A2(AddRoundKeyOutput[42]), .ZN(SubCellInst_LFInst_10_LFInst_3_n12 )
         );
  XNOR2_X1 SubCellInst_LFInst_10_LFInst_3_U4  ( .A(AddRoundKeyOutput[40]), 
        .B(SubCellInst_LFInst_10_LFInst_3_n11 ), .ZN(
        SubCellInst_LFInst_10_LFInst_3_n13 ) );
  OR2_X1 SubCellInst_LFInst_10_LFInst_3_U3  ( .A1(AddRoundKeyOutput[43]), 
        .A2(AddRoundKeyOutput[41]), .ZN(SubCellInst_LFInst_10_LFInst_3_n11 )
         );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_0_U6  ( .A1(AddRoundKeyOutput[46]), 
        .A2(SubCellInst_LFInst_11_LFInst_0_n4 ), .ZN(
        SubCellInst_LFInst_11_LFInst_0_n5 ) );
  INV_X1 SubCellInst_LFInst_11_LFInst_0_U5  ( .A(AddRoundKeyOutput[45]), .ZN(
        SubCellInst_LFInst_11_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst_LFInst_11_LFInst_0_U4  ( .A(AddRoundKeyOutput[44]), .B(
        AddRoundKeyOutput[47]), .Z(SubCellInst_LFInst_11_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst_LFInst_11_LFInst_0_U3  ( .A(
        SubCellInst_LFInst_11_LFInst_0_n6 ), .B(
        SubCellInst_LFInst_11_LFInst_0_n5 ), .ZN(MCInst_MC3_v1_0 [0]) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_1_U12  ( .A1(
        SubCellInst_LFInst_11_LFInst_1_n18 ), .A2(
        SubCellInst_LFInst_11_LFInst_1_n17 ), .ZN(MCInst_MC3_v1_3 [2]) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_1_U11  ( .A1(AddRoundKeyOutput[45]), 
        .A2(SubCellInst_LFInst_11_LFInst_1_n16 ), .ZN(
        SubCellInst_LFInst_11_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst_LFInst_11_LFInst_1_U10  ( .A1(AddRoundKeyOutput[47]), 
        .A2(SubCellInst_LFInst_11_LFInst_1_n15 ), .ZN(
        SubCellInst_LFInst_11_LFInst_1_n16 ) );
  AND2_X1 SubCellInst_LFInst_11_LFInst_1_U9  ( .A1(AddRoundKeyOutput[44]), 
        .A2(AddRoundKeyOutput[46]), .ZN(SubCellInst_LFInst_11_LFInst_1_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_1_U8  ( .A1(AddRoundKeyOutput[47]), 
        .A2(SubCellInst_LFInst_11_LFInst_1_n14 ), .ZN(
        SubCellInst_LFInst_11_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_1_U7  ( .A1(
        SubCellInst_LFInst_11_LFInst_1_n13 ), .A2(
        SubCellInst_LFInst_11_LFInst_1_n12 ), .ZN(
        SubCellInst_LFInst_11_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_1_U6  ( .A1(AddRoundKeyOutput[44]), 
        .A2(AddRoundKeyOutput[46]), .ZN(SubCellInst_LFInst_11_LFInst_1_n12 )
         );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_1_U5  ( .A1(
        SubCellInst_LFInst_11_LFInst_1_n11 ), .A2(
        SubCellInst_LFInst_11_LFInst_1_n10 ), .ZN(
        SubCellInst_LFInst_11_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_1_U4  ( .A1(AddRoundKeyOutput[44]), 
        .A2(AddRoundKeyOutput[45]), .ZN(SubCellInst_LFInst_11_LFInst_1_n10 )
         );
  INV_X1 SubCellInst_LFInst_11_LFInst_1_U3  ( .A(AddRoundKeyOutput[46]), .ZN(
        SubCellInst_LFInst_11_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_2_U11  ( .A1(
        SubCellInst_LFInst_11_LFInst_2_n22 ), .A2(
        SubCellInst_LFInst_11_LFInst_2_n21 ), .ZN(Red_MCInst_MC3_v1_1[0] )
         );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_2_U10  ( .A1(AddRoundKeyOutput[46]), 
        .A2(SubCellInst_LFInst_11_LFInst_2_n20 ), .ZN(
        SubCellInst_LFInst_11_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst_LFInst_11_LFInst_2_U9  ( .A1(AddRoundKeyOutput[45]), 
        .A2(SubCellInst_LFInst_11_LFInst_2_n19 ), .ZN(
        SubCellInst_LFInst_11_LFInst_2_n20 ) );
  INV_X1 SubCellInst_LFInst_11_LFInst_2_U8  ( .A(AddRoundKeyOutput[47]), .ZN(
        SubCellInst_LFInst_11_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_2_U7  ( .A1(
        SubCellInst_LFInst_11_LFInst_2_n18 ), .A2(
        SubCellInst_LFInst_11_LFInst_2_n17 ), .ZN(
        SubCellInst_LFInst_11_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst_LFInst_11_LFInst_2_U6  ( .A(
        SubCellInst_LFInst_11_LFInst_2_n16 ), .B(AddRoundKeyOutput[46]), .Z(
        SubCellInst_LFInst_11_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_2_U5  ( .A1(AddRoundKeyOutput[44]), 
        .A2(AddRoundKeyOutput[45]), .ZN(SubCellInst_LFInst_11_LFInst_2_n16 )
         );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_2_U4  ( .A1(
        SubCellInst_LFInst_11_LFInst_2_n15 ), .A2(AddRoundKeyOutput[47]), 
        .ZN(SubCellInst_LFInst_11_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst_LFInst_11_LFInst_2_U3  ( .A(AddRoundKeyOutput[44]), 
        .B(AddRoundKeyOutput[45]), .ZN(SubCellInst_LFInst_11_LFInst_2_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_3_U9  ( .A1(
        SubCellInst_LFInst_11_LFInst_3_n16 ), .A2(
        SubCellInst_LFInst_11_LFInst_3_n15 ), .ZN(MCInst_MC3_v1_0 [3]) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_3_U8  ( .A1(AddRoundKeyOutput[45]), 
        .A2(SubCellInst_LFInst_11_LFInst_3_n14 ), .ZN(
        SubCellInst_LFInst_11_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst_LFInst_11_LFInst_3_U7  ( .A(AddRoundKeyOutput[47]), .B(
        AddRoundKeyOutput[46]), .Z(SubCellInst_LFInst_11_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_3_U6  ( .A1(
        SubCellInst_LFInst_11_LFInst_3_n13 ), .A2(
        SubCellInst_LFInst_11_LFInst_3_n12 ), .ZN(
        SubCellInst_LFInst_11_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_3_U5  ( .A1(AddRoundKeyOutput[44]), 
        .A2(AddRoundKeyOutput[46]), .ZN(SubCellInst_LFInst_11_LFInst_3_n12 )
         );
  XNOR2_X1 SubCellInst_LFInst_11_LFInst_3_U4  ( .A(AddRoundKeyOutput[44]), 
        .B(SubCellInst_LFInst_11_LFInst_3_n11 ), .ZN(
        SubCellInst_LFInst_11_LFInst_3_n13 ) );
  OR2_X1 SubCellInst_LFInst_11_LFInst_3_U3  ( .A1(AddRoundKeyOutput[47]), 
        .A2(AddRoundKeyOutput[45]), .ZN(SubCellInst_LFInst_11_LFInst_3_n11 )
         );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_0_U6  ( .A1(AddRoundKeyOutput[50]), 
        .A2(SubCellInst_LFInst_12_LFInst_0_n4 ), .ZN(
        SubCellInst_LFInst_12_LFInst_0_n5 ) );
  INV_X1 SubCellInst_LFInst_12_LFInst_0_U5  ( .A(AddRoundKeyOutput[49]), .ZN(
        SubCellInst_LFInst_12_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst_LFInst_12_LFInst_0_U4  ( .A(AddRoundKeyOutput[48]), .B(
        AddRoundKeyOutput[51]), .Z(SubCellInst_LFInst_12_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst_LFInst_12_LFInst_0_U3  ( .A(
        SubCellInst_LFInst_12_LFInst_0_n6 ), .B(
        SubCellInst_LFInst_12_LFInst_0_n5 ), .ZN(Red_MCInst_MC3_v0_1[0] ) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_1_U12  ( .A1(
        SubCellInst_LFInst_12_LFInst_1_n18 ), .A2(
        SubCellInst_LFInst_12_LFInst_1_n17 ), .ZN(MCInst_MC3_v0_0 [3]) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_1_U11  ( .A1(AddRoundKeyOutput[49]), 
        .A2(SubCellInst_LFInst_12_LFInst_1_n16 ), .ZN(
        SubCellInst_LFInst_12_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst_LFInst_12_LFInst_1_U10  ( .A1(AddRoundKeyOutput[51]), 
        .A2(SubCellInst_LFInst_12_LFInst_1_n15 ), .ZN(
        SubCellInst_LFInst_12_LFInst_1_n16 ) );
  AND2_X1 SubCellInst_LFInst_12_LFInst_1_U9  ( .A1(AddRoundKeyOutput[48]), 
        .A2(AddRoundKeyOutput[50]), .ZN(SubCellInst_LFInst_12_LFInst_1_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_1_U8  ( .A1(AddRoundKeyOutput[51]), 
        .A2(SubCellInst_LFInst_12_LFInst_1_n14 ), .ZN(
        SubCellInst_LFInst_12_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_1_U7  ( .A1(
        SubCellInst_LFInst_12_LFInst_1_n13 ), .A2(
        SubCellInst_LFInst_12_LFInst_1_n12 ), .ZN(
        SubCellInst_LFInst_12_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_1_U6  ( .A1(AddRoundKeyOutput[48]), 
        .A2(AddRoundKeyOutput[50]), .ZN(SubCellInst_LFInst_12_LFInst_1_n12 )
         );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_1_U5  ( .A1(
        SubCellInst_LFInst_12_LFInst_1_n11 ), .A2(
        SubCellInst_LFInst_12_LFInst_1_n10 ), .ZN(
        SubCellInst_LFInst_12_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_1_U4  ( .A1(AddRoundKeyOutput[48]), 
        .A2(AddRoundKeyOutput[49]), .ZN(SubCellInst_LFInst_12_LFInst_1_n10 )
         );
  INV_X1 SubCellInst_LFInst_12_LFInst_1_U3  ( .A(AddRoundKeyOutput[50]), .ZN(
        SubCellInst_LFInst_12_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_2_U11  ( .A1(
        SubCellInst_LFInst_12_LFInst_2_n22 ), .A2(
        SubCellInst_LFInst_12_LFInst_2_n21 ), .ZN(MCInst_MC3_v0_3 [3]) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_2_U10  ( .A1(AddRoundKeyOutput[50]), 
        .A2(SubCellInst_LFInst_12_LFInst_2_n20 ), .ZN(
        SubCellInst_LFInst_12_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst_LFInst_12_LFInst_2_U9  ( .A1(AddRoundKeyOutput[49]), 
        .A2(SubCellInst_LFInst_12_LFInst_2_n19 ), .ZN(
        SubCellInst_LFInst_12_LFInst_2_n20 ) );
  INV_X1 SubCellInst_LFInst_12_LFInst_2_U8  ( .A(AddRoundKeyOutput[51]), .ZN(
        SubCellInst_LFInst_12_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_2_U7  ( .A1(
        SubCellInst_LFInst_12_LFInst_2_n18 ), .A2(
        SubCellInst_LFInst_12_LFInst_2_n17 ), .ZN(
        SubCellInst_LFInst_12_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst_LFInst_12_LFInst_2_U6  ( .A(
        SubCellInst_LFInst_12_LFInst_2_n16 ), .B(AddRoundKeyOutput[50]), .Z(
        SubCellInst_LFInst_12_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_2_U5  ( .A1(AddRoundKeyOutput[48]), 
        .A2(AddRoundKeyOutput[49]), .ZN(SubCellInst_LFInst_12_LFInst_2_n16 )
         );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_2_U4  ( .A1(
        SubCellInst_LFInst_12_LFInst_2_n15 ), .A2(AddRoundKeyOutput[51]), 
        .ZN(SubCellInst_LFInst_12_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst_LFInst_12_LFInst_2_U3  ( .A(AddRoundKeyOutput[48]), 
        .B(AddRoundKeyOutput[49]), .ZN(SubCellInst_LFInst_12_LFInst_2_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_3_U9  ( .A1(
        SubCellInst_LFInst_12_LFInst_3_n16 ), .A2(
        SubCellInst_LFInst_12_LFInst_3_n15 ), .ZN(MCInst_MC3_v0_3 [0]) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_3_U8  ( .A1(AddRoundKeyOutput[49]), 
        .A2(SubCellInst_LFInst_12_LFInst_3_n14 ), .ZN(
        SubCellInst_LFInst_12_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst_LFInst_12_LFInst_3_U7  ( .A(AddRoundKeyOutput[51]), .B(
        AddRoundKeyOutput[50]), .Z(SubCellInst_LFInst_12_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_3_U6  ( .A1(
        SubCellInst_LFInst_12_LFInst_3_n13 ), .A2(
        SubCellInst_LFInst_12_LFInst_3_n12 ), .ZN(
        SubCellInst_LFInst_12_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_3_U5  ( .A1(AddRoundKeyOutput[48]), 
        .A2(AddRoundKeyOutput[50]), .ZN(SubCellInst_LFInst_12_LFInst_3_n12 )
         );
  XNOR2_X1 SubCellInst_LFInst_12_LFInst_3_U4  ( .A(AddRoundKeyOutput[48]), 
        .B(SubCellInst_LFInst_12_LFInst_3_n11 ), .ZN(
        SubCellInst_LFInst_12_LFInst_3_n13 ) );
  OR2_X1 SubCellInst_LFInst_12_LFInst_3_U3  ( .A1(AddRoundKeyOutput[51]), 
        .A2(AddRoundKeyOutput[49]), .ZN(SubCellInst_LFInst_12_LFInst_3_n11 )
         );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_0_U6  ( .A1(AddRoundKeyOutput[54]), 
        .A2(SubCellInst_LFInst_13_LFInst_0_n4 ), .ZN(
        SubCellInst_LFInst_13_LFInst_0_n5 ) );
  INV_X1 SubCellInst_LFInst_13_LFInst_0_U5  ( .A(AddRoundKeyOutput[53]), .ZN(
        SubCellInst_LFInst_13_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst_LFInst_13_LFInst_0_U4  ( .A(AddRoundKeyOutput[52]), .B(
        AddRoundKeyOutput[55]), .Z(SubCellInst_LFInst_13_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst_LFInst_13_LFInst_0_U3  ( .A(
        SubCellInst_LFInst_13_LFInst_0_n6 ), .B(
        SubCellInst_LFInst_13_LFInst_0_n5 ), .ZN(Red_MCInst_MC2_v0_1[0] ) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_1_U12  ( .A1(
        SubCellInst_LFInst_13_LFInst_1_n18 ), .A2(
        SubCellInst_LFInst_13_LFInst_1_n17 ), .ZN(MCInst_MC2_v0_0 [3]) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_1_U11  ( .A1(AddRoundKeyOutput[53]), 
        .A2(SubCellInst_LFInst_13_LFInst_1_n16 ), .ZN(
        SubCellInst_LFInst_13_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst_LFInst_13_LFInst_1_U10  ( .A1(AddRoundKeyOutput[55]), 
        .A2(SubCellInst_LFInst_13_LFInst_1_n15 ), .ZN(
        SubCellInst_LFInst_13_LFInst_1_n16 ) );
  AND2_X1 SubCellInst_LFInst_13_LFInst_1_U9  ( .A1(AddRoundKeyOutput[52]), 
        .A2(AddRoundKeyOutput[54]), .ZN(SubCellInst_LFInst_13_LFInst_1_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_1_U8  ( .A1(AddRoundKeyOutput[55]), 
        .A2(SubCellInst_LFInst_13_LFInst_1_n14 ), .ZN(
        SubCellInst_LFInst_13_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_1_U7  ( .A1(
        SubCellInst_LFInst_13_LFInst_1_n13 ), .A2(
        SubCellInst_LFInst_13_LFInst_1_n12 ), .ZN(
        SubCellInst_LFInst_13_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_1_U6  ( .A1(AddRoundKeyOutput[52]), 
        .A2(AddRoundKeyOutput[54]), .ZN(SubCellInst_LFInst_13_LFInst_1_n12 )
         );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_1_U5  ( .A1(
        SubCellInst_LFInst_13_LFInst_1_n11 ), .A2(
        SubCellInst_LFInst_13_LFInst_1_n10 ), .ZN(
        SubCellInst_LFInst_13_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_1_U4  ( .A1(AddRoundKeyOutput[52]), 
        .A2(AddRoundKeyOutput[53]), .ZN(SubCellInst_LFInst_13_LFInst_1_n10 )
         );
  INV_X1 SubCellInst_LFInst_13_LFInst_1_U3  ( .A(AddRoundKeyOutput[54]), .ZN(
        SubCellInst_LFInst_13_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_2_U11  ( .A1(
        SubCellInst_LFInst_13_LFInst_2_n22 ), .A2(
        SubCellInst_LFInst_13_LFInst_2_n21 ), .ZN(MCInst_MC2_v0_3 [3]) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_2_U10  ( .A1(AddRoundKeyOutput[54]), 
        .A2(SubCellInst_LFInst_13_LFInst_2_n20 ), .ZN(
        SubCellInst_LFInst_13_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst_LFInst_13_LFInst_2_U9  ( .A1(AddRoundKeyOutput[53]), 
        .A2(SubCellInst_LFInst_13_LFInst_2_n19 ), .ZN(
        SubCellInst_LFInst_13_LFInst_2_n20 ) );
  INV_X1 SubCellInst_LFInst_13_LFInst_2_U8  ( .A(AddRoundKeyOutput[55]), .ZN(
        SubCellInst_LFInst_13_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_2_U7  ( .A1(
        SubCellInst_LFInst_13_LFInst_2_n18 ), .A2(
        SubCellInst_LFInst_13_LFInst_2_n17 ), .ZN(
        SubCellInst_LFInst_13_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst_LFInst_13_LFInst_2_U6  ( .A(
        SubCellInst_LFInst_13_LFInst_2_n16 ), .B(AddRoundKeyOutput[54]), .Z(
        SubCellInst_LFInst_13_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_2_U5  ( .A1(AddRoundKeyOutput[52]), 
        .A2(AddRoundKeyOutput[53]), .ZN(SubCellInst_LFInst_13_LFInst_2_n16 )
         );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_2_U4  ( .A1(
        SubCellInst_LFInst_13_LFInst_2_n15 ), .A2(AddRoundKeyOutput[55]), 
        .ZN(SubCellInst_LFInst_13_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst_LFInst_13_LFInst_2_U3  ( .A(AddRoundKeyOutput[52]), 
        .B(AddRoundKeyOutput[53]), .ZN(SubCellInst_LFInst_13_LFInst_2_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_3_U9  ( .A1(
        SubCellInst_LFInst_13_LFInst_3_n16 ), .A2(
        SubCellInst_LFInst_13_LFInst_3_n15 ), .ZN(MCInst_MC2_v0_3 [0]) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_3_U8  ( .A1(AddRoundKeyOutput[53]), 
        .A2(SubCellInst_LFInst_13_LFInst_3_n14 ), .ZN(
        SubCellInst_LFInst_13_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst_LFInst_13_LFInst_3_U7  ( .A(AddRoundKeyOutput[55]), .B(
        AddRoundKeyOutput[54]), .Z(SubCellInst_LFInst_13_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_3_U6  ( .A1(
        SubCellInst_LFInst_13_LFInst_3_n13 ), .A2(
        SubCellInst_LFInst_13_LFInst_3_n12 ), .ZN(
        SubCellInst_LFInst_13_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_3_U5  ( .A1(AddRoundKeyOutput[52]), 
        .A2(AddRoundKeyOutput[54]), .ZN(SubCellInst_LFInst_13_LFInst_3_n12 )
         );
  XNOR2_X1 SubCellInst_LFInst_13_LFInst_3_U4  ( .A(AddRoundKeyOutput[52]), 
        .B(SubCellInst_LFInst_13_LFInst_3_n11 ), .ZN(
        SubCellInst_LFInst_13_LFInst_3_n13 ) );
  OR2_X1 SubCellInst_LFInst_13_LFInst_3_U3  ( .A1(AddRoundKeyOutput[55]), 
        .A2(AddRoundKeyOutput[53]), .ZN(SubCellInst_LFInst_13_LFInst_3_n11 )
         );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_0_U6  ( .A1(AddRoundKeyOutput[58]), 
        .A2(SubCellInst_LFInst_14_LFInst_0_n4 ), .ZN(
        SubCellInst_LFInst_14_LFInst_0_n5 ) );
  INV_X1 SubCellInst_LFInst_14_LFInst_0_U5  ( .A(AddRoundKeyOutput[57]), .ZN(
        SubCellInst_LFInst_14_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst_LFInst_14_LFInst_0_U4  ( .A(AddRoundKeyOutput[56]), .B(
        AddRoundKeyOutput[59]), .Z(SubCellInst_LFInst_14_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst_LFInst_14_LFInst_0_U3  ( .A(
        SubCellInst_LFInst_14_LFInst_0_n6 ), .B(
        SubCellInst_LFInst_14_LFInst_0_n5 ), .ZN(Red_MCInst_MC1_v0_1[0] ) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_1_U12  ( .A1(
        SubCellInst_LFInst_14_LFInst_1_n18 ), .A2(
        SubCellInst_LFInst_14_LFInst_1_n17 ), .ZN(MCInst_MC1_v0_0 [3]) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_1_U11  ( .A1(AddRoundKeyOutput[57]), 
        .A2(SubCellInst_LFInst_14_LFInst_1_n16 ), .ZN(
        SubCellInst_LFInst_14_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst_LFInst_14_LFInst_1_U10  ( .A1(AddRoundKeyOutput[59]), 
        .A2(SubCellInst_LFInst_14_LFInst_1_n15 ), .ZN(
        SubCellInst_LFInst_14_LFInst_1_n16 ) );
  AND2_X1 SubCellInst_LFInst_14_LFInst_1_U9  ( .A1(AddRoundKeyOutput[56]), 
        .A2(AddRoundKeyOutput[58]), .ZN(SubCellInst_LFInst_14_LFInst_1_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_1_U8  ( .A1(AddRoundKeyOutput[59]), 
        .A2(SubCellInst_LFInst_14_LFInst_1_n14 ), .ZN(
        SubCellInst_LFInst_14_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_1_U7  ( .A1(
        SubCellInst_LFInst_14_LFInst_1_n13 ), .A2(
        SubCellInst_LFInst_14_LFInst_1_n12 ), .ZN(
        SubCellInst_LFInst_14_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_1_U6  ( .A1(AddRoundKeyOutput[56]), 
        .A2(AddRoundKeyOutput[58]), .ZN(SubCellInst_LFInst_14_LFInst_1_n12 )
         );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_1_U5  ( .A1(
        SubCellInst_LFInst_14_LFInst_1_n11 ), .A2(
        SubCellInst_LFInst_14_LFInst_1_n10 ), .ZN(
        SubCellInst_LFInst_14_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_1_U4  ( .A1(AddRoundKeyOutput[56]), 
        .A2(AddRoundKeyOutput[57]), .ZN(SubCellInst_LFInst_14_LFInst_1_n10 )
         );
  INV_X1 SubCellInst_LFInst_14_LFInst_1_U3  ( .A(AddRoundKeyOutput[58]), .ZN(
        SubCellInst_LFInst_14_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_2_U11  ( .A1(
        SubCellInst_LFInst_14_LFInst_2_n22 ), .A2(
        SubCellInst_LFInst_14_LFInst_2_n21 ), .ZN(MCInst_MC1_v0_3 [3]) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_2_U10  ( .A1(AddRoundKeyOutput[58]), 
        .A2(SubCellInst_LFInst_14_LFInst_2_n20 ), .ZN(
        SubCellInst_LFInst_14_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst_LFInst_14_LFInst_2_U9  ( .A1(AddRoundKeyOutput[57]), 
        .A2(SubCellInst_LFInst_14_LFInst_2_n19 ), .ZN(
        SubCellInst_LFInst_14_LFInst_2_n20 ) );
  INV_X1 SubCellInst_LFInst_14_LFInst_2_U8  ( .A(AddRoundKeyOutput[59]), .ZN(
        SubCellInst_LFInst_14_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_2_U7  ( .A1(
        SubCellInst_LFInst_14_LFInst_2_n18 ), .A2(
        SubCellInst_LFInst_14_LFInst_2_n17 ), .ZN(
        SubCellInst_LFInst_14_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst_LFInst_14_LFInst_2_U6  ( .A(
        SubCellInst_LFInst_14_LFInst_2_n16 ), .B(AddRoundKeyOutput[58]), .Z(
        SubCellInst_LFInst_14_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_2_U5  ( .A1(AddRoundKeyOutput[56]), 
        .A2(AddRoundKeyOutput[57]), .ZN(SubCellInst_LFInst_14_LFInst_2_n16 )
         );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_2_U4  ( .A1(
        SubCellInst_LFInst_14_LFInst_2_n15 ), .A2(AddRoundKeyOutput[59]), 
        .ZN(SubCellInst_LFInst_14_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst_LFInst_14_LFInst_2_U3  ( .A(AddRoundKeyOutput[56]), 
        .B(AddRoundKeyOutput[57]), .ZN(SubCellInst_LFInst_14_LFInst_2_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_3_U9  ( .A1(
        SubCellInst_LFInst_14_LFInst_3_n16 ), .A2(
        SubCellInst_LFInst_14_LFInst_3_n15 ), .ZN(MCInst_MC1_v0_3 [0]) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_3_U8  ( .A1(AddRoundKeyOutput[57]), 
        .A2(SubCellInst_LFInst_14_LFInst_3_n14 ), .ZN(
        SubCellInst_LFInst_14_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst_LFInst_14_LFInst_3_U7  ( .A(AddRoundKeyOutput[59]), .B(
        AddRoundKeyOutput[58]), .Z(SubCellInst_LFInst_14_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_3_U6  ( .A1(
        SubCellInst_LFInst_14_LFInst_3_n13 ), .A2(
        SubCellInst_LFInst_14_LFInst_3_n12 ), .ZN(
        SubCellInst_LFInst_14_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_3_U5  ( .A1(AddRoundKeyOutput[56]), 
        .A2(AddRoundKeyOutput[58]), .ZN(SubCellInst_LFInst_14_LFInst_3_n12 )
         );
  XNOR2_X1 SubCellInst_LFInst_14_LFInst_3_U4  ( .A(AddRoundKeyOutput[56]), 
        .B(SubCellInst_LFInst_14_LFInst_3_n11 ), .ZN(
        SubCellInst_LFInst_14_LFInst_3_n13 ) );
  OR2_X1 SubCellInst_LFInst_14_LFInst_3_U3  ( .A1(AddRoundKeyOutput[59]), 
        .A2(AddRoundKeyOutput[57]), .ZN(SubCellInst_LFInst_14_LFInst_3_n11 )
         );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_0_U6  ( .A1(AddRoundKeyOutput[62]), 
        .A2(SubCellInst_LFInst_15_LFInst_0_n4 ), .ZN(
        SubCellInst_LFInst_15_LFInst_0_n5 ) );
  INV_X1 SubCellInst_LFInst_15_LFInst_0_U5  ( .A(AddRoundKeyOutput[61]), .ZN(
        SubCellInst_LFInst_15_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst_LFInst_15_LFInst_0_U4  ( .A(AddRoundKeyOutput[60]), .B(
        AddRoundKeyOutput[63]), .Z(SubCellInst_LFInst_15_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst_LFInst_15_LFInst_0_U3  ( .A(
        SubCellInst_LFInst_15_LFInst_0_n6 ), .B(
        SubCellInst_LFInst_15_LFInst_0_n5 ), .ZN(Red_MCInst_MC0_v0_1[0] ) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_1_U12  ( .A1(
        SubCellInst_LFInst_15_LFInst_1_n18 ), .A2(
        SubCellInst_LFInst_15_LFInst_1_n17 ), .ZN(MCInst_MC0_v0_0 [3]) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_1_U11  ( .A1(AddRoundKeyOutput[61]), 
        .A2(SubCellInst_LFInst_15_LFInst_1_n16 ), .ZN(
        SubCellInst_LFInst_15_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst_LFInst_15_LFInst_1_U10  ( .A1(AddRoundKeyOutput[63]), 
        .A2(SubCellInst_LFInst_15_LFInst_1_n15 ), .ZN(
        SubCellInst_LFInst_15_LFInst_1_n16 ) );
  AND2_X1 SubCellInst_LFInst_15_LFInst_1_U9  ( .A1(AddRoundKeyOutput[60]), 
        .A2(AddRoundKeyOutput[62]), .ZN(SubCellInst_LFInst_15_LFInst_1_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_1_U8  ( .A1(AddRoundKeyOutput[63]), 
        .A2(SubCellInst_LFInst_15_LFInst_1_n14 ), .ZN(
        SubCellInst_LFInst_15_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_1_U7  ( .A1(
        SubCellInst_LFInst_15_LFInst_1_n13 ), .A2(
        SubCellInst_LFInst_15_LFInst_1_n12 ), .ZN(
        SubCellInst_LFInst_15_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_1_U6  ( .A1(AddRoundKeyOutput[60]), 
        .A2(AddRoundKeyOutput[62]), .ZN(SubCellInst_LFInst_15_LFInst_1_n12 )
         );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_1_U5  ( .A1(
        SubCellInst_LFInst_15_LFInst_1_n11 ), .A2(
        SubCellInst_LFInst_15_LFInst_1_n10 ), .ZN(
        SubCellInst_LFInst_15_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_1_U4  ( .A1(AddRoundKeyOutput[60]), 
        .A2(AddRoundKeyOutput[61]), .ZN(SubCellInst_LFInst_15_LFInst_1_n10 )
         );
  INV_X1 SubCellInst_LFInst_15_LFInst_1_U3  ( .A(AddRoundKeyOutput[62]), .ZN(
        SubCellInst_LFInst_15_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_2_U11  ( .A1(
        SubCellInst_LFInst_15_LFInst_2_n22 ), .A2(
        SubCellInst_LFInst_15_LFInst_2_n21 ), .ZN(MCInst_MC0_v0_3 [3]) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_2_U10  ( .A1(AddRoundKeyOutput[62]), 
        .A2(SubCellInst_LFInst_15_LFInst_2_n20 ), .ZN(
        SubCellInst_LFInst_15_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst_LFInst_15_LFInst_2_U9  ( .A1(AddRoundKeyOutput[61]), 
        .A2(SubCellInst_LFInst_15_LFInst_2_n19 ), .ZN(
        SubCellInst_LFInst_15_LFInst_2_n20 ) );
  INV_X1 SubCellInst_LFInst_15_LFInst_2_U8  ( .A(AddRoundKeyOutput[63]), .ZN(
        SubCellInst_LFInst_15_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_2_U7  ( .A1(
        SubCellInst_LFInst_15_LFInst_2_n18 ), .A2(
        SubCellInst_LFInst_15_LFInst_2_n17 ), .ZN(
        SubCellInst_LFInst_15_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst_LFInst_15_LFInst_2_U6  ( .A(
        SubCellInst_LFInst_15_LFInst_2_n16 ), .B(AddRoundKeyOutput[62]), .Z(
        SubCellInst_LFInst_15_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_2_U5  ( .A1(AddRoundKeyOutput[60]), 
        .A2(AddRoundKeyOutput[61]), .ZN(SubCellInst_LFInst_15_LFInst_2_n16 )
         );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_2_U4  ( .A1(
        SubCellInst_LFInst_15_LFInst_2_n15 ), .A2(AddRoundKeyOutput[63]), 
        .ZN(SubCellInst_LFInst_15_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst_LFInst_15_LFInst_2_U3  ( .A(AddRoundKeyOutput[60]), 
        .B(AddRoundKeyOutput[61]), .ZN(SubCellInst_LFInst_15_LFInst_2_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_3_U9  ( .A1(
        SubCellInst_LFInst_15_LFInst_3_n16 ), .A2(
        SubCellInst_LFInst_15_LFInst_3_n15 ), .ZN(MCInst_MC0_v0_3 [0]) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_3_U8  ( .A1(AddRoundKeyOutput[61]), 
        .A2(SubCellInst_LFInst_15_LFInst_3_n14 ), .ZN(
        SubCellInst_LFInst_15_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst_LFInst_15_LFInst_3_U7  ( .A(AddRoundKeyOutput[63]), .B(
        AddRoundKeyOutput[62]), .Z(SubCellInst_LFInst_15_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_3_U6  ( .A1(
        SubCellInst_LFInst_15_LFInst_3_n13 ), .A2(
        SubCellInst_LFInst_15_LFInst_3_n12 ), .ZN(
        SubCellInst_LFInst_15_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_3_U5  ( .A1(AddRoundKeyOutput[60]), 
        .A2(AddRoundKeyOutput[62]), .ZN(SubCellInst_LFInst_15_LFInst_3_n12 )
         );
  XNOR2_X1 SubCellInst_LFInst_15_LFInst_3_U4  ( .A(AddRoundKeyOutput[60]), 
        .B(SubCellInst_LFInst_15_LFInst_3_n11 ), .ZN(
        SubCellInst_LFInst_15_LFInst_3_n13 ) );
  OR2_X1 SubCellInst_LFInst_15_LFInst_3_U3  ( .A1(AddRoundKeyOutput[63]), 
        .A2(AddRoundKeyOutput[61]), .ZN(SubCellInst_LFInst_15_LFInst_3_n11 )
         );
  XNOR2_X1 MCInst_MC0_v0_2Inst_0_U4  ( .A(MCInst_MC0_v0_2Inst_0_n2 ), .B(
        MCInst_MC0_v0_0 [3]), .ZN(MCInst_MC0_v0_2 [0]) );
  XNOR2_X1 MCInst_MC0_v0_2Inst_0_U3  ( .A(MCInst_MC0_v0_3 [0]), .B(
        Red_MCInst_MC0_v0_1[0] ), .ZN(MCInst_MC0_v0_2Inst_0_n2 ) );
  XOR2_X1 MCInst_MC0_v1_1Inst_0_U3  ( .A(Red_MCInst_MC0_v1_1[0] ), .B(
        MCInst_MC0_v1_0 [3]), .Z(MCInst_MC0_v1_1 [0]) );
  XNOR2_X1 MCInst_MC0_v1_2Inst_0_U4  ( .A(MCInst_MC0_v1_2Inst_0_n2 ), .B(
        Red_MCInst_MC0_v1_1[0] ), .ZN(MCInst_MC0_v1_2 [0]) );
  XNOR2_X1 MCInst_MC0_v1_2Inst_0_U3  ( .A(MCInst_MC0_v1_0 [3]), .B(
        MCInst_MC0_v1_3 [2]), .ZN(MCInst_MC0_v1_2Inst_0_n2 ) );
  XOR2_X1 MCInst_MC0_v2_1Inst_0_U3  ( .A(MCInst_MC0_v2_3 [1]), .B(
        MCInst_MC0_v2_0 [3]), .Z(MCInst_MC0_v2_1 [0]) );
  XOR2_X1 MCInst_MC0_v2_2Inst_0_U3  ( .A(MCInst_MC0_v2_0 [2]), .B(
        MCInst_MC0_v2_0 [0]), .Z(MCInst_MC0_v2_2 [0]) );
  XNOR2_X1 MCInst_MC0_v2_3Inst_0_U5  ( .A(MCInst_MC0_v2_3Inst_0_n4 ), .B(
        MCInst_MC0_v2_3Inst_0_n3 ), .ZN(MCInst_MC0_v2_3 [0]) );
  XNOR2_X1 MCInst_MC0_v2_3Inst_0_U4  ( .A(MCInst_MC0_v2_0 [2]), .B(
        MCInst_MC0_v2_3 [1]), .ZN(MCInst_MC0_v2_3Inst_0_n3 ) );
  XOR2_X1 MCInst_MC0_v2_3Inst_0_U3  ( .A(MCInst_MC0_v2_0 [3]), .B(
        MCInst_MC0_v2_0 [0]), .Z(MCInst_MC0_v2_3Inst_0_n4 ) );
  XOR2_X1 MCInst_MC0_v3_1Inst_0_U3  ( .A(Red_MCInst_MC0_v3_1[0] ), .B(
        MCInst_MC0_v3_2 [2]), .Z(MCInst_MC0_v3_1 [0]) );
  XOR2_X1 MCInst_MC0_v3_2Inst_0_U3  ( .A(MCInst_MC0_v3_2 [3]), .B(
        MCInst_MC0_v3_0 [2]), .Z(MCInst_MC0_v3_2 [0]) );
  XNOR2_X1 MCInst_MC0_v3_3Inst_0_U4  ( .A(MCInst_MC0_v3_3Inst_0_n2 ), .B(
        MCInst_MC0_v3_0 [2]), .ZN(MCInst_MC0_v3_3 [0]) );
  XNOR2_X1 MCInst_MC0_v3_3Inst_0_U3  ( .A(MCInst_MC0_v3_2 [2]), .B(
        MCInst_MC0_v3_2 [3]), .ZN(MCInst_MC0_v3_3Inst_0_n2 ) );
  XOR2_X1 MCInst_MC0_v0_0Inst_1_U3  ( .A(MCInst_MC0_v0_3 [3]), .B(
        MCInst_MC0_v0_3 [0]), .Z(MCInst_MC0_v0_0 [1]) );
  XOR2_X1 MCInst_MC0_v0_1Inst_1_U3  ( .A(MCInst_MC0_v0_0 [3]), .B(
        MCInst_MC0_v0_3 [3]), .Z(MCInst_MC0_v0_1 [1]) );
  XNOR2_X1 MCInst_MC0_v0_2Inst_1_U4  ( .A(MCInst_MC0_v0_2Inst_1_n2 ), .B(
        MCInst_MC0_v0_3 [3]), .ZN(MCInst_MC0_v0_2 [1]) );
  XNOR2_X1 MCInst_MC0_v0_2Inst_1_U3  ( .A(MCInst_MC0_v0_3 [0]), .B(
        Red_MCInst_MC0_v0_1[0] ), .ZN(MCInst_MC0_v0_2Inst_1_n2 ) );
  XOR2_X1 MCInst_MC0_v0_3Inst_1_U3  ( .A(Red_MCInst_MC0_v0_1[0] ), .B(
        MCInst_MC0_v0_3 [0]), .Z(MCInst_MC0_v0_3 [1]) );
  XOR2_X1 MCInst_MC0_v1_1Inst_1_U3  ( .A(MCInst_MC0_v1_0 [0]), .B(
        Red_MCInst_MC0_v1_1[0] ), .Z(MCInst_MC0_v1_1 [1]) );
  XOR2_X1 MCInst_MC0_v1_2Inst_1_U3  ( .A(MCInst_MC0_v1_0 [0]), .B(
        MCInst_MC0_v1_3 [2]), .Z(MCInst_MC0_v1_2 [1]) );
  XOR2_X1 MCInst_MC0_v1_3Inst_1_U3  ( .A(MCInst_MC0_v1_0 [0]), .B(
        MCInst_MC0_v1_0 [3]), .Z(MCInst_MC0_v1_3 [1]) );
  XOR2_X1 MCInst_MC0_v2_0Inst_1_U3  ( .A(MCInst_MC0_v2_3 [1]), .B(
        MCInst_MC0_v2_0 [0]), .Z(MCInst_MC0_v2_0 [1]) );
  XNOR2_X1 MCInst_MC0_v2_1Inst_1_U4  ( .A(MCInst_MC0_v2_1Inst_1_n2 ), .B(
        MCInst_MC0_v2_0 [3]), .ZN(MCInst_MC0_v2_1 [1]) );
  XNOR2_X1 MCInst_MC0_v2_1Inst_1_U3  ( .A(MCInst_MC0_v2_0 [0]), .B(
        MCInst_MC0_v2_0 [2]), .ZN(MCInst_MC0_v2_1Inst_1_n2 ) );
  XNOR2_X1 MCInst_MC0_v2_2Inst_1_U5  ( .A(MCInst_MC0_v2_2Inst_1_n4 ), .B(
        MCInst_MC0_v2_2Inst_1_n3 ), .ZN(MCInst_MC0_v2_2 [1]) );
  XNOR2_X1 MCInst_MC0_v2_2Inst_1_U4  ( .A(MCInst_MC0_v2_0 [2]), .B(
        MCInst_MC0_v2_3 [1]), .ZN(MCInst_MC0_v2_2Inst_1_n3 ) );
  XOR2_X1 MCInst_MC0_v2_2Inst_1_U3  ( .A(MCInst_MC0_v2_0 [3]), .B(
        MCInst_MC0_v2_0 [0]), .Z(MCInst_MC0_v2_2Inst_1_n4 ) );
  XOR2_X1 MCInst_MC0_v3_0Inst_1_U3  ( .A(MCInst_MC0_v3_2 [3]), .B(
        MCInst_MC0_v3_2 [2]), .Z(MCInst_MC0_v3_0 [1]) );
  XOR2_X1 MCInst_MC0_v3_1Inst_1_U3  ( .A(MCInst_MC0_v3_2 [3]), .B(
        Red_MCInst_MC0_v3_1[0] ), .Z(MCInst_MC0_v3_1 [1]) );
  XNOR2_X1 MCInst_MC0_v3_3Inst_1_U4  ( .A(MCInst_MC0_v3_3Inst_1_n2 ), .B(
        Red_MCInst_MC0_v3_1[0] ), .ZN(MCInst_MC0_v3_3 [1]) );
  XNOR2_X1 MCInst_MC0_v3_3Inst_1_U3  ( .A(MCInst_MC0_v3_2 [2]), .B(
        MCInst_MC0_v3_2 [3]), .ZN(MCInst_MC0_v3_3Inst_1_n2 ) );
  XOR2_X1 MCInst_MC0_v0_0Inst_2_U3  ( .A(Red_MCInst_MC0_v0_1[0] ), .B(
        MCInst_MC0_v0_3 [0]), .Z(MCInst_MC0_v0_0 [2]) );
  XOR2_X1 MCInst_MC0_v0_1Inst_2_U3  ( .A(MCInst_MC0_v0_3 [3]), .B(
        MCInst_MC0_v0_3 [0]), .Z(MCInst_MC0_v0_1 [2]) );
  XOR2_X1 MCInst_MC0_v0_2Inst_2_U3  ( .A(MCInst_MC0_v0_0 [3]), .B(
        MCInst_MC0_v0_3 [0]), .Z(MCInst_MC0_v0_2 [2]) );
  XNOR2_X1 MCInst_MC0_v1_1Inst_2_U4  ( .A(MCInst_MC0_v1_1Inst_2_n2 ), .B(
        MCInst_MC0_v1_3 [2]), .ZN(MCInst_MC0_v1_1 [2]) );
  XNOR2_X1 MCInst_MC0_v1_1Inst_2_U3  ( .A(MCInst_MC0_v1_0 [3]), .B(
        MCInst_MC0_v1_0 [0]), .ZN(MCInst_MC0_v1_1Inst_2_n2 ) );
  XNOR2_X1 MCInst_MC0_v1_2Inst_2_U4  ( .A(MCInst_MC0_v1_2Inst_2_n2 ), .B(
        MCInst_MC0_v1_3 [2]), .ZN(MCInst_MC0_v1_2 [2]) );
  XNOR2_X1 MCInst_MC0_v1_2Inst_2_U3  ( .A(Red_MCInst_MC0_v1_1[0] ), .B(
        MCInst_MC0_v1_0 [0]), .ZN(MCInst_MC0_v1_2Inst_2_n2 ) );
  XNOR2_X1 MCInst_MC0_v2_1Inst_2_U4  ( .A(MCInst_MC0_v2_1Inst_2_n2 ), .B(
        MCInst_MC0_v2_0 [3]), .ZN(MCInst_MC0_v2_1 [2]) );
  XNOR2_X1 MCInst_MC0_v2_1Inst_2_U3  ( .A(MCInst_MC0_v2_0 [0]), .B(
        MCInst_MC0_v2_3 [1]), .ZN(MCInst_MC0_v2_1Inst_2_n2 ) );
  XNOR2_X1 MCInst_MC0_v2_2Inst_2_U4  ( .A(MCInst_MC0_v2_2Inst_2_n2 ), .B(
        MCInst_MC0_v2_0 [3]), .ZN(MCInst_MC0_v2_2 [2]) );
  XNOR2_X1 MCInst_MC0_v2_2Inst_2_U3  ( .A(MCInst_MC0_v2_0 [0]), .B(
        MCInst_MC0_v2_0 [2]), .ZN(MCInst_MC0_v2_2Inst_2_n2 ) );
  XOR2_X1 MCInst_MC0_v2_3Inst_2_U3  ( .A(MCInst_MC0_v2_3 [1]), .B(
        MCInst_MC0_v2_0 [2]), .Z(MCInst_MC0_v2_3 [2]) );
  XNOR2_X1 MCInst_MC0_v3_1Inst_2_U4  ( .A(MCInst_MC0_v3_1Inst_2_n2 ), .B(
        MCInst_MC0_v3_0 [2]), .ZN(MCInst_MC0_v3_1 [2]) );
  XNOR2_X1 MCInst_MC0_v3_1Inst_2_U3  ( .A(MCInst_MC0_v3_2 [2]), .B(
        MCInst_MC0_v3_2 [3]), .ZN(MCInst_MC0_v3_1Inst_2_n2 ) );
  XOR2_X1 MCInst_MC0_v3_3Inst_2_U3  ( .A(MCInst_MC0_v3_0 [2]), .B(
        MCInst_MC0_v3_2 [2]), .Z(MCInst_MC0_v3_3 [2]) );
  XOR2_X1 MCInst_MC0_v0_1Inst_3_U3  ( .A(Red_MCInst_MC0_v0_1[0] ), .B(
        MCInst_MC0_v0_3 [0]), .Z(MCInst_MC0_v0_1 [3]) );
  XOR2_X1 MCInst_MC0_v0_2Inst_3_U3  ( .A(Red_MCInst_MC0_v0_1[0] ), .B(
        MCInst_MC0_v0_3 [3]), .Z(MCInst_MC0_v0_2 [3]) );
  XOR2_X1 MCInst_MC0_v1_1Inst_3_U3  ( .A(MCInst_MC0_v1_3 [2]), .B(
        Red_MCInst_MC0_v1_1[0] ), .Z(MCInst_MC0_v1_1 [3]) );
  XNOR2_X1 MCInst_MC0_v1_2Inst_3_U5  ( .A(MCInst_MC0_v1_2Inst_3_n4 ), .B(
        MCInst_MC0_v1_2Inst_3_n3 ), .ZN(MCInst_MC0_v1_2 [3]) );
  XNOR2_X1 MCInst_MC0_v1_2Inst_3_U4  ( .A(MCInst_MC0_v1_3 [2]), .B(
        MCInst_MC0_v1_0 [0]), .ZN(MCInst_MC0_v1_2Inst_3_n3 ) );
  XOR2_X1 MCInst_MC0_v1_2Inst_3_U3  ( .A(Red_MCInst_MC0_v1_1[0] ), .B(
        MCInst_MC0_v1_0 [3]), .Z(MCInst_MC0_v1_2Inst_3_n4 ) );
  XOR2_X1 MCInst_MC0_v2_1Inst_3_U3  ( .A(MCInst_MC0_v2_0 [2]), .B(
        MCInst_MC0_v2_0 [0]), .Z(MCInst_MC0_v2_1 [3]) );
  XNOR2_X1 MCInst_MC0_v2_2Inst_3_U4  ( .A(MCInst_MC0_v2_2Inst_3_n2 ), .B(
        MCInst_MC0_v2_0 [3]), .ZN(MCInst_MC0_v2_2 [3]) );
  XNOR2_X1 MCInst_MC0_v2_2Inst_3_U3  ( .A(MCInst_MC0_v2_0 [0]), .B(
        MCInst_MC0_v2_3 [1]), .ZN(MCInst_MC0_v2_2Inst_3_n2 ) );
  XNOR2_X1 MCInst_MC0_v2_3Inst_3_U4  ( .A(MCInst_MC0_v2_3Inst_3_n2 ), .B(
        MCInst_MC0_v2_0 [2]), .ZN(MCInst_MC0_v2_3 [3]) );
  XNOR2_X1 MCInst_MC0_v2_3Inst_3_U3  ( .A(MCInst_MC0_v2_0 [3]), .B(
        MCInst_MC0_v2_3 [1]), .ZN(MCInst_MC0_v2_3Inst_3_n2 ) );
  XOR2_X1 MCInst_MC0_v3_1Inst_3_U3  ( .A(MCInst_MC0_v3_0 [2]), .B(
        Red_MCInst_MC0_v3_1[0] ), .Z(MCInst_MC0_v3_1 [3]) );
  XOR2_X1 MCInst_MC0_v3_3Inst_3_U3  ( .A(MCInst_MC0_v3_2 [3]), .B(
        Red_MCInst_MC0_v3_1[0] ), .Z(MCInst_MC0_v3_3 [3]) );
  XNOR2_X1 MCInst_MC0_r0Inst_XORInst_0_0_U3  ( .A(
        MCInst_MC0_r0Inst_XORInst_0_0_n5 ), .B(
        MCInst_MC0_r0Inst_XORInst_0_0_n4 ), .ZN(Feedback[60]) );
  XNOR2_X1 MCInst_MC0_r0Inst_XORInst_0_0_U2  ( .A(MCInst_MC0_v3_2 [2]), .B(
        MCInst_MC0_v2_0 [0]), .ZN(MCInst_MC0_r0Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst_MC0_r0Inst_XORInst_0_0_U1  ( .A(MCInst_MC0_v0_3 [3]), .B(
        MCInst_MC0_v1_0 [0]), .Z(MCInst_MC0_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst_MC0_r0Inst_XORInst_0_1_U3  ( .A(
        MCInst_MC0_r0Inst_XORInst_0_1_n5 ), .B(
        MCInst_MC0_r0Inst_XORInst_0_1_n4 ), .ZN(Feedback[61]) );
  XNOR2_X1 MCInst_MC0_r0Inst_XORInst_0_1_U2  ( .A(MCInst_MC0_v3_0 [1]), .B(
        MCInst_MC0_v2_0 [1]), .ZN(MCInst_MC0_r0Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst_MC0_r0Inst_XORInst_0_1_U1  ( .A(MCInst_MC0_v0_0 [1]), .B(
        MCInst_MC0_v1_3 [2]), .Z(MCInst_MC0_r0Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst_MC0_r0Inst_XORInst_0_2_U3  ( .A(
        MCInst_MC0_r0Inst_XORInst_0_2_n5 ), .B(
        MCInst_MC0_r0Inst_XORInst_0_2_n4 ), .ZN(Feedback[62]) );
  XNOR2_X1 MCInst_MC0_r0Inst_XORInst_0_2_U2  ( .A(MCInst_MC0_v3_0 [2]), .B(
        MCInst_MC0_v2_0 [2]), .ZN(MCInst_MC0_r0Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst_MC0_r0Inst_XORInst_0_2_U1  ( .A(MCInst_MC0_v0_0 [2]), .B(
        Red_MCInst_MC0_v1_1[0] ), .Z(MCInst_MC0_r0Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst_MC0_r0Inst_XORInst_0_3_U3  ( .A(
        MCInst_MC0_r0Inst_XORInst_0_3_n5 ), .B(
        MCInst_MC0_r0Inst_XORInst_0_3_n4 ), .ZN(Feedback[63]) );
  XNOR2_X1 MCInst_MC0_r0Inst_XORInst_0_3_U2  ( .A(Red_MCInst_MC0_v3_1[0] ), 
        .B(MCInst_MC0_v2_0 [3]), .ZN(MCInst_MC0_r0Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst_MC0_r0Inst_XORInst_0_3_U1  ( .A(MCInst_MC0_v0_0 [3]), .B(
        MCInst_MC0_v1_0 [3]), .Z(MCInst_MC0_r0Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst_MC0_r1Inst_XORInst_0_0_U3  ( .A(
        MCInst_MC0_r1Inst_XORInst_0_0_n5 ), .B(
        MCInst_MC0_r1Inst_XORInst_0_0_n4 ), .ZN(Feedback[44]) );
  XNOR2_X1 MCInst_MC0_r1Inst_XORInst_0_0_U2  ( .A(MCInst_MC0_v3_1 [0]), .B(
        MCInst_MC0_v2_1 [0]), .ZN(MCInst_MC0_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst_MC0_r1Inst_XORInst_0_0_U1  ( .A(MCInst_MC0_v0_0 [3]), .B(
        MCInst_MC0_v1_1 [0]), .Z(MCInst_MC0_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst_MC0_r1Inst_XORInst_0_1_U3  ( .A(
        MCInst_MC0_r1Inst_XORInst_0_1_n5 ), .B(
        MCInst_MC0_r1Inst_XORInst_0_1_n4 ), .ZN(Feedback[45]) );
  XNOR2_X1 MCInst_MC0_r1Inst_XORInst_0_1_U2  ( .A(MCInst_MC0_v3_1 [1]), .B(
        MCInst_MC0_v2_1 [1]), .ZN(MCInst_MC0_r1Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst_MC0_r1Inst_XORInst_0_1_U1  ( .A(MCInst_MC0_v0_1 [1]), .B(
        MCInst_MC0_v1_1 [1]), .Z(MCInst_MC0_r1Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst_MC0_r1Inst_XORInst_0_2_U3  ( .A(
        MCInst_MC0_r1Inst_XORInst_0_2_n5 ), .B(
        MCInst_MC0_r1Inst_XORInst_0_2_n4 ), .ZN(Feedback[46]) );
  XNOR2_X1 MCInst_MC0_r1Inst_XORInst_0_2_U2  ( .A(MCInst_MC0_v3_1 [2]), .B(
        MCInst_MC0_v2_1 [2]), .ZN(MCInst_MC0_r1Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst_MC0_r1Inst_XORInst_0_2_U1  ( .A(MCInst_MC0_v0_1 [2]), .B(
        MCInst_MC0_v1_1 [2]), .Z(MCInst_MC0_r1Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst_MC0_r1Inst_XORInst_0_3_U3  ( .A(
        MCInst_MC0_r1Inst_XORInst_0_3_n5 ), .B(
        MCInst_MC0_r1Inst_XORInst_0_3_n4 ), .ZN(Feedback[47]) );
  XNOR2_X1 MCInst_MC0_r1Inst_XORInst_0_3_U2  ( .A(MCInst_MC0_v3_1 [3]), .B(
        MCInst_MC0_v2_1 [3]), .ZN(MCInst_MC0_r1Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst_MC0_r1Inst_XORInst_0_3_U1  ( .A(MCInst_MC0_v0_1 [3]), .B(
        MCInst_MC0_v1_1 [3]), .Z(MCInst_MC0_r1Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst_MC0_r2Inst_XORInst_0_0_U3  ( .A(
        MCInst_MC0_r2Inst_XORInst_0_0_n5 ), .B(
        MCInst_MC0_r2Inst_XORInst_0_0_n4 ), .ZN(Feedback[28]) );
  XNOR2_X1 MCInst_MC0_r2Inst_XORInst_0_0_U2  ( .A(MCInst_MC0_v3_2 [0]), .B(
        MCInst_MC0_v2_2 [0]), .ZN(MCInst_MC0_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst_MC0_r2Inst_XORInst_0_0_U1  ( .A(MCInst_MC0_v0_2 [0]), .B(
        MCInst_MC0_v1_2 [0]), .Z(MCInst_MC0_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst_MC0_r2Inst_XORInst_0_1_U3  ( .A(
        MCInst_MC0_r2Inst_XORInst_0_1_n5 ), .B(
        MCInst_MC0_r2Inst_XORInst_0_1_n4 ), .ZN(Feedback[29]) );
  XNOR2_X1 MCInst_MC0_r2Inst_XORInst_0_1_U2  ( .A(Red_MCInst_MC0_v3_1[0] ), 
        .B(MCInst_MC0_v2_2 [1]), .ZN(MCInst_MC0_r2Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst_MC0_r2Inst_XORInst_0_1_U1  ( .A(MCInst_MC0_v0_2 [1]), .B(
        MCInst_MC0_v1_2 [1]), .Z(MCInst_MC0_r2Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst_MC0_r2Inst_XORInst_0_2_U3  ( .A(
        MCInst_MC0_r2Inst_XORInst_0_2_n5 ), .B(
        MCInst_MC0_r2Inst_XORInst_0_2_n4 ), .ZN(Feedback[30]) );
  XNOR2_X1 MCInst_MC0_r2Inst_XORInst_0_2_U2  ( .A(MCInst_MC0_v3_2 [2]), .B(
        MCInst_MC0_v2_2 [2]), .ZN(MCInst_MC0_r2Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst_MC0_r2Inst_XORInst_0_2_U1  ( .A(MCInst_MC0_v0_2 [2]), .B(
        MCInst_MC0_v1_2 [2]), .Z(MCInst_MC0_r2Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst_MC0_r2Inst_XORInst_0_3_U3  ( .A(
        MCInst_MC0_r2Inst_XORInst_0_3_n5 ), .B(
        MCInst_MC0_r2Inst_XORInst_0_3_n4 ), .ZN(Feedback[31]) );
  XNOR2_X1 MCInst_MC0_r2Inst_XORInst_0_3_U2  ( .A(MCInst_MC0_v3_2 [3]), .B(
        MCInst_MC0_v2_2 [3]), .ZN(MCInst_MC0_r2Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst_MC0_r2Inst_XORInst_0_3_U1  ( .A(MCInst_MC0_v0_2 [3]), .B(
        MCInst_MC0_v1_2 [3]), .Z(MCInst_MC0_r2Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst_MC0_r3Inst_XORInst_0_0_U3  ( .A(
        MCInst_MC0_r3Inst_XORInst_0_0_n5 ), .B(
        MCInst_MC0_r3Inst_XORInst_0_0_n4 ), .ZN(Feedback[12]) );
  XNOR2_X1 MCInst_MC0_r3Inst_XORInst_0_0_U2  ( .A(MCInst_MC0_v3_3 [0]), .B(
        MCInst_MC0_v2_3 [0]), .ZN(MCInst_MC0_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst_MC0_r3Inst_XORInst_0_0_U1  ( .A(MCInst_MC0_v0_3 [0]), .B(
        MCInst_MC0_v1_0 [3]), .Z(MCInst_MC0_r3Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst_MC0_r3Inst_XORInst_0_1_U3  ( .A(
        MCInst_MC0_r3Inst_XORInst_0_1_n5 ), .B(
        MCInst_MC0_r3Inst_XORInst_0_1_n4 ), .ZN(Feedback[13]) );
  XNOR2_X1 MCInst_MC0_r3Inst_XORInst_0_1_U2  ( .A(MCInst_MC0_v3_3 [1]), .B(
        MCInst_MC0_v2_3 [1]), .ZN(MCInst_MC0_r3Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst_MC0_r3Inst_XORInst_0_1_U1  ( .A(MCInst_MC0_v0_3 [1]), .B(
        MCInst_MC0_v1_3 [1]), .Z(MCInst_MC0_r3Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst_MC0_r3Inst_XORInst_0_2_U3  ( .A(
        MCInst_MC0_r3Inst_XORInst_0_2_n5 ), .B(
        MCInst_MC0_r3Inst_XORInst_0_2_n4 ), .ZN(Feedback[14]) );
  XNOR2_X1 MCInst_MC0_r3Inst_XORInst_0_2_U2  ( .A(MCInst_MC0_v3_3 [2]), .B(
        MCInst_MC0_v2_3 [2]), .ZN(MCInst_MC0_r3Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst_MC0_r3Inst_XORInst_0_2_U1  ( .A(MCInst_MC0_v0_0 [3]), .B(
        MCInst_MC0_v1_3 [2]), .Z(MCInst_MC0_r3Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst_MC0_r3Inst_XORInst_0_3_U3  ( .A(
        MCInst_MC0_r3Inst_XORInst_0_3_n5 ), .B(
        MCInst_MC0_r3Inst_XORInst_0_3_n4 ), .ZN(Feedback[15]) );
  XNOR2_X1 MCInst_MC0_r3Inst_XORInst_0_3_U2  ( .A(MCInst_MC0_v3_3 [3]), .B(
        MCInst_MC0_v2_3 [3]), .ZN(MCInst_MC0_r3Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst_MC0_r3Inst_XORInst_0_3_U1  ( .A(MCInst_MC0_v0_3 [3]), .B(
        Red_MCInst_MC0_v1_1[0] ), .Z(MCInst_MC0_r3Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst_MC1_v0_2Inst_0_U4  ( .A(MCInst_MC1_v0_2Inst_0_n2 ), .B(
        MCInst_MC1_v0_0 [3]), .ZN(MCInst_MC1_v0_2 [0]) );
  XNOR2_X1 MCInst_MC1_v0_2Inst_0_U3  ( .A(MCInst_MC1_v0_3 [0]), .B(
        Red_MCInst_MC1_v0_1[0] ), .ZN(MCInst_MC1_v0_2Inst_0_n2 ) );
  XOR2_X1 MCInst_MC1_v1_1Inst_0_U3  ( .A(Red_MCInst_MC1_v1_1[0] ), .B(
        MCInst_MC1_v1_0 [3]), .Z(MCInst_MC1_v1_1 [0]) );
  XNOR2_X1 MCInst_MC1_v1_2Inst_0_U4  ( .A(MCInst_MC1_v1_2Inst_0_n2 ), .B(
        Red_MCInst_MC1_v1_1[0] ), .ZN(MCInst_MC1_v1_2 [0]) );
  XNOR2_X1 MCInst_MC1_v1_2Inst_0_U3  ( .A(MCInst_MC1_v1_0 [3]), .B(
        MCInst_MC1_v1_3 [2]), .ZN(MCInst_MC1_v1_2Inst_0_n2 ) );
  XOR2_X1 MCInst_MC1_v2_1Inst_0_U3  ( .A(MCInst_MC1_v2_3 [1]), .B(
        MCInst_MC1_v2_0 [3]), .Z(MCInst_MC1_v2_1 [0]) );
  XOR2_X1 MCInst_MC1_v2_2Inst_0_U3  ( .A(MCInst_MC1_v2_0 [2]), .B(
        MCInst_MC1_v2_0 [0]), .Z(MCInst_MC1_v2_2 [0]) );
  XNOR2_X1 MCInst_MC1_v2_3Inst_0_U5  ( .A(MCInst_MC1_v2_3Inst_0_n4 ), .B(
        MCInst_MC1_v2_3Inst_0_n3 ), .ZN(MCInst_MC1_v2_3 [0]) );
  XNOR2_X1 MCInst_MC1_v2_3Inst_0_U4  ( .A(MCInst_MC1_v2_0 [2]), .B(
        MCInst_MC1_v2_3 [1]), .ZN(MCInst_MC1_v2_3Inst_0_n3 ) );
  XOR2_X1 MCInst_MC1_v2_3Inst_0_U3  ( .A(MCInst_MC1_v2_0 [3]), .B(
        MCInst_MC1_v2_0 [0]), .Z(MCInst_MC1_v2_3Inst_0_n4 ) );
  XOR2_X1 MCInst_MC1_v3_1Inst_0_U3  ( .A(Red_MCInst_MC1_v3_1[0] ), .B(
        MCInst_MC1_v3_2 [2]), .Z(MCInst_MC1_v3_1 [0]) );
  XOR2_X1 MCInst_MC1_v3_2Inst_0_U3  ( .A(MCInst_MC1_v3_2 [3]), .B(
        MCInst_MC1_v3_0 [2]), .Z(MCInst_MC1_v3_2 [0]) );
  XNOR2_X1 MCInst_MC1_v3_3Inst_0_U4  ( .A(MCInst_MC1_v3_3Inst_0_n2 ), .B(
        MCInst_MC1_v3_0 [2]), .ZN(MCInst_MC1_v3_3 [0]) );
  XNOR2_X1 MCInst_MC1_v3_3Inst_0_U3  ( .A(MCInst_MC1_v3_2 [2]), .B(
        MCInst_MC1_v3_2 [3]), .ZN(MCInst_MC1_v3_3Inst_0_n2 ) );
  XOR2_X1 MCInst_MC1_v0_0Inst_1_U3  ( .A(MCInst_MC1_v0_3 [3]), .B(
        MCInst_MC1_v0_3 [0]), .Z(MCInst_MC1_v0_0 [1]) );
  XOR2_X1 MCInst_MC1_v0_1Inst_1_U3  ( .A(MCInst_MC1_v0_0 [3]), .B(
        MCInst_MC1_v0_3 [3]), .Z(MCInst_MC1_v0_1 [1]) );
  XNOR2_X1 MCInst_MC1_v0_2Inst_1_U4  ( .A(MCInst_MC1_v0_2Inst_1_n2 ), .B(
        MCInst_MC1_v0_3 [3]), .ZN(MCInst_MC1_v0_2 [1]) );
  XNOR2_X1 MCInst_MC1_v0_2Inst_1_U3  ( .A(MCInst_MC1_v0_3 [0]), .B(
        Red_MCInst_MC1_v0_1[0] ), .ZN(MCInst_MC1_v0_2Inst_1_n2 ) );
  XOR2_X1 MCInst_MC1_v0_3Inst_1_U3  ( .A(Red_MCInst_MC1_v0_1[0] ), .B(
        MCInst_MC1_v0_3 [0]), .Z(MCInst_MC1_v0_3 [1]) );
  XOR2_X1 MCInst_MC1_v1_1Inst_1_U3  ( .A(MCInst_MC1_v1_0 [0]), .B(
        Red_MCInst_MC1_v1_1[0] ), .Z(MCInst_MC1_v1_1 [1]) );
  XOR2_X1 MCInst_MC1_v1_2Inst_1_U3  ( .A(MCInst_MC1_v1_0 [0]), .B(
        MCInst_MC1_v1_3 [2]), .Z(MCInst_MC1_v1_2 [1]) );
  XOR2_X1 MCInst_MC1_v1_3Inst_1_U3  ( .A(MCInst_MC1_v1_0 [0]), .B(
        MCInst_MC1_v1_0 [3]), .Z(MCInst_MC1_v1_3 [1]) );
  XOR2_X1 MCInst_MC1_v2_0Inst_1_U3  ( .A(MCInst_MC1_v2_3 [1]), .B(
        MCInst_MC1_v2_0 [0]), .Z(MCInst_MC1_v2_0 [1]) );
  XNOR2_X1 MCInst_MC1_v2_1Inst_1_U4  ( .A(MCInst_MC1_v2_1Inst_1_n2 ), .B(
        MCInst_MC1_v2_0 [3]), .ZN(MCInst_MC1_v2_1 [1]) );
  XNOR2_X1 MCInst_MC1_v2_1Inst_1_U3  ( .A(MCInst_MC1_v2_0 [0]), .B(
        MCInst_MC1_v2_0 [2]), .ZN(MCInst_MC1_v2_1Inst_1_n2 ) );
  XNOR2_X1 MCInst_MC1_v2_2Inst_1_U5  ( .A(MCInst_MC1_v2_2Inst_1_n4 ), .B(
        MCInst_MC1_v2_2Inst_1_n3 ), .ZN(MCInst_MC1_v2_2 [1]) );
  XNOR2_X1 MCInst_MC1_v2_2Inst_1_U4  ( .A(MCInst_MC1_v2_0 [2]), .B(
        MCInst_MC1_v2_3 [1]), .ZN(MCInst_MC1_v2_2Inst_1_n3 ) );
  XOR2_X1 MCInst_MC1_v2_2Inst_1_U3  ( .A(MCInst_MC1_v2_0 [3]), .B(
        MCInst_MC1_v2_0 [0]), .Z(MCInst_MC1_v2_2Inst_1_n4 ) );
  XOR2_X1 MCInst_MC1_v3_0Inst_1_U3  ( .A(MCInst_MC1_v3_2 [3]), .B(
        MCInst_MC1_v3_2 [2]), .Z(MCInst_MC1_v3_0 [1]) );
  XOR2_X1 MCInst_MC1_v3_1Inst_1_U3  ( .A(MCInst_MC1_v3_2 [3]), .B(
        Red_MCInst_MC1_v3_1[0] ), .Z(MCInst_MC1_v3_1 [1]) );
  XNOR2_X1 MCInst_MC1_v3_3Inst_1_U4  ( .A(MCInst_MC1_v3_3Inst_1_n2 ), .B(
        Red_MCInst_MC1_v3_1[0] ), .ZN(MCInst_MC1_v3_3 [1]) );
  XNOR2_X1 MCInst_MC1_v3_3Inst_1_U3  ( .A(MCInst_MC1_v3_2 [2]), .B(
        MCInst_MC1_v3_2 [3]), .ZN(MCInst_MC1_v3_3Inst_1_n2 ) );
  XOR2_X1 MCInst_MC1_v0_0Inst_2_U3  ( .A(Red_MCInst_MC1_v0_1[0] ), .B(
        MCInst_MC1_v0_3 [0]), .Z(MCInst_MC1_v0_0 [2]) );
  XOR2_X1 MCInst_MC1_v0_1Inst_2_U3  ( .A(MCInst_MC1_v0_3 [3]), .B(
        MCInst_MC1_v0_3 [0]), .Z(MCInst_MC1_v0_1 [2]) );
  XOR2_X1 MCInst_MC1_v0_2Inst_2_U3  ( .A(MCInst_MC1_v0_0 [3]), .B(
        MCInst_MC1_v0_3 [0]), .Z(MCInst_MC1_v0_2 [2]) );
  XNOR2_X1 MCInst_MC1_v1_1Inst_2_U4  ( .A(MCInst_MC1_v1_1Inst_2_n2 ), .B(
        MCInst_MC1_v1_3 [2]), .ZN(MCInst_MC1_v1_1 [2]) );
  XNOR2_X1 MCInst_MC1_v1_1Inst_2_U3  ( .A(MCInst_MC1_v1_0 [3]), .B(
        MCInst_MC1_v1_0 [0]), .ZN(MCInst_MC1_v1_1Inst_2_n2 ) );
  XNOR2_X1 MCInst_MC1_v1_2Inst_2_U4  ( .A(MCInst_MC1_v1_2Inst_2_n2 ), .B(
        MCInst_MC1_v1_3 [2]), .ZN(MCInst_MC1_v1_2 [2]) );
  XNOR2_X1 MCInst_MC1_v1_2Inst_2_U3  ( .A(Red_MCInst_MC1_v1_1[0] ), .B(
        MCInst_MC1_v1_0 [0]), .ZN(MCInst_MC1_v1_2Inst_2_n2 ) );
  XNOR2_X1 MCInst_MC1_v2_1Inst_2_U4  ( .A(MCInst_MC1_v2_1Inst_2_n2 ), .B(
        MCInst_MC1_v2_0 [3]), .ZN(MCInst_MC1_v2_1 [2]) );
  XNOR2_X1 MCInst_MC1_v2_1Inst_2_U3  ( .A(MCInst_MC1_v2_0 [0]), .B(
        MCInst_MC1_v2_3 [1]), .ZN(MCInst_MC1_v2_1Inst_2_n2 ) );
  XNOR2_X1 MCInst_MC1_v2_2Inst_2_U4  ( .A(MCInst_MC1_v2_2Inst_2_n2 ), .B(
        MCInst_MC1_v2_0 [3]), .ZN(MCInst_MC1_v2_2 [2]) );
  XNOR2_X1 MCInst_MC1_v2_2Inst_2_U3  ( .A(MCInst_MC1_v2_0 [0]), .B(
        MCInst_MC1_v2_0 [2]), .ZN(MCInst_MC1_v2_2Inst_2_n2 ) );
  XOR2_X1 MCInst_MC1_v2_3Inst_2_U3  ( .A(MCInst_MC1_v2_3 [1]), .B(
        MCInst_MC1_v2_0 [2]), .Z(MCInst_MC1_v2_3 [2]) );
  XNOR2_X1 MCInst_MC1_v3_1Inst_2_U4  ( .A(MCInst_MC1_v3_1Inst_2_n2 ), .B(
        MCInst_MC1_v3_0 [2]), .ZN(MCInst_MC1_v3_1 [2]) );
  XNOR2_X1 MCInst_MC1_v3_1Inst_2_U3  ( .A(MCInst_MC1_v3_2 [2]), .B(
        MCInst_MC1_v3_2 [3]), .ZN(MCInst_MC1_v3_1Inst_2_n2 ) );
  XOR2_X1 MCInst_MC1_v3_3Inst_2_U3  ( .A(MCInst_MC1_v3_0 [2]), .B(
        MCInst_MC1_v3_2 [2]), .Z(MCInst_MC1_v3_3 [2]) );
  XOR2_X1 MCInst_MC1_v0_1Inst_3_U3  ( .A(Red_MCInst_MC1_v0_1[0] ), .B(
        MCInst_MC1_v0_3 [0]), .Z(MCInst_MC1_v0_1 [3]) );
  XOR2_X1 MCInst_MC1_v0_2Inst_3_U3  ( .A(Red_MCInst_MC1_v0_1[0] ), .B(
        MCInst_MC1_v0_3 [3]), .Z(MCInst_MC1_v0_2 [3]) );
  XOR2_X1 MCInst_MC1_v1_1Inst_3_U3  ( .A(MCInst_MC1_v1_3 [2]), .B(
        Red_MCInst_MC1_v1_1[0] ), .Z(MCInst_MC1_v1_1 [3]) );
  XNOR2_X1 MCInst_MC1_v1_2Inst_3_U5  ( .A(MCInst_MC1_v1_2Inst_3_n4 ), .B(
        MCInst_MC1_v1_2Inst_3_n3 ), .ZN(MCInst_MC1_v1_2 [3]) );
  XNOR2_X1 MCInst_MC1_v1_2Inst_3_U4  ( .A(MCInst_MC1_v1_3 [2]), .B(
        MCInst_MC1_v1_0 [0]), .ZN(MCInst_MC1_v1_2Inst_3_n3 ) );
  XOR2_X1 MCInst_MC1_v1_2Inst_3_U3  ( .A(Red_MCInst_MC1_v1_1[0] ), .B(
        MCInst_MC1_v1_0 [3]), .Z(MCInst_MC1_v1_2Inst_3_n4 ) );
  XOR2_X1 MCInst_MC1_v2_1Inst_3_U3  ( .A(MCInst_MC1_v2_0 [2]), .B(
        MCInst_MC1_v2_0 [0]), .Z(MCInst_MC1_v2_1 [3]) );
  XNOR2_X1 MCInst_MC1_v2_2Inst_3_U4  ( .A(MCInst_MC1_v2_2Inst_3_n2 ), .B(
        MCInst_MC1_v2_0 [3]), .ZN(MCInst_MC1_v2_2 [3]) );
  XNOR2_X1 MCInst_MC1_v2_2Inst_3_U3  ( .A(MCInst_MC1_v2_0 [0]), .B(
        MCInst_MC1_v2_3 [1]), .ZN(MCInst_MC1_v2_2Inst_3_n2 ) );
  XNOR2_X1 MCInst_MC1_v2_3Inst_3_U4  ( .A(MCInst_MC1_v2_3Inst_3_n2 ), .B(
        MCInst_MC1_v2_0 [2]), .ZN(MCInst_MC1_v2_3 [3]) );
  XNOR2_X1 MCInst_MC1_v2_3Inst_3_U3  ( .A(MCInst_MC1_v2_0 [3]), .B(
        MCInst_MC1_v2_3 [1]), .ZN(MCInst_MC1_v2_3Inst_3_n2 ) );
  XOR2_X1 MCInst_MC1_v3_1Inst_3_U3  ( .A(MCInst_MC1_v3_0 [2]), .B(
        Red_MCInst_MC1_v3_1[0] ), .Z(MCInst_MC1_v3_1 [3]) );
  XOR2_X1 MCInst_MC1_v3_3Inst_3_U3  ( .A(MCInst_MC1_v3_2 [3]), .B(
        Red_MCInst_MC1_v3_1[0] ), .Z(MCInst_MC1_v3_3 [3]) );
  XNOR2_X1 MCInst_MC1_r0Inst_XORInst_0_0_U3  ( .A(
        MCInst_MC1_r0Inst_XORInst_0_0_n5 ), .B(
        MCInst_MC1_r0Inst_XORInst_0_0_n4 ), .ZN(Feedback[56]) );
  XNOR2_X1 MCInst_MC1_r0Inst_XORInst_0_0_U2  ( .A(MCInst_MC1_v3_2 [2]), .B(
        MCInst_MC1_v2_0 [0]), .ZN(MCInst_MC1_r0Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst_MC1_r0Inst_XORInst_0_0_U1  ( .A(MCInst_MC1_v0_3 [3]), .B(
        MCInst_MC1_v1_0 [0]), .Z(MCInst_MC1_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst_MC1_r0Inst_XORInst_0_1_U3  ( .A(
        MCInst_MC1_r0Inst_XORInst_0_1_n5 ), .B(
        MCInst_MC1_r0Inst_XORInst_0_1_n4 ), .ZN(Feedback[57]) );
  XNOR2_X1 MCInst_MC1_r0Inst_XORInst_0_1_U2  ( .A(MCInst_MC1_v3_0 [1]), .B(
        MCInst_MC1_v2_0 [1]), .ZN(MCInst_MC1_r0Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst_MC1_r0Inst_XORInst_0_1_U1  ( .A(MCInst_MC1_v0_0 [1]), .B(
        MCInst_MC1_v1_3 [2]), .Z(MCInst_MC1_r0Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst_MC1_r0Inst_XORInst_0_2_U3  ( .A(
        MCInst_MC1_r0Inst_XORInst_0_2_n5 ), .B(
        MCInst_MC1_r0Inst_XORInst_0_2_n4 ), .ZN(Feedback[58]) );
  XNOR2_X1 MCInst_MC1_r0Inst_XORInst_0_2_U2  ( .A(MCInst_MC1_v3_0 [2]), .B(
        MCInst_MC1_v2_0 [2]), .ZN(MCInst_MC1_r0Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst_MC1_r0Inst_XORInst_0_2_U1  ( .A(MCInst_MC1_v0_0 [2]), .B(
        Red_MCInst_MC1_v1_1[0] ), .Z(MCInst_MC1_r0Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst_MC1_r0Inst_XORInst_0_3_U3  ( .A(
        MCInst_MC1_r0Inst_XORInst_0_3_n5 ), .B(
        MCInst_MC1_r0Inst_XORInst_0_3_n4 ), .ZN(Feedback[59]) );
  XNOR2_X1 MCInst_MC1_r0Inst_XORInst_0_3_U2  ( .A(Red_MCInst_MC1_v3_1[0] ), 
        .B(MCInst_MC1_v2_0 [3]), .ZN(MCInst_MC1_r0Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst_MC1_r0Inst_XORInst_0_3_U1  ( .A(MCInst_MC1_v0_0 [3]), .B(
        MCInst_MC1_v1_0 [3]), .Z(MCInst_MC1_r0Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst_MC1_r1Inst_XORInst_0_0_U3  ( .A(
        MCInst_MC1_r1Inst_XORInst_0_0_n5 ), .B(
        MCInst_MC1_r1Inst_XORInst_0_0_n4 ), .ZN(Feedback[40]) );
  XNOR2_X1 MCInst_MC1_r1Inst_XORInst_0_0_U2  ( .A(MCInst_MC1_v3_1 [0]), .B(
        MCInst_MC1_v2_1 [0]), .ZN(MCInst_MC1_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst_MC1_r1Inst_XORInst_0_0_U1  ( .A(MCInst_MC1_v0_0 [3]), .B(
        MCInst_MC1_v1_1 [0]), .Z(MCInst_MC1_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst_MC1_r1Inst_XORInst_0_1_U3  ( .A(
        MCInst_MC1_r1Inst_XORInst_0_1_n5 ), .B(
        MCInst_MC1_r1Inst_XORInst_0_1_n4 ), .ZN(Feedback[41]) );
  XNOR2_X1 MCInst_MC1_r1Inst_XORInst_0_1_U2  ( .A(MCInst_MC1_v3_1 [1]), .B(
        MCInst_MC1_v2_1 [1]), .ZN(MCInst_MC1_r1Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst_MC1_r1Inst_XORInst_0_1_U1  ( .A(MCInst_MC1_v0_1 [1]), .B(
        MCInst_MC1_v1_1 [1]), .Z(MCInst_MC1_r1Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst_MC1_r1Inst_XORInst_0_2_U3  ( .A(
        MCInst_MC1_r1Inst_XORInst_0_2_n5 ), .B(
        MCInst_MC1_r1Inst_XORInst_0_2_n4 ), .ZN(Feedback[42]) );
  XNOR2_X1 MCInst_MC1_r1Inst_XORInst_0_2_U2  ( .A(MCInst_MC1_v3_1 [2]), .B(
        MCInst_MC1_v2_1 [2]), .ZN(MCInst_MC1_r1Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst_MC1_r1Inst_XORInst_0_2_U1  ( .A(MCInst_MC1_v0_1 [2]), .B(
        MCInst_MC1_v1_1 [2]), .Z(MCInst_MC1_r1Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst_MC1_r1Inst_XORInst_0_3_U3  ( .A(
        MCInst_MC1_r1Inst_XORInst_0_3_n5 ), .B(
        MCInst_MC1_r1Inst_XORInst_0_3_n4 ), .ZN(Feedback[43]) );
  XNOR2_X1 MCInst_MC1_r1Inst_XORInst_0_3_U2  ( .A(MCInst_MC1_v3_1 [3]), .B(
        MCInst_MC1_v2_1 [3]), .ZN(MCInst_MC1_r1Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst_MC1_r1Inst_XORInst_0_3_U1  ( .A(MCInst_MC1_v0_1 [3]), .B(
        MCInst_MC1_v1_1 [3]), .Z(MCInst_MC1_r1Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst_MC1_r2Inst_XORInst_0_0_U3  ( .A(
        MCInst_MC1_r2Inst_XORInst_0_0_n5 ), .B(
        MCInst_MC1_r2Inst_XORInst_0_0_n4 ), .ZN(Feedback[24]) );
  XNOR2_X1 MCInst_MC1_r2Inst_XORInst_0_0_U2  ( .A(MCInst_MC1_v3_2 [0]), .B(
        MCInst_MC1_v2_2 [0]), .ZN(MCInst_MC1_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst_MC1_r2Inst_XORInst_0_0_U1  ( .A(MCInst_MC1_v0_2 [0]), .B(
        MCInst_MC1_v1_2 [0]), .Z(MCInst_MC1_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst_MC1_r2Inst_XORInst_0_1_U3  ( .A(
        MCInst_MC1_r2Inst_XORInst_0_1_n5 ), .B(
        MCInst_MC1_r2Inst_XORInst_0_1_n4 ), .ZN(Feedback[25]) );
  XNOR2_X1 MCInst_MC1_r2Inst_XORInst_0_1_U2  ( .A(Red_MCInst_MC1_v3_1[0] ), 
        .B(MCInst_MC1_v2_2 [1]), .ZN(MCInst_MC1_r2Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst_MC1_r2Inst_XORInst_0_1_U1  ( .A(MCInst_MC1_v0_2 [1]), .B(
        MCInst_MC1_v1_2 [1]), .Z(MCInst_MC1_r2Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst_MC1_r2Inst_XORInst_0_2_U3  ( .A(
        MCInst_MC1_r2Inst_XORInst_0_2_n5 ), .B(
        MCInst_MC1_r2Inst_XORInst_0_2_n4 ), .ZN(Feedback[26]) );
  XNOR2_X1 MCInst_MC1_r2Inst_XORInst_0_2_U2  ( .A(MCInst_MC1_v3_2 [2]), .B(
        MCInst_MC1_v2_2 [2]), .ZN(MCInst_MC1_r2Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst_MC1_r2Inst_XORInst_0_2_U1  ( .A(MCInst_MC1_v0_2 [2]), .B(
        MCInst_MC1_v1_2 [2]), .Z(MCInst_MC1_r2Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst_MC1_r2Inst_XORInst_0_3_U3  ( .A(
        MCInst_MC1_r2Inst_XORInst_0_3_n5 ), .B(
        MCInst_MC1_r2Inst_XORInst_0_3_n4 ), .ZN(Feedback[27]) );
  XNOR2_X1 MCInst_MC1_r2Inst_XORInst_0_3_U2  ( .A(MCInst_MC1_v3_2 [3]), .B(
        MCInst_MC1_v2_2 [3]), .ZN(MCInst_MC1_r2Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst_MC1_r2Inst_XORInst_0_3_U1  ( .A(MCInst_MC1_v0_2 [3]), .B(
        MCInst_MC1_v1_2 [3]), .Z(MCInst_MC1_r2Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst_MC1_r3Inst_XORInst_0_0_U3  ( .A(
        MCInst_MC1_r3Inst_XORInst_0_0_n5 ), .B(
        MCInst_MC1_r3Inst_XORInst_0_0_n4 ), .ZN(Feedback[8]) );
  XNOR2_X1 MCInst_MC1_r3Inst_XORInst_0_0_U2  ( .A(MCInst_MC1_v3_3 [0]), .B(
        MCInst_MC1_v2_3 [0]), .ZN(MCInst_MC1_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst_MC1_r3Inst_XORInst_0_0_U1  ( .A(MCInst_MC1_v0_3 [0]), .B(
        MCInst_MC1_v1_0 [3]), .Z(MCInst_MC1_r3Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst_MC1_r3Inst_XORInst_0_1_U3  ( .A(
        MCInst_MC1_r3Inst_XORInst_0_1_n5 ), .B(
        MCInst_MC1_r3Inst_XORInst_0_1_n4 ), .ZN(Feedback[9]) );
  XNOR2_X1 MCInst_MC1_r3Inst_XORInst_0_1_U2  ( .A(MCInst_MC1_v3_3 [1]), .B(
        MCInst_MC1_v2_3 [1]), .ZN(MCInst_MC1_r3Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst_MC1_r3Inst_XORInst_0_1_U1  ( .A(MCInst_MC1_v0_3 [1]), .B(
        MCInst_MC1_v1_3 [1]), .Z(MCInst_MC1_r3Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst_MC1_r3Inst_XORInst_0_2_U3  ( .A(
        MCInst_MC1_r3Inst_XORInst_0_2_n5 ), .B(
        MCInst_MC1_r3Inst_XORInst_0_2_n4 ), .ZN(Feedback[10]) );
  XNOR2_X1 MCInst_MC1_r3Inst_XORInst_0_2_U2  ( .A(MCInst_MC1_v3_3 [2]), .B(
        MCInst_MC1_v2_3 [2]), .ZN(MCInst_MC1_r3Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst_MC1_r3Inst_XORInst_0_2_U1  ( .A(MCInst_MC1_v0_0 [3]), .B(
        MCInst_MC1_v1_3 [2]), .Z(MCInst_MC1_r3Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst_MC1_r3Inst_XORInst_0_3_U3  ( .A(
        MCInst_MC1_r3Inst_XORInst_0_3_n5 ), .B(
        MCInst_MC1_r3Inst_XORInst_0_3_n4 ), .ZN(Feedback[11]) );
  XNOR2_X1 MCInst_MC1_r3Inst_XORInst_0_3_U2  ( .A(MCInst_MC1_v3_3 [3]), .B(
        MCInst_MC1_v2_3 [3]), .ZN(MCInst_MC1_r3Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst_MC1_r3Inst_XORInst_0_3_U1  ( .A(MCInst_MC1_v0_3 [3]), .B(
        Red_MCInst_MC1_v1_1[0] ), .Z(MCInst_MC1_r3Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst_MC2_v0_2Inst_0_U4  ( .A(MCInst_MC2_v0_2Inst_0_n2 ), .B(
        MCInst_MC2_v0_0 [3]), .ZN(MCInst_MC2_v0_2 [0]) );
  XNOR2_X1 MCInst_MC2_v0_2Inst_0_U3  ( .A(MCInst_MC2_v0_3 [0]), .B(
        Red_MCInst_MC2_v0_1[0] ), .ZN(MCInst_MC2_v0_2Inst_0_n2 ) );
  XOR2_X1 MCInst_MC2_v1_1Inst_0_U3  ( .A(Red_MCInst_MC2_v1_1[0] ), .B(
        MCInst_MC2_v1_0 [3]), .Z(MCInst_MC2_v1_1 [0]) );
  XNOR2_X1 MCInst_MC2_v1_2Inst_0_U4  ( .A(MCInst_MC2_v1_2Inst_0_n2 ), .B(
        Red_MCInst_MC2_v1_1[0] ), .ZN(MCInst_MC2_v1_2 [0]) );
  XNOR2_X1 MCInst_MC2_v1_2Inst_0_U3  ( .A(MCInst_MC2_v1_0 [3]), .B(
        MCInst_MC2_v1_3 [2]), .ZN(MCInst_MC2_v1_2Inst_0_n2 ) );
  XOR2_X1 MCInst_MC2_v2_1Inst_0_U3  ( .A(MCInst_MC2_v2_3 [1]), .B(
        MCInst_MC2_v2_0 [3]), .Z(MCInst_MC2_v2_1 [0]) );
  XOR2_X1 MCInst_MC2_v2_2Inst_0_U3  ( .A(MCInst_MC2_v2_0 [2]), .B(
        MCInst_MC2_v2_0 [0]), .Z(MCInst_MC2_v2_2 [0]) );
  XNOR2_X1 MCInst_MC2_v2_3Inst_0_U5  ( .A(MCInst_MC2_v2_3Inst_0_n4 ), .B(
        MCInst_MC2_v2_3Inst_0_n3 ), .ZN(MCInst_MC2_v2_3 [0]) );
  XNOR2_X1 MCInst_MC2_v2_3Inst_0_U4  ( .A(MCInst_MC2_v2_0 [2]), .B(
        MCInst_MC2_v2_3 [1]), .ZN(MCInst_MC2_v2_3Inst_0_n3 ) );
  XOR2_X1 MCInst_MC2_v2_3Inst_0_U3  ( .A(MCInst_MC2_v2_0 [3]), .B(
        MCInst_MC2_v2_0 [0]), .Z(MCInst_MC2_v2_3Inst_0_n4 ) );
  XOR2_X1 MCInst_MC2_v3_1Inst_0_U3  ( .A(Red_MCInst_MC2_v3_1[0] ), .B(
        MCInst_MC2_v3_2 [2]), .Z(MCInst_MC2_v3_1 [0]) );
  XOR2_X1 MCInst_MC2_v3_2Inst_0_U3  ( .A(MCInst_MC2_v3_2 [3]), .B(
        MCInst_MC2_v3_0 [2]), .Z(MCInst_MC2_v3_2 [0]) );
  XNOR2_X1 MCInst_MC2_v3_3Inst_0_U4  ( .A(MCInst_MC2_v3_3Inst_0_n2 ), .B(
        MCInst_MC2_v3_0 [2]), .ZN(MCInst_MC2_v3_3 [0]) );
  XNOR2_X1 MCInst_MC2_v3_3Inst_0_U3  ( .A(MCInst_MC2_v3_2 [2]), .B(
        MCInst_MC2_v3_2 [3]), .ZN(MCInst_MC2_v3_3Inst_0_n2 ) );
  XOR2_X1 MCInst_MC2_v0_0Inst_1_U3  ( .A(MCInst_MC2_v0_3 [3]), .B(
        MCInst_MC2_v0_3 [0]), .Z(MCInst_MC2_v0_0 [1]) );
  XOR2_X1 MCInst_MC2_v0_1Inst_1_U3  ( .A(MCInst_MC2_v0_0 [3]), .B(
        MCInst_MC2_v0_3 [3]), .Z(MCInst_MC2_v0_1 [1]) );
  XNOR2_X1 MCInst_MC2_v0_2Inst_1_U4  ( .A(MCInst_MC2_v0_2Inst_1_n2 ), .B(
        MCInst_MC2_v0_3 [3]), .ZN(MCInst_MC2_v0_2 [1]) );
  XNOR2_X1 MCInst_MC2_v0_2Inst_1_U3  ( .A(MCInst_MC2_v0_3 [0]), .B(
        Red_MCInst_MC2_v0_1[0] ), .ZN(MCInst_MC2_v0_2Inst_1_n2 ) );
  XOR2_X1 MCInst_MC2_v0_3Inst_1_U3  ( .A(Red_MCInst_MC2_v0_1[0] ), .B(
        MCInst_MC2_v0_3 [0]), .Z(MCInst_MC2_v0_3 [1]) );
  XOR2_X1 MCInst_MC2_v1_1Inst_1_U3  ( .A(MCInst_MC2_v1_0 [0]), .B(
        Red_MCInst_MC2_v1_1[0] ), .Z(MCInst_MC2_v1_1 [1]) );
  XOR2_X1 MCInst_MC2_v1_2Inst_1_U3  ( .A(MCInst_MC2_v1_0 [0]), .B(
        MCInst_MC2_v1_3 [2]), .Z(MCInst_MC2_v1_2 [1]) );
  XOR2_X1 MCInst_MC2_v1_3Inst_1_U3  ( .A(MCInst_MC2_v1_0 [0]), .B(
        MCInst_MC2_v1_0 [3]), .Z(MCInst_MC2_v1_3 [1]) );
  XOR2_X1 MCInst_MC2_v2_0Inst_1_U3  ( .A(MCInst_MC2_v2_3 [1]), .B(
        MCInst_MC2_v2_0 [0]), .Z(MCInst_MC2_v2_0 [1]) );
  XNOR2_X1 MCInst_MC2_v2_1Inst_1_U4  ( .A(MCInst_MC2_v2_1Inst_1_n2 ), .B(
        MCInst_MC2_v2_0 [3]), .ZN(MCInst_MC2_v2_1 [1]) );
  XNOR2_X1 MCInst_MC2_v2_1Inst_1_U3  ( .A(MCInst_MC2_v2_0 [0]), .B(
        MCInst_MC2_v2_0 [2]), .ZN(MCInst_MC2_v2_1Inst_1_n2 ) );
  XNOR2_X1 MCInst_MC2_v2_2Inst_1_U5  ( .A(MCInst_MC2_v2_2Inst_1_n4 ), .B(
        MCInst_MC2_v2_2Inst_1_n3 ), .ZN(MCInst_MC2_v2_2 [1]) );
  XNOR2_X1 MCInst_MC2_v2_2Inst_1_U4  ( .A(MCInst_MC2_v2_0 [2]), .B(
        MCInst_MC2_v2_3 [1]), .ZN(MCInst_MC2_v2_2Inst_1_n3 ) );
  XOR2_X1 MCInst_MC2_v2_2Inst_1_U3  ( .A(MCInst_MC2_v2_0 [3]), .B(
        MCInst_MC2_v2_0 [0]), .Z(MCInst_MC2_v2_2Inst_1_n4 ) );
  XOR2_X1 MCInst_MC2_v3_0Inst_1_U3  ( .A(MCInst_MC2_v3_2 [3]), .B(
        MCInst_MC2_v3_2 [2]), .Z(MCInst_MC2_v3_0 [1]) );
  XOR2_X1 MCInst_MC2_v3_1Inst_1_U3  ( .A(MCInst_MC2_v3_2 [3]), .B(
        Red_MCInst_MC2_v3_1[0] ), .Z(MCInst_MC2_v3_1 [1]) );
  XNOR2_X1 MCInst_MC2_v3_3Inst_1_U4  ( .A(MCInst_MC2_v3_3Inst_1_n2 ), .B(
        Red_MCInst_MC2_v3_1[0] ), .ZN(MCInst_MC2_v3_3 [1]) );
  XNOR2_X1 MCInst_MC2_v3_3Inst_1_U3  ( .A(MCInst_MC2_v3_2 [2]), .B(
        MCInst_MC2_v3_2 [3]), .ZN(MCInst_MC2_v3_3Inst_1_n2 ) );
  XOR2_X1 MCInst_MC2_v0_0Inst_2_U3  ( .A(Red_MCInst_MC2_v0_1[0] ), .B(
        MCInst_MC2_v0_3 [0]), .Z(MCInst_MC2_v0_0 [2]) );
  XOR2_X1 MCInst_MC2_v0_1Inst_2_U3  ( .A(MCInst_MC2_v0_3 [3]), .B(
        MCInst_MC2_v0_3 [0]), .Z(MCInst_MC2_v0_1 [2]) );
  XOR2_X1 MCInst_MC2_v0_2Inst_2_U3  ( .A(MCInst_MC2_v0_0 [3]), .B(
        MCInst_MC2_v0_3 [0]), .Z(MCInst_MC2_v0_2 [2]) );
  XNOR2_X1 MCInst_MC2_v1_1Inst_2_U4  ( .A(MCInst_MC2_v1_1Inst_2_n2 ), .B(
        MCInst_MC2_v1_3 [2]), .ZN(MCInst_MC2_v1_1 [2]) );
  XNOR2_X1 MCInst_MC2_v1_1Inst_2_U3  ( .A(MCInst_MC2_v1_0 [3]), .B(
        MCInst_MC2_v1_0 [0]), .ZN(MCInst_MC2_v1_1Inst_2_n2 ) );
  XNOR2_X1 MCInst_MC2_v1_2Inst_2_U4  ( .A(MCInst_MC2_v1_2Inst_2_n2 ), .B(
        MCInst_MC2_v1_3 [2]), .ZN(MCInst_MC2_v1_2 [2]) );
  XNOR2_X1 MCInst_MC2_v1_2Inst_2_U3  ( .A(Red_MCInst_MC2_v1_1[0] ), .B(
        MCInst_MC2_v1_0 [0]), .ZN(MCInst_MC2_v1_2Inst_2_n2 ) );
  XNOR2_X1 MCInst_MC2_v2_1Inst_2_U4  ( .A(MCInst_MC2_v2_1Inst_2_n2 ), .B(
        MCInst_MC2_v2_0 [3]), .ZN(MCInst_MC2_v2_1 [2]) );
  XNOR2_X1 MCInst_MC2_v2_1Inst_2_U3  ( .A(MCInst_MC2_v2_0 [0]), .B(
        MCInst_MC2_v2_3 [1]), .ZN(MCInst_MC2_v2_1Inst_2_n2 ) );
  XNOR2_X1 MCInst_MC2_v2_2Inst_2_U4  ( .A(MCInst_MC2_v2_2Inst_2_n2 ), .B(
        MCInst_MC2_v2_0 [3]), .ZN(MCInst_MC2_v2_2 [2]) );
  XNOR2_X1 MCInst_MC2_v2_2Inst_2_U3  ( .A(MCInst_MC2_v2_0 [0]), .B(
        MCInst_MC2_v2_0 [2]), .ZN(MCInst_MC2_v2_2Inst_2_n2 ) );
  XOR2_X1 MCInst_MC2_v2_3Inst_2_U3  ( .A(MCInst_MC2_v2_3 [1]), .B(
        MCInst_MC2_v2_0 [2]), .Z(MCInst_MC2_v2_3 [2]) );
  XNOR2_X1 MCInst_MC2_v3_1Inst_2_U4  ( .A(MCInst_MC2_v3_1Inst_2_n2 ), .B(
        MCInst_MC2_v3_0 [2]), .ZN(MCInst_MC2_v3_1 [2]) );
  XNOR2_X1 MCInst_MC2_v3_1Inst_2_U3  ( .A(MCInst_MC2_v3_2 [2]), .B(
        MCInst_MC2_v3_2 [3]), .ZN(MCInst_MC2_v3_1Inst_2_n2 ) );
  XOR2_X1 MCInst_MC2_v3_3Inst_2_U3  ( .A(MCInst_MC2_v3_0 [2]), .B(
        MCInst_MC2_v3_2 [2]), .Z(MCInst_MC2_v3_3 [2]) );
  XOR2_X1 MCInst_MC2_v0_1Inst_3_U3  ( .A(Red_MCInst_MC2_v0_1[0] ), .B(
        MCInst_MC2_v0_3 [0]), .Z(MCInst_MC2_v0_1 [3]) );
  XOR2_X1 MCInst_MC2_v0_2Inst_3_U3  ( .A(Red_MCInst_MC2_v0_1[0] ), .B(
        MCInst_MC2_v0_3 [3]), .Z(MCInst_MC2_v0_2 [3]) );
  XOR2_X1 MCInst_MC2_v1_1Inst_3_U3  ( .A(MCInst_MC2_v1_3 [2]), .B(
        Red_MCInst_MC2_v1_1[0] ), .Z(MCInst_MC2_v1_1 [3]) );
  XNOR2_X1 MCInst_MC2_v1_2Inst_3_U5  ( .A(MCInst_MC2_v1_2Inst_3_n4 ), .B(
        MCInst_MC2_v1_2Inst_3_n3 ), .ZN(MCInst_MC2_v1_2 [3]) );
  XNOR2_X1 MCInst_MC2_v1_2Inst_3_U4  ( .A(MCInst_MC2_v1_3 [2]), .B(
        MCInst_MC2_v1_0 [0]), .ZN(MCInst_MC2_v1_2Inst_3_n3 ) );
  XOR2_X1 MCInst_MC2_v1_2Inst_3_U3  ( .A(Red_MCInst_MC2_v1_1[0] ), .B(
        MCInst_MC2_v1_0 [3]), .Z(MCInst_MC2_v1_2Inst_3_n4 ) );
  XOR2_X1 MCInst_MC2_v2_1Inst_3_U3  ( .A(MCInst_MC2_v2_0 [2]), .B(
        MCInst_MC2_v2_0 [0]), .Z(MCInst_MC2_v2_1 [3]) );
  XNOR2_X1 MCInst_MC2_v2_2Inst_3_U4  ( .A(MCInst_MC2_v2_2Inst_3_n2 ), .B(
        MCInst_MC2_v2_0 [3]), .ZN(MCInst_MC2_v2_2 [3]) );
  XNOR2_X1 MCInst_MC2_v2_2Inst_3_U3  ( .A(MCInst_MC2_v2_0 [0]), .B(
        MCInst_MC2_v2_3 [1]), .ZN(MCInst_MC2_v2_2Inst_3_n2 ) );
  XNOR2_X1 MCInst_MC2_v2_3Inst_3_U4  ( .A(MCInst_MC2_v2_3Inst_3_n2 ), .B(
        MCInst_MC2_v2_0 [2]), .ZN(MCInst_MC2_v2_3 [3]) );
  XNOR2_X1 MCInst_MC2_v2_3Inst_3_U3  ( .A(MCInst_MC2_v2_0 [3]), .B(
        MCInst_MC2_v2_3 [1]), .ZN(MCInst_MC2_v2_3Inst_3_n2 ) );
  XOR2_X1 MCInst_MC2_v3_1Inst_3_U3  ( .A(MCInst_MC2_v3_0 [2]), .B(
        Red_MCInst_MC2_v3_1[0] ), .Z(MCInst_MC2_v3_1 [3]) );
  XOR2_X1 MCInst_MC2_v3_3Inst_3_U3  ( .A(MCInst_MC2_v3_2 [3]), .B(
        Red_MCInst_MC2_v3_1[0] ), .Z(MCInst_MC2_v3_3 [3]) );
  XNOR2_X1 MCInst_MC2_r0Inst_XORInst_0_0_U3  ( .A(
        MCInst_MC2_r0Inst_XORInst_0_0_n5 ), .B(
        MCInst_MC2_r0Inst_XORInst_0_0_n4 ), .ZN(Feedback[52]) );
  XNOR2_X1 MCInst_MC2_r0Inst_XORInst_0_0_U2  ( .A(MCInst_MC2_v3_2 [2]), .B(
        MCInst_MC2_v2_0 [0]), .ZN(MCInst_MC2_r0Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst_MC2_r0Inst_XORInst_0_0_U1  ( .A(MCInst_MC2_v0_3 [3]), .B(
        MCInst_MC2_v1_0 [0]), .Z(MCInst_MC2_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst_MC2_r0Inst_XORInst_0_1_U3  ( .A(
        MCInst_MC2_r0Inst_XORInst_0_1_n5 ), .B(
        MCInst_MC2_r0Inst_XORInst_0_1_n4 ), .ZN(Feedback[53]) );
  XNOR2_X1 MCInst_MC2_r0Inst_XORInst_0_1_U2  ( .A(MCInst_MC2_v3_0 [1]), .B(
        MCInst_MC2_v2_0 [1]), .ZN(MCInst_MC2_r0Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst_MC2_r0Inst_XORInst_0_1_U1  ( .A(MCInst_MC2_v0_0 [1]), .B(
        MCInst_MC2_v1_3 [2]), .Z(MCInst_MC2_r0Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst_MC2_r0Inst_XORInst_0_2_U3  ( .A(
        MCInst_MC2_r0Inst_XORInst_0_2_n5 ), .B(
        MCInst_MC2_r0Inst_XORInst_0_2_n4 ), .ZN(Feedback[54]) );
  XNOR2_X1 MCInst_MC2_r0Inst_XORInst_0_2_U2  ( .A(MCInst_MC2_v3_0 [2]), .B(
        MCInst_MC2_v2_0 [2]), .ZN(MCInst_MC2_r0Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst_MC2_r0Inst_XORInst_0_2_U1  ( .A(MCInst_MC2_v0_0 [2]), .B(
        Red_MCInst_MC2_v1_1[0] ), .Z(MCInst_MC2_r0Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst_MC2_r0Inst_XORInst_0_3_U3  ( .A(
        MCInst_MC2_r0Inst_XORInst_0_3_n5 ), .B(
        MCInst_MC2_r0Inst_XORInst_0_3_n4 ), .ZN(Feedback[55]) );
  XNOR2_X1 MCInst_MC2_r0Inst_XORInst_0_3_U2  ( .A(Red_MCInst_MC2_v3_1[0] ), 
        .B(MCInst_MC2_v2_0 [3]), .ZN(MCInst_MC2_r0Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst_MC2_r0Inst_XORInst_0_3_U1  ( .A(MCInst_MC2_v0_0 [3]), .B(
        MCInst_MC2_v1_0 [3]), .Z(MCInst_MC2_r0Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst_MC2_r1Inst_XORInst_0_0_U3  ( .A(
        MCInst_MC2_r1Inst_XORInst_0_0_n5 ), .B(
        MCInst_MC2_r1Inst_XORInst_0_0_n4 ), .ZN(Feedback[36]) );
  XNOR2_X1 MCInst_MC2_r1Inst_XORInst_0_0_U2  ( .A(MCInst_MC2_v3_1 [0]), .B(
        MCInst_MC2_v2_1 [0]), .ZN(MCInst_MC2_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst_MC2_r1Inst_XORInst_0_0_U1  ( .A(MCInst_MC2_v0_0 [3]), .B(
        MCInst_MC2_v1_1 [0]), .Z(MCInst_MC2_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst_MC2_r1Inst_XORInst_0_1_U3  ( .A(
        MCInst_MC2_r1Inst_XORInst_0_1_n5 ), .B(
        MCInst_MC2_r1Inst_XORInst_0_1_n4 ), .ZN(Feedback[37]) );
  XNOR2_X1 MCInst_MC2_r1Inst_XORInst_0_1_U2  ( .A(MCInst_MC2_v3_1 [1]), .B(
        MCInst_MC2_v2_1 [1]), .ZN(MCInst_MC2_r1Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst_MC2_r1Inst_XORInst_0_1_U1  ( .A(MCInst_MC2_v0_1 [1]), .B(
        MCInst_MC2_v1_1 [1]), .Z(MCInst_MC2_r1Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst_MC2_r1Inst_XORInst_0_2_U3  ( .A(
        MCInst_MC2_r1Inst_XORInst_0_2_n5 ), .B(
        MCInst_MC2_r1Inst_XORInst_0_2_n4 ), .ZN(Feedback[38]) );
  XNOR2_X1 MCInst_MC2_r1Inst_XORInst_0_2_U2  ( .A(MCInst_MC2_v3_1 [2]), .B(
        MCInst_MC2_v2_1 [2]), .ZN(MCInst_MC2_r1Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst_MC2_r1Inst_XORInst_0_2_U1  ( .A(MCInst_MC2_v0_1 [2]), .B(
        MCInst_MC2_v1_1 [2]), .Z(MCInst_MC2_r1Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst_MC2_r1Inst_XORInst_0_3_U3  ( .A(
        MCInst_MC2_r1Inst_XORInst_0_3_n5 ), .B(
        MCInst_MC2_r1Inst_XORInst_0_3_n4 ), .ZN(Feedback[39]) );
  XNOR2_X1 MCInst_MC2_r1Inst_XORInst_0_3_U2  ( .A(MCInst_MC2_v3_1 [3]), .B(
        MCInst_MC2_v2_1 [3]), .ZN(MCInst_MC2_r1Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst_MC2_r1Inst_XORInst_0_3_U1  ( .A(MCInst_MC2_v0_1 [3]), .B(
        MCInst_MC2_v1_1 [3]), .Z(MCInst_MC2_r1Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst_MC2_r2Inst_XORInst_0_0_U3  ( .A(
        MCInst_MC2_r2Inst_XORInst_0_0_n5 ), .B(
        MCInst_MC2_r2Inst_XORInst_0_0_n4 ), .ZN(Feedback[20]) );
  XNOR2_X1 MCInst_MC2_r2Inst_XORInst_0_0_U2  ( .A(MCInst_MC2_v3_2 [0]), .B(
        MCInst_MC2_v2_2 [0]), .ZN(MCInst_MC2_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst_MC2_r2Inst_XORInst_0_0_U1  ( .A(MCInst_MC2_v0_2 [0]), .B(
        MCInst_MC2_v1_2 [0]), .Z(MCInst_MC2_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst_MC2_r2Inst_XORInst_0_1_U3  ( .A(
        MCInst_MC2_r2Inst_XORInst_0_1_n5 ), .B(
        MCInst_MC2_r2Inst_XORInst_0_1_n4 ), .ZN(Feedback[21]) );
  XNOR2_X1 MCInst_MC2_r2Inst_XORInst_0_1_U2  ( .A(Red_MCInst_MC2_v3_1[0] ), 
        .B(MCInst_MC2_v2_2 [1]), .ZN(MCInst_MC2_r2Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst_MC2_r2Inst_XORInst_0_1_U1  ( .A(MCInst_MC2_v0_2 [1]), .B(
        MCInst_MC2_v1_2 [1]), .Z(MCInst_MC2_r2Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst_MC2_r2Inst_XORInst_0_2_U3  ( .A(
        MCInst_MC2_r2Inst_XORInst_0_2_n5 ), .B(
        MCInst_MC2_r2Inst_XORInst_0_2_n4 ), .ZN(Feedback[22]) );
  XNOR2_X1 MCInst_MC2_r2Inst_XORInst_0_2_U2  ( .A(MCInst_MC2_v3_2 [2]), .B(
        MCInst_MC2_v2_2 [2]), .ZN(MCInst_MC2_r2Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst_MC2_r2Inst_XORInst_0_2_U1  ( .A(MCInst_MC2_v0_2 [2]), .B(
        MCInst_MC2_v1_2 [2]), .Z(MCInst_MC2_r2Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst_MC2_r2Inst_XORInst_0_3_U3  ( .A(
        MCInst_MC2_r2Inst_XORInst_0_3_n5 ), .B(
        MCInst_MC2_r2Inst_XORInst_0_3_n4 ), .ZN(Feedback[23]) );
  XNOR2_X1 MCInst_MC2_r2Inst_XORInst_0_3_U2  ( .A(MCInst_MC2_v3_2 [3]), .B(
        MCInst_MC2_v2_2 [3]), .ZN(MCInst_MC2_r2Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst_MC2_r2Inst_XORInst_0_3_U1  ( .A(MCInst_MC2_v0_2 [3]), .B(
        MCInst_MC2_v1_2 [3]), .Z(MCInst_MC2_r2Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst_MC2_r3Inst_XORInst_0_0_U3  ( .A(
        MCInst_MC2_r3Inst_XORInst_0_0_n5 ), .B(
        MCInst_MC2_r3Inst_XORInst_0_0_n4 ), .ZN(Feedback[4]) );
  XNOR2_X1 MCInst_MC2_r3Inst_XORInst_0_0_U2  ( .A(MCInst_MC2_v3_3 [0]), .B(
        MCInst_MC2_v2_3 [0]), .ZN(MCInst_MC2_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst_MC2_r3Inst_XORInst_0_0_U1  ( .A(MCInst_MC2_v0_3 [0]), .B(
        MCInst_MC2_v1_0 [3]), .Z(MCInst_MC2_r3Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst_MC2_r3Inst_XORInst_0_1_U3  ( .A(
        MCInst_MC2_r3Inst_XORInst_0_1_n5 ), .B(
        MCInst_MC2_r3Inst_XORInst_0_1_n4 ), .ZN(Feedback[5]) );
  XNOR2_X1 MCInst_MC2_r3Inst_XORInst_0_1_U2  ( .A(MCInst_MC2_v3_3 [1]), .B(
        MCInst_MC2_v2_3 [1]), .ZN(MCInst_MC2_r3Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst_MC2_r3Inst_XORInst_0_1_U1  ( .A(MCInst_MC2_v0_3 [1]), .B(
        MCInst_MC2_v1_3 [1]), .Z(MCInst_MC2_r3Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst_MC2_r3Inst_XORInst_0_2_U3  ( .A(
        MCInst_MC2_r3Inst_XORInst_0_2_n5 ), .B(
        MCInst_MC2_r3Inst_XORInst_0_2_n4 ), .ZN(Feedback[6]) );
  XNOR2_X1 MCInst_MC2_r3Inst_XORInst_0_2_U2  ( .A(MCInst_MC2_v3_3 [2]), .B(
        MCInst_MC2_v2_3 [2]), .ZN(MCInst_MC2_r3Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst_MC2_r3Inst_XORInst_0_2_U1  ( .A(MCInst_MC2_v0_0 [3]), .B(
        MCInst_MC2_v1_3 [2]), .Z(MCInst_MC2_r3Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst_MC2_r3Inst_XORInst_0_3_U3  ( .A(
        MCInst_MC2_r3Inst_XORInst_0_3_n5 ), .B(
        MCInst_MC2_r3Inst_XORInst_0_3_n4 ), .ZN(Feedback[7]) );
  XNOR2_X1 MCInst_MC2_r3Inst_XORInst_0_3_U2  ( .A(MCInst_MC2_v3_3 [3]), .B(
        MCInst_MC2_v2_3 [3]), .ZN(MCInst_MC2_r3Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst_MC2_r3Inst_XORInst_0_3_U1  ( .A(MCInst_MC2_v0_3 [3]), .B(
        Red_MCInst_MC2_v1_1[0] ), .Z(MCInst_MC2_r3Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst_MC3_v0_2Inst_0_U4  ( .A(MCInst_MC3_v0_2Inst_0_n2 ), .B(
        MCInst_MC3_v0_0 [3]), .ZN(MCInst_MC3_v0_2 [0]) );
  XNOR2_X1 MCInst_MC3_v0_2Inst_0_U3  ( .A(MCInst_MC3_v0_3 [0]), .B(
        Red_MCInst_MC3_v0_1[0] ), .ZN(MCInst_MC3_v0_2Inst_0_n2 ) );
  XOR2_X1 MCInst_MC3_v1_1Inst_0_U3  ( .A(Red_MCInst_MC3_v1_1[0] ), .B(
        MCInst_MC3_v1_0 [3]), .Z(MCInst_MC3_v1_1 [0]) );
  XNOR2_X1 MCInst_MC3_v1_2Inst_0_U4  ( .A(MCInst_MC3_v1_2Inst_0_n2 ), .B(
        Red_MCInst_MC3_v1_1[0] ), .ZN(MCInst_MC3_v1_2 [0]) );
  XNOR2_X1 MCInst_MC3_v1_2Inst_0_U3  ( .A(MCInst_MC3_v1_0 [3]), .B(
        MCInst_MC3_v1_3 [2]), .ZN(MCInst_MC3_v1_2Inst_0_n2 ) );
  XOR2_X1 MCInst_MC3_v2_1Inst_0_U3  ( .A(MCInst_MC3_v2_3 [1]), .B(
        MCInst_MC3_v2_0 [3]), .Z(MCInst_MC3_v2_1 [0]) );
  XOR2_X1 MCInst_MC3_v2_2Inst_0_U3  ( .A(MCInst_MC3_v2_0 [2]), .B(
        MCInst_MC3_v2_0 [0]), .Z(MCInst_MC3_v2_2 [0]) );
  XNOR2_X1 MCInst_MC3_v2_3Inst_0_U5  ( .A(MCInst_MC3_v2_3Inst_0_n4 ), .B(
        MCInst_MC3_v2_3Inst_0_n3 ), .ZN(MCInst_MC3_v2_3 [0]) );
  XNOR2_X1 MCInst_MC3_v2_3Inst_0_U4  ( .A(MCInst_MC3_v2_0 [2]), .B(
        MCInst_MC3_v2_3 [1]), .ZN(MCInst_MC3_v2_3Inst_0_n3 ) );
  XOR2_X1 MCInst_MC3_v2_3Inst_0_U3  ( .A(MCInst_MC3_v2_0 [3]), .B(
        MCInst_MC3_v2_0 [0]), .Z(MCInst_MC3_v2_3Inst_0_n4 ) );
  XOR2_X1 MCInst_MC3_v3_1Inst_0_U3  ( .A(Red_MCInst_MC3_v3_1[0] ), .B(
        MCInst_MC3_v3_2 [2]), .Z(MCInst_MC3_v3_1 [0]) );
  XOR2_X1 MCInst_MC3_v3_2Inst_0_U3  ( .A(MCInst_MC3_v3_2 [3]), .B(
        MCInst_MC3_v3_0 [2]), .Z(MCInst_MC3_v3_2 [0]) );
  XNOR2_X1 MCInst_MC3_v3_3Inst_0_U4  ( .A(MCInst_MC3_v3_3Inst_0_n2 ), .B(
        MCInst_MC3_v3_0 [2]), .ZN(MCInst_MC3_v3_3 [0]) );
  XNOR2_X1 MCInst_MC3_v3_3Inst_0_U3  ( .A(MCInst_MC3_v3_2 [2]), .B(
        MCInst_MC3_v3_2 [3]), .ZN(MCInst_MC3_v3_3Inst_0_n2 ) );
  XOR2_X1 MCInst_MC3_v0_0Inst_1_U3  ( .A(MCInst_MC3_v0_3 [3]), .B(
        MCInst_MC3_v0_3 [0]), .Z(MCInst_MC3_v0_0 [1]) );
  XOR2_X1 MCInst_MC3_v0_1Inst_1_U3  ( .A(MCInst_MC3_v0_0 [3]), .B(
        MCInst_MC3_v0_3 [3]), .Z(MCInst_MC3_v0_1 [1]) );
  XNOR2_X1 MCInst_MC3_v0_2Inst_1_U4  ( .A(MCInst_MC3_v0_2Inst_1_n2 ), .B(
        MCInst_MC3_v0_3 [3]), .ZN(MCInst_MC3_v0_2 [1]) );
  XNOR2_X1 MCInst_MC3_v0_2Inst_1_U3  ( .A(MCInst_MC3_v0_3 [0]), .B(
        Red_MCInst_MC3_v0_1[0] ), .ZN(MCInst_MC3_v0_2Inst_1_n2 ) );
  XOR2_X1 MCInst_MC3_v0_3Inst_1_U3  ( .A(Red_MCInst_MC3_v0_1[0] ), .B(
        MCInst_MC3_v0_3 [0]), .Z(MCInst_MC3_v0_3 [1]) );
  XOR2_X1 MCInst_MC3_v1_1Inst_1_U3  ( .A(MCInst_MC3_v1_0 [0]), .B(
        Red_MCInst_MC3_v1_1[0] ), .Z(MCInst_MC3_v1_1 [1]) );
  XOR2_X1 MCInst_MC3_v1_2Inst_1_U3  ( .A(MCInst_MC3_v1_0 [0]), .B(
        MCInst_MC3_v1_3 [2]), .Z(MCInst_MC3_v1_2 [1]) );
  XOR2_X1 MCInst_MC3_v1_3Inst_1_U3  ( .A(MCInst_MC3_v1_0 [0]), .B(
        MCInst_MC3_v1_0 [3]), .Z(MCInst_MC3_v1_3 [1]) );
  XOR2_X1 MCInst_MC3_v2_0Inst_1_U3  ( .A(MCInst_MC3_v2_3 [1]), .B(
        MCInst_MC3_v2_0 [0]), .Z(MCInst_MC3_v2_0 [1]) );
  XNOR2_X1 MCInst_MC3_v2_1Inst_1_U4  ( .A(MCInst_MC3_v2_1Inst_1_n2 ), .B(
        MCInst_MC3_v2_0 [3]), .ZN(MCInst_MC3_v2_1 [1]) );
  XNOR2_X1 MCInst_MC3_v2_1Inst_1_U3  ( .A(MCInst_MC3_v2_0 [0]), .B(
        MCInst_MC3_v2_0 [2]), .ZN(MCInst_MC3_v2_1Inst_1_n2 ) );
  XNOR2_X1 MCInst_MC3_v2_2Inst_1_U5  ( .A(MCInst_MC3_v2_2Inst_1_n4 ), .B(
        MCInst_MC3_v2_2Inst_1_n3 ), .ZN(MCInst_MC3_v2_2 [1]) );
  XNOR2_X1 MCInst_MC3_v2_2Inst_1_U4  ( .A(MCInst_MC3_v2_0 [2]), .B(
        MCInst_MC3_v2_3 [1]), .ZN(MCInst_MC3_v2_2Inst_1_n3 ) );
  XOR2_X1 MCInst_MC3_v2_2Inst_1_U3  ( .A(MCInst_MC3_v2_0 [3]), .B(
        MCInst_MC3_v2_0 [0]), .Z(MCInst_MC3_v2_2Inst_1_n4 ) );
  XOR2_X1 MCInst_MC3_v3_0Inst_1_U3  ( .A(MCInst_MC3_v3_2 [3]), .B(
        MCInst_MC3_v3_2 [2]), .Z(MCInst_MC3_v3_0 [1]) );
  XOR2_X1 MCInst_MC3_v3_1Inst_1_U3  ( .A(MCInst_MC3_v3_2 [3]), .B(
        Red_MCInst_MC3_v3_1[0] ), .Z(MCInst_MC3_v3_1 [1]) );
  XNOR2_X1 MCInst_MC3_v3_3Inst_1_U4  ( .A(MCInst_MC3_v3_3Inst_1_n2 ), .B(
        Red_MCInst_MC3_v3_1[0] ), .ZN(MCInst_MC3_v3_3 [1]) );
  XNOR2_X1 MCInst_MC3_v3_3Inst_1_U3  ( .A(MCInst_MC3_v3_2 [2]), .B(
        MCInst_MC3_v3_2 [3]), .ZN(MCInst_MC3_v3_3Inst_1_n2 ) );
  XOR2_X1 MCInst_MC3_v0_0Inst_2_U3  ( .A(Red_MCInst_MC3_v0_1[0] ), .B(
        MCInst_MC3_v0_3 [0]), .Z(MCInst_MC3_v0_0 [2]) );
  XOR2_X1 MCInst_MC3_v0_1Inst_2_U3  ( .A(MCInst_MC3_v0_3 [3]), .B(
        MCInst_MC3_v0_3 [0]), .Z(MCInst_MC3_v0_1 [2]) );
  XOR2_X1 MCInst_MC3_v0_2Inst_2_U3  ( .A(MCInst_MC3_v0_0 [3]), .B(
        MCInst_MC3_v0_3 [0]), .Z(MCInst_MC3_v0_2 [2]) );
  XNOR2_X1 MCInst_MC3_v1_1Inst_2_U4  ( .A(MCInst_MC3_v1_1Inst_2_n2 ), .B(
        MCInst_MC3_v1_3 [2]), .ZN(MCInst_MC3_v1_1 [2]) );
  XNOR2_X1 MCInst_MC3_v1_1Inst_2_U3  ( .A(MCInst_MC3_v1_0 [3]), .B(
        MCInst_MC3_v1_0 [0]), .ZN(MCInst_MC3_v1_1Inst_2_n2 ) );
  XNOR2_X1 MCInst_MC3_v1_2Inst_2_U4  ( .A(MCInst_MC3_v1_2Inst_2_n2 ), .B(
        MCInst_MC3_v1_3 [2]), .ZN(MCInst_MC3_v1_2 [2]) );
  XNOR2_X1 MCInst_MC3_v1_2Inst_2_U3  ( .A(Red_MCInst_MC3_v1_1[0] ), .B(
        MCInst_MC3_v1_0 [0]), .ZN(MCInst_MC3_v1_2Inst_2_n2 ) );
  XNOR2_X1 MCInst_MC3_v2_1Inst_2_U4  ( .A(MCInst_MC3_v2_1Inst_2_n2 ), .B(
        MCInst_MC3_v2_0 [3]), .ZN(MCInst_MC3_v2_1 [2]) );
  XNOR2_X1 MCInst_MC3_v2_1Inst_2_U3  ( .A(MCInst_MC3_v2_0 [0]), .B(
        MCInst_MC3_v2_3 [1]), .ZN(MCInst_MC3_v2_1Inst_2_n2 ) );
  XNOR2_X1 MCInst_MC3_v2_2Inst_2_U4  ( .A(MCInst_MC3_v2_2Inst_2_n2 ), .B(
        MCInst_MC3_v2_0 [3]), .ZN(MCInst_MC3_v2_2 [2]) );
  XNOR2_X1 MCInst_MC3_v2_2Inst_2_U3  ( .A(MCInst_MC3_v2_0 [0]), .B(
        MCInst_MC3_v2_0 [2]), .ZN(MCInst_MC3_v2_2Inst_2_n2 ) );
  XOR2_X1 MCInst_MC3_v2_3Inst_2_U3  ( .A(MCInst_MC3_v2_3 [1]), .B(
        MCInst_MC3_v2_0 [2]), .Z(MCInst_MC3_v2_3 [2]) );
  XNOR2_X1 MCInst_MC3_v3_1Inst_2_U4  ( .A(MCInst_MC3_v3_1Inst_2_n2 ), .B(
        MCInst_MC3_v3_0 [2]), .ZN(MCInst_MC3_v3_1 [2]) );
  XNOR2_X1 MCInst_MC3_v3_1Inst_2_U3  ( .A(MCInst_MC3_v3_2 [2]), .B(
        MCInst_MC3_v3_2 [3]), .ZN(MCInst_MC3_v3_1Inst_2_n2 ) );
  XOR2_X1 MCInst_MC3_v3_3Inst_2_U3  ( .A(MCInst_MC3_v3_0 [2]), .B(
        MCInst_MC3_v3_2 [2]), .Z(MCInst_MC3_v3_3 [2]) );
  XOR2_X1 MCInst_MC3_v0_1Inst_3_U3  ( .A(Red_MCInst_MC3_v0_1[0] ), .B(
        MCInst_MC3_v0_3 [0]), .Z(MCInst_MC3_v0_1 [3]) );
  XOR2_X1 MCInst_MC3_v0_2Inst_3_U3  ( .A(Red_MCInst_MC3_v0_1[0] ), .B(
        MCInst_MC3_v0_3 [3]), .Z(MCInst_MC3_v0_2 [3]) );
  XOR2_X1 MCInst_MC3_v1_1Inst_3_U3  ( .A(MCInst_MC3_v1_3 [2]), .B(
        Red_MCInst_MC3_v1_1[0] ), .Z(MCInst_MC3_v1_1 [3]) );
  XNOR2_X1 MCInst_MC3_v1_2Inst_3_U5  ( .A(MCInst_MC3_v1_2Inst_3_n4 ), .B(
        MCInst_MC3_v1_2Inst_3_n3 ), .ZN(MCInst_MC3_v1_2 [3]) );
  XNOR2_X1 MCInst_MC3_v1_2Inst_3_U4  ( .A(MCInst_MC3_v1_3 [2]), .B(
        MCInst_MC3_v1_0 [0]), .ZN(MCInst_MC3_v1_2Inst_3_n3 ) );
  XOR2_X1 MCInst_MC3_v1_2Inst_3_U3  ( .A(Red_MCInst_MC3_v1_1[0] ), .B(
        MCInst_MC3_v1_0 [3]), .Z(MCInst_MC3_v1_2Inst_3_n4 ) );
  XOR2_X1 MCInst_MC3_v2_1Inst_3_U3  ( .A(MCInst_MC3_v2_0 [2]), .B(
        MCInst_MC3_v2_0 [0]), .Z(MCInst_MC3_v2_1 [3]) );
  XNOR2_X1 MCInst_MC3_v2_2Inst_3_U4  ( .A(MCInst_MC3_v2_2Inst_3_n2 ), .B(
        MCInst_MC3_v2_0 [3]), .ZN(MCInst_MC3_v2_2 [3]) );
  XNOR2_X1 MCInst_MC3_v2_2Inst_3_U3  ( .A(MCInst_MC3_v2_0 [0]), .B(
        MCInst_MC3_v2_3 [1]), .ZN(MCInst_MC3_v2_2Inst_3_n2 ) );
  XNOR2_X1 MCInst_MC3_v2_3Inst_3_U4  ( .A(MCInst_MC3_v2_3Inst_3_n2 ), .B(
        MCInst_MC3_v2_0 [2]), .ZN(MCInst_MC3_v2_3 [3]) );
  XNOR2_X1 MCInst_MC3_v2_3Inst_3_U3  ( .A(MCInst_MC3_v2_0 [3]), .B(
        MCInst_MC3_v2_3 [1]), .ZN(MCInst_MC3_v2_3Inst_3_n2 ) );
  XOR2_X1 MCInst_MC3_v3_1Inst_3_U3  ( .A(MCInst_MC3_v3_0 [2]), .B(
        Red_MCInst_MC3_v3_1[0] ), .Z(MCInst_MC3_v3_1 [3]) );
  XOR2_X1 MCInst_MC3_v3_3Inst_3_U3  ( .A(MCInst_MC3_v3_2 [3]), .B(
        Red_MCInst_MC3_v3_1[0] ), .Z(MCInst_MC3_v3_3 [3]) );
  XNOR2_X1 MCInst_MC3_r0Inst_XORInst_0_0_U3  ( .A(
        MCInst_MC3_r0Inst_XORInst_0_0_n5 ), .B(
        MCInst_MC3_r0Inst_XORInst_0_0_n4 ), .ZN(Feedback[48]) );
  XNOR2_X1 MCInst_MC3_r0Inst_XORInst_0_0_U2  ( .A(MCInst_MC3_v3_2 [2]), .B(
        MCInst_MC3_v2_0 [0]), .ZN(MCInst_MC3_r0Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst_MC3_r0Inst_XORInst_0_0_U1  ( .A(MCInst_MC3_v0_3 [3]), .B(
        MCInst_MC3_v1_0 [0]), .Z(MCInst_MC3_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst_MC3_r0Inst_XORInst_0_1_U3  ( .A(
        MCInst_MC3_r0Inst_XORInst_0_1_n5 ), .B(
        MCInst_MC3_r0Inst_XORInst_0_1_n4 ), .ZN(Feedback[49]) );
  XNOR2_X1 MCInst_MC3_r0Inst_XORInst_0_1_U2  ( .A(MCInst_MC3_v3_0 [1]), .B(
        MCInst_MC3_v2_0 [1]), .ZN(MCInst_MC3_r0Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst_MC3_r0Inst_XORInst_0_1_U1  ( .A(MCInst_MC3_v0_0 [1]), .B(
        MCInst_MC3_v1_3 [2]), .Z(MCInst_MC3_r0Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst_MC3_r0Inst_XORInst_0_2_U3  ( .A(
        MCInst_MC3_r0Inst_XORInst_0_2_n5 ), .B(
        MCInst_MC3_r0Inst_XORInst_0_2_n4 ), .ZN(Feedback[50]) );
  XNOR2_X1 MCInst_MC3_r0Inst_XORInst_0_2_U2  ( .A(MCInst_MC3_v3_0 [2]), .B(
        MCInst_MC3_v2_0 [2]), .ZN(MCInst_MC3_r0Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst_MC3_r0Inst_XORInst_0_2_U1  ( .A(MCInst_MC3_v0_0 [2]), .B(
        Red_MCInst_MC3_v1_1[0] ), .Z(MCInst_MC3_r0Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst_MC3_r0Inst_XORInst_0_3_U3  ( .A(
        MCInst_MC3_r0Inst_XORInst_0_3_n5 ), .B(
        MCInst_MC3_r0Inst_XORInst_0_3_n4 ), .ZN(Feedback[51]) );
  XNOR2_X1 MCInst_MC3_r0Inst_XORInst_0_3_U2  ( .A(Red_MCInst_MC3_v3_1[0] ), 
        .B(MCInst_MC3_v2_0 [3]), .ZN(MCInst_MC3_r0Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst_MC3_r0Inst_XORInst_0_3_U1  ( .A(MCInst_MC3_v0_0 [3]), .B(
        MCInst_MC3_v1_0 [3]), .Z(MCInst_MC3_r0Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst_MC3_r1Inst_XORInst_0_0_U3  ( .A(
        MCInst_MC3_r1Inst_XORInst_0_0_n5 ), .B(
        MCInst_MC3_r1Inst_XORInst_0_0_n4 ), .ZN(Feedback[32]) );
  XNOR2_X1 MCInst_MC3_r1Inst_XORInst_0_0_U2  ( .A(MCInst_MC3_v3_1 [0]), .B(
        MCInst_MC3_v2_1 [0]), .ZN(MCInst_MC3_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst_MC3_r1Inst_XORInst_0_0_U1  ( .A(MCInst_MC3_v0_0 [3]), .B(
        MCInst_MC3_v1_1 [0]), .Z(MCInst_MC3_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst_MC3_r1Inst_XORInst_0_1_U3  ( .A(
        MCInst_MC3_r1Inst_XORInst_0_1_n5 ), .B(
        MCInst_MC3_r1Inst_XORInst_0_1_n4 ), .ZN(Feedback[33]) );
  XNOR2_X1 MCInst_MC3_r1Inst_XORInst_0_1_U2  ( .A(MCInst_MC3_v3_1 [1]), .B(
        MCInst_MC3_v2_1 [1]), .ZN(MCInst_MC3_r1Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst_MC3_r1Inst_XORInst_0_1_U1  ( .A(MCInst_MC3_v0_1 [1]), .B(
        MCInst_MC3_v1_1 [1]), .Z(MCInst_MC3_r1Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst_MC3_r1Inst_XORInst_0_2_U3  ( .A(
        MCInst_MC3_r1Inst_XORInst_0_2_n5 ), .B(
        MCInst_MC3_r1Inst_XORInst_0_2_n4 ), .ZN(Feedback[34]) );
  XNOR2_X1 MCInst_MC3_r1Inst_XORInst_0_2_U2  ( .A(MCInst_MC3_v3_1 [2]), .B(
        MCInst_MC3_v2_1 [2]), .ZN(MCInst_MC3_r1Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst_MC3_r1Inst_XORInst_0_2_U1  ( .A(MCInst_MC3_v0_1 [2]), .B(
        MCInst_MC3_v1_1 [2]), .Z(MCInst_MC3_r1Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst_MC3_r1Inst_XORInst_0_3_U3  ( .A(
        MCInst_MC3_r1Inst_XORInst_0_3_n5 ), .B(
        MCInst_MC3_r1Inst_XORInst_0_3_n4 ), .ZN(Feedback[35]) );
  XNOR2_X1 MCInst_MC3_r1Inst_XORInst_0_3_U2  ( .A(MCInst_MC3_v3_1 [3]), .B(
        MCInst_MC3_v2_1 [3]), .ZN(MCInst_MC3_r1Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst_MC3_r1Inst_XORInst_0_3_U1  ( .A(MCInst_MC3_v0_1 [3]), .B(
        MCInst_MC3_v1_1 [3]), .Z(MCInst_MC3_r1Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst_MC3_r2Inst_XORInst_0_0_U3  ( .A(
        MCInst_MC3_r2Inst_XORInst_0_0_n5 ), .B(
        MCInst_MC3_r2Inst_XORInst_0_0_n4 ), .ZN(Feedback[16]) );
  XNOR2_X1 MCInst_MC3_r2Inst_XORInst_0_0_U2  ( .A(MCInst_MC3_v3_2 [0]), .B(
        MCInst_MC3_v2_2 [0]), .ZN(MCInst_MC3_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst_MC3_r2Inst_XORInst_0_0_U1  ( .A(MCInst_MC3_v0_2 [0]), .B(
        MCInst_MC3_v1_2 [0]), .Z(MCInst_MC3_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst_MC3_r2Inst_XORInst_0_1_U3  ( .A(
        MCInst_MC3_r2Inst_XORInst_0_1_n5 ), .B(
        MCInst_MC3_r2Inst_XORInst_0_1_n4 ), .ZN(Feedback[17]) );
  XNOR2_X1 MCInst_MC3_r2Inst_XORInst_0_1_U2  ( .A(Red_MCInst_MC3_v3_1[0] ), 
        .B(MCInst_MC3_v2_2 [1]), .ZN(MCInst_MC3_r2Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst_MC3_r2Inst_XORInst_0_1_U1  ( .A(MCInst_MC3_v0_2 [1]), .B(
        MCInst_MC3_v1_2 [1]), .Z(MCInst_MC3_r2Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst_MC3_r2Inst_XORInst_0_2_U3  ( .A(
        MCInst_MC3_r2Inst_XORInst_0_2_n5 ), .B(
        MCInst_MC3_r2Inst_XORInst_0_2_n4 ), .ZN(Feedback[18]) );
  XNOR2_X1 MCInst_MC3_r2Inst_XORInst_0_2_U2  ( .A(MCInst_MC3_v3_2 [2]), .B(
        MCInst_MC3_v2_2 [2]), .ZN(MCInst_MC3_r2Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst_MC3_r2Inst_XORInst_0_2_U1  ( .A(MCInst_MC3_v0_2 [2]), .B(
        MCInst_MC3_v1_2 [2]), .Z(MCInst_MC3_r2Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst_MC3_r2Inst_XORInst_0_3_U3  ( .A(
        MCInst_MC3_r2Inst_XORInst_0_3_n5 ), .B(
        MCInst_MC3_r2Inst_XORInst_0_3_n4 ), .ZN(Feedback[19]) );
  XNOR2_X1 MCInst_MC3_r2Inst_XORInst_0_3_U2  ( .A(MCInst_MC3_v3_2 [3]), .B(
        MCInst_MC3_v2_2 [3]), .ZN(MCInst_MC3_r2Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst_MC3_r2Inst_XORInst_0_3_U1  ( .A(MCInst_MC3_v0_2 [3]), .B(
        MCInst_MC3_v1_2 [3]), .Z(MCInst_MC3_r2Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst_MC3_r3Inst_XORInst_0_0_U3  ( .A(
        MCInst_MC3_r3Inst_XORInst_0_0_n5 ), .B(
        MCInst_MC3_r3Inst_XORInst_0_0_n4 ), .ZN(Feedback[0]) );
  XNOR2_X1 MCInst_MC3_r3Inst_XORInst_0_0_U2  ( .A(MCInst_MC3_v3_3 [0]), .B(
        MCInst_MC3_v2_3 [0]), .ZN(MCInst_MC3_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst_MC3_r3Inst_XORInst_0_0_U1  ( .A(MCInst_MC3_v0_3 [0]), .B(
        MCInst_MC3_v1_0 [3]), .Z(MCInst_MC3_r3Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst_MC3_r3Inst_XORInst_0_1_U3  ( .A(
        MCInst_MC3_r3Inst_XORInst_0_1_n5 ), .B(
        MCInst_MC3_r3Inst_XORInst_0_1_n4 ), .ZN(Feedback[1]) );
  XNOR2_X1 MCInst_MC3_r3Inst_XORInst_0_1_U2  ( .A(MCInst_MC3_v3_3 [1]), .B(
        MCInst_MC3_v2_3 [1]), .ZN(MCInst_MC3_r3Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst_MC3_r3Inst_XORInst_0_1_U1  ( .A(MCInst_MC3_v0_3 [1]), .B(
        MCInst_MC3_v1_3 [1]), .Z(MCInst_MC3_r3Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst_MC3_r3Inst_XORInst_0_2_U3  ( .A(
        MCInst_MC3_r3Inst_XORInst_0_2_n5 ), .B(
        MCInst_MC3_r3Inst_XORInst_0_2_n4 ), .ZN(Feedback[2]) );
  XNOR2_X1 MCInst_MC3_r3Inst_XORInst_0_2_U2  ( .A(MCInst_MC3_v3_3 [2]), .B(
        MCInst_MC3_v2_3 [2]), .ZN(MCInst_MC3_r3Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst_MC3_r3Inst_XORInst_0_2_U1  ( .A(MCInst_MC3_v0_0 [3]), .B(
        MCInst_MC3_v1_3 [2]), .Z(MCInst_MC3_r3Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst_MC3_r3Inst_XORInst_0_3_U3  ( .A(
        MCInst_MC3_r3Inst_XORInst_0_3_n5 ), .B(
        MCInst_MC3_r3Inst_XORInst_0_3_n4 ), .ZN(Feedback[3]) );
  XNOR2_X1 MCInst_MC3_r3Inst_XORInst_0_3_U2  ( .A(MCInst_MC3_v3_3 [3]), .B(
        MCInst_MC3_v2_3 [3]), .ZN(MCInst_MC3_r3Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst_MC3_r3Inst_XORInst_0_3_U1  ( .A(MCInst_MC3_v0_3 [3]), .B(
        Red_MCInst_MC3_v1_1[0] ), .Z(MCInst_MC3_r3Inst_XORInst_0_3_n5 ) );
  DFF_X1 StateReg_s_current_state_reg[0]  ( .D(Feedback[0]), .CK(clk), .Q(
        SubCellInput[0]) );
  DFF_X1 StateReg_s_current_state_reg[1]  ( .D(Feedback[1]), .CK(clk), .Q(
        SubCellInput[1]) );
  DFF_X1 StateReg_s_current_state_reg[2]  ( .D(Feedback[2]), .CK(clk), .Q(
        SubCellInput[2]) );
  DFF_X1 StateReg_s_current_state_reg[3]  ( .D(Feedback[3]), .CK(clk), .Q(
        SubCellInput[3]) );
  DFF_X1 StateReg_s_current_state_reg[4]  ( .D(Feedback[4]), .CK(clk), .Q(
        SubCellInput[4]) );
  DFF_X1 StateReg_s_current_state_reg[5]  ( .D(Feedback[5]), .CK(clk), .Q(
        SubCellInput[5]) );
  DFF_X1 StateReg_s_current_state_reg[6]  ( .D(Feedback[6]), .CK(clk), .Q(
        SubCellInput[6]) );
  DFF_X1 StateReg_s_current_state_reg[7]  ( .D(Feedback[7]), .CK(clk), .Q(
        SubCellInput[7]) );
  DFF_X1 StateReg_s_current_state_reg[8]  ( .D(Feedback[8]), .CK(clk), .Q(
        SubCellInput[8]) );
  DFF_X1 StateReg_s_current_state_reg[9]  ( .D(Feedback[9]), .CK(clk), .Q(
        SubCellInput[9]) );
  DFF_X1 StateReg_s_current_state_reg[10]  ( .D(Feedback[10]), .CK(clk), .Q(
        SubCellInput[10]) );
  DFF_X1 StateReg_s_current_state_reg[11]  ( .D(Feedback[11]), .CK(clk), .Q(
        SubCellInput[11]) );
  DFF_X1 StateReg_s_current_state_reg[12]  ( .D(Feedback[12]), .CK(clk), .Q(
        SubCellInput[12]) );
  DFF_X1 StateReg_s_current_state_reg[13]  ( .D(Feedback[13]), .CK(clk), .Q(
        SubCellInput[13]) );
  DFF_X1 StateReg_s_current_state_reg[14]  ( .D(Feedback[14]), .CK(clk), .Q(
        SubCellInput[14]) );
  DFF_X1 StateReg_s_current_state_reg[15]  ( .D(Feedback[15]), .CK(clk), .Q(
        SubCellInput[15]) );
  DFF_X1 StateReg_s_current_state_reg[16]  ( .D(Feedback[16]), .CK(clk), .Q(
        SubCellInput[16]) );
  DFF_X1 StateReg_s_current_state_reg[17]  ( .D(Feedback[17]), .CK(clk), .Q(
        SubCellInput[17]) );
  DFF_X1 StateReg_s_current_state_reg[18]  ( .D(Feedback[18]), .CK(clk), .Q(
        SubCellInput[18]) );
  DFF_X1 StateReg_s_current_state_reg[19]  ( .D(Feedback[19]), .CK(clk), .Q(
        SubCellInput[19]) );
  DFF_X1 StateReg_s_current_state_reg[20]  ( .D(Feedback[20]), .CK(clk), .Q(
        SubCellInput[20]) );
  DFF_X1 StateReg_s_current_state_reg[21]  ( .D(Feedback[21]), .CK(clk), .Q(
        SubCellInput[21]) );
  DFF_X1 StateReg_s_current_state_reg[22]  ( .D(Feedback[22]), .CK(clk), .Q(
        SubCellInput[22]) );
  DFF_X1 StateReg_s_current_state_reg[23]  ( .D(Feedback[23]), .CK(clk), .Q(
        SubCellInput[23]) );
  DFF_X1 StateReg_s_current_state_reg[24]  ( .D(Feedback[24]), .CK(clk), .Q(
        SubCellInput[24]) );
  DFF_X1 StateReg_s_current_state_reg[25]  ( .D(Feedback[25]), .CK(clk), .Q(
        SubCellInput[25]) );
  DFF_X1 StateReg_s_current_state_reg[26]  ( .D(Feedback[26]), .CK(clk), .Q(
        SubCellInput[26]) );
  DFF_X1 StateReg_s_current_state_reg[27]  ( .D(Feedback[27]), .CK(clk), .Q(
        SubCellInput[27]) );
  DFF_X1 StateReg_s_current_state_reg[28]  ( .D(Feedback[28]), .CK(clk), .Q(
        SubCellInput[28]) );
  DFF_X1 StateReg_s_current_state_reg[29]  ( .D(Feedback[29]), .CK(clk), .Q(
        SubCellInput[29]) );
  DFF_X1 StateReg_s_current_state_reg[30]  ( .D(Feedback[30]), .CK(clk), .Q(
        SubCellInput[30]) );
  DFF_X1 StateReg_s_current_state_reg[31]  ( .D(Feedback[31]), .CK(clk), .Q(
        SubCellInput[31]) );
  DFF_X1 StateReg_s_current_state_reg[32]  ( .D(Feedback[32]), .CK(clk), .Q(
        SubCellInput[32]) );
  DFF_X1 StateReg_s_current_state_reg[33]  ( .D(Feedback[33]), .CK(clk), .Q(
        SubCellInput[33]) );
  DFF_X1 StateReg_s_current_state_reg[34]  ( .D(Feedback[34]), .CK(clk), .Q(
        SubCellInput[34]) );
  DFF_X1 StateReg_s_current_state_reg[35]  ( .D(Feedback[35]), .CK(clk), .Q(
        SubCellInput[35]) );
  DFF_X1 StateReg_s_current_state_reg[36]  ( .D(Feedback[36]), .CK(clk), .Q(
        SubCellInput[36]) );
  DFF_X1 StateReg_s_current_state_reg[37]  ( .D(Feedback[37]), .CK(clk), .Q(
        SubCellInput[37]) );
  DFF_X1 StateReg_s_current_state_reg[38]  ( .D(Feedback[38]), .CK(clk), .Q(
        SubCellInput[38]) );
  DFF_X1 StateReg_s_current_state_reg[39]  ( .D(Feedback[39]), .CK(clk), .Q(
        SubCellInput[39]) );
  DFF_X1 StateReg_s_current_state_reg[40]  ( .D(Feedback[40]), .CK(clk), .Q(
        SubCellInput[40]) );
  DFF_X1 StateReg_s_current_state_reg[41]  ( .D(Feedback[41]), .CK(clk), .Q(
        SubCellInput[41]) );
  DFF_X1 StateReg_s_current_state_reg[42]  ( .D(Feedback[42]), .CK(clk), .Q(
        SubCellInput[42]) );
  DFF_X1 StateReg_s_current_state_reg[43]  ( .D(Feedback[43]), .CK(clk), .Q(
        SubCellInput[43]) );
  DFF_X1 StateReg_s_current_state_reg[44]  ( .D(Feedback[44]), .CK(clk), .Q(
        SubCellInput[44]) );
  DFF_X1 StateReg_s_current_state_reg[45]  ( .D(Feedback[45]), .CK(clk), .Q(
        SubCellInput[45]) );
  DFF_X1 StateReg_s_current_state_reg[46]  ( .D(Feedback[46]), .CK(clk), .Q(
        SubCellInput[46]) );
  DFF_X1 StateReg_s_current_state_reg[47]  ( .D(Feedback[47]), .CK(clk), .Q(
        SubCellInput[47]) );
  DFF_X1 StateReg_s_current_state_reg[48]  ( .D(Feedback[48]), .CK(clk), .Q(
        SubCellInput[48]) );
  DFF_X1 StateReg_s_current_state_reg[49]  ( .D(Feedback[49]), .CK(clk), .Q(
        SubCellInput[49]) );
  DFF_X1 StateReg_s_current_state_reg[50]  ( .D(Feedback[50]), .CK(clk), .Q(
        SubCellInput[50]) );
  DFF_X1 StateReg_s_current_state_reg[51]  ( .D(Feedback[51]), .CK(clk), .Q(
        SubCellInput[51]) );
  DFF_X1 StateReg_s_current_state_reg[52]  ( .D(Feedback[52]), .CK(clk), .Q(
        SubCellInput[52]) );
  DFF_X1 StateReg_s_current_state_reg[53]  ( .D(Feedback[53]), .CK(clk), .Q(
        SubCellInput[53]) );
  DFF_X1 StateReg_s_current_state_reg[54]  ( .D(Feedback[54]), .CK(clk), .Q(
        SubCellInput[54]) );
  DFF_X1 StateReg_s_current_state_reg[55]  ( .D(Feedback[55]), .CK(clk), .Q(
        SubCellInput[55]) );
  DFF_X1 StateReg_s_current_state_reg[56]  ( .D(Feedback[56]), .CK(clk), .Q(
        SubCellInput[56]) );
  DFF_X1 StateReg_s_current_state_reg[57]  ( .D(Feedback[57]), .CK(clk), .Q(
        SubCellInput[57]) );
  DFF_X1 StateReg_s_current_state_reg[58]  ( .D(Feedback[58]), .CK(clk), .Q(
        SubCellInput[58]) );
  DFF_X1 StateReg_s_current_state_reg[59]  ( .D(Feedback[59]), .CK(clk), .Q(
        SubCellInput[59]) );
  DFF_X1 StateReg_s_current_state_reg[60]  ( .D(Feedback[60]), .CK(clk), .Q(
        SubCellInput[60]) );
  DFF_X1 StateReg_s_current_state_reg[61]  ( .D(Feedback[61]), .CK(clk), .Q(
        SubCellInput[61]) );
  DFF_X1 StateReg_s_current_state_reg[62]  ( .D(Feedback[62]), .CK(clk), .Q(
        SubCellInput[62]) );
  DFF_X1 StateReg_s_current_state_reg[63]  ( .D(Feedback[63]), .CK(clk), .Q(
        SubCellInput[63]) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_0_U6  ( .A1(SubCellInput[2]), .A2(
        SubCellInst2_LFInst_0_LFInst_0_n4 ), .ZN(
        SubCellInst2_LFInst_0_LFInst_0_n5 ) );
  INV_X1 SubCellInst2_LFInst_0_LFInst_0_U5  ( .A(SubCellInput[1]), .ZN(
        SubCellInst2_LFInst_0_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst2_LFInst_0_LFInst_0_U4  ( .A(SubCellInput[0]), .B(
        SubCellInput[3]), .Z(SubCellInst2_LFInst_0_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst2_LFInst_0_LFInst_0_U3  ( .A(
        SubCellInst2_LFInst_0_LFInst_0_n6 ), .B(
        SubCellInst2_LFInst_0_LFInst_0_n5 ), .ZN(MCInst2_MC0_v3_2 [3]) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_1_U12  ( .A1(
        SubCellInst2_LFInst_0_LFInst_1_n18 ), .A2(
        SubCellInst2_LFInst_0_LFInst_1_n17 ), .ZN(MCInst2_MC0_v3_0 [2]) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_1_U11  ( .A1(SubCellInput[1]), .A2(
        SubCellInst2_LFInst_0_LFInst_1_n16 ), .ZN(
        SubCellInst2_LFInst_0_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst2_LFInst_0_LFInst_1_U10  ( .A1(SubCellInput[3]), .A2(
        SubCellInst2_LFInst_0_LFInst_1_n15 ), .ZN(
        SubCellInst2_LFInst_0_LFInst_1_n16 ) );
  AND2_X1 SubCellInst2_LFInst_0_LFInst_1_U9  ( .A1(SubCellInput[0]), .A2(
        SubCellInput[2]), .ZN(SubCellInst2_LFInst_0_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_1_U8  ( .A1(SubCellInput[3]), .A2(
        SubCellInst2_LFInst_0_LFInst_1_n14 ), .ZN(
        SubCellInst2_LFInst_0_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_1_U7  ( .A1(
        SubCellInst2_LFInst_0_LFInst_1_n13 ), .A2(
        SubCellInst2_LFInst_0_LFInst_1_n12 ), .ZN(
        SubCellInst2_LFInst_0_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_1_U6  ( .A1(SubCellInput[0]), .A2(
        SubCellInput[2]), .ZN(SubCellInst2_LFInst_0_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_1_U5  ( .A1(
        SubCellInst2_LFInst_0_LFInst_1_n11 ), .A2(
        SubCellInst2_LFInst_0_LFInst_1_n10 ), .ZN(
        SubCellInst2_LFInst_0_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_1_U4  ( .A1(SubCellInput[0]), .A2(
        SubCellInput[1]), .ZN(SubCellInst2_LFInst_0_LFInst_1_n10 ) );
  INV_X1 SubCellInst2_LFInst_0_LFInst_1_U3  ( .A(SubCellInput[2]), .ZN(
        SubCellInst2_LFInst_0_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_2_U11  ( .A1(
        SubCellInst2_LFInst_0_LFInst_2_n22 ), .A2(
        SubCellInst2_LFInst_0_LFInst_2_n21 ), .ZN(Red_MCInst2_MC0_v3_1[0] )
         );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_2_U10  ( .A1(SubCellInput[2]), .A2(
        SubCellInst2_LFInst_0_LFInst_2_n20 ), .ZN(
        SubCellInst2_LFInst_0_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst2_LFInst_0_LFInst_2_U9  ( .A1(SubCellInput[1]), .A2(
        SubCellInst2_LFInst_0_LFInst_2_n19 ), .ZN(
        SubCellInst2_LFInst_0_LFInst_2_n20 ) );
  INV_X1 SubCellInst2_LFInst_0_LFInst_2_U8  ( .A(SubCellInput[3]), .ZN(
        SubCellInst2_LFInst_0_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_2_U7  ( .A1(
        SubCellInst2_LFInst_0_LFInst_2_n18 ), .A2(
        SubCellInst2_LFInst_0_LFInst_2_n17 ), .ZN(
        SubCellInst2_LFInst_0_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst2_LFInst_0_LFInst_2_U6  ( .A(
        SubCellInst2_LFInst_0_LFInst_2_n16 ), .B(SubCellInput[2]), .Z(
        SubCellInst2_LFInst_0_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_2_U5  ( .A1(SubCellInput[0]), .A2(
        SubCellInput[1]), .ZN(SubCellInst2_LFInst_0_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_2_U4  ( .A1(
        SubCellInst2_LFInst_0_LFInst_2_n15 ), .A2(SubCellInput[3]), .ZN(
        SubCellInst2_LFInst_0_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst2_LFInst_0_LFInst_2_U3  ( .A(SubCellInput[0]), .B(
        SubCellInput[1]), .ZN(SubCellInst2_LFInst_0_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_3_U9  ( .A1(
        SubCellInst2_LFInst_0_LFInst_3_n16 ), .A2(
        SubCellInst2_LFInst_0_LFInst_3_n15 ), .ZN(MCInst2_MC0_v3_2 [2]) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_3_U8  ( .A1(SubCellInput[1]), .A2(
        SubCellInst2_LFInst_0_LFInst_3_n14 ), .ZN(
        SubCellInst2_LFInst_0_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst2_LFInst_0_LFInst_3_U7  ( .A(SubCellInput[3]), .B(
        SubCellInput[2]), .Z(SubCellInst2_LFInst_0_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_3_U6  ( .A1(
        SubCellInst2_LFInst_0_LFInst_3_n13 ), .A2(
        SubCellInst2_LFInst_0_LFInst_3_n12 ), .ZN(
        SubCellInst2_LFInst_0_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_0_LFInst_3_U5  ( .A1(SubCellInput[0]), .A2(
        SubCellInput[2]), .ZN(SubCellInst2_LFInst_0_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst2_LFInst_0_LFInst_3_U4  ( .A(SubCellInput[0]), .B(
        SubCellInst2_LFInst_0_LFInst_3_n11 ), .ZN(
        SubCellInst2_LFInst_0_LFInst_3_n13 ) );
  OR2_X1 SubCellInst2_LFInst_0_LFInst_3_U3  ( .A1(SubCellInput[3]), .A2(
        SubCellInput[1]), .ZN(SubCellInst2_LFInst_0_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_0_U6  ( .A1(SubCellInput[6]), .A2(
        SubCellInst2_LFInst_1_LFInst_0_n4 ), .ZN(
        SubCellInst2_LFInst_1_LFInst_0_n5 ) );
  INV_X1 SubCellInst2_LFInst_1_LFInst_0_U5  ( .A(SubCellInput[5]), .ZN(
        SubCellInst2_LFInst_1_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst2_LFInst_1_LFInst_0_U4  ( .A(SubCellInput[4]), .B(
        SubCellInput[7]), .Z(SubCellInst2_LFInst_1_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst2_LFInst_1_LFInst_0_U3  ( .A(
        SubCellInst2_LFInst_1_LFInst_0_n6 ), .B(
        SubCellInst2_LFInst_1_LFInst_0_n5 ), .ZN(MCInst2_MC3_v3_2 [3]) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_1_U12  ( .A1(
        SubCellInst2_LFInst_1_LFInst_1_n18 ), .A2(
        SubCellInst2_LFInst_1_LFInst_1_n17 ), .ZN(MCInst2_MC3_v3_0 [2]) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_1_U11  ( .A1(SubCellInput[5]), .A2(
        SubCellInst2_LFInst_1_LFInst_1_n16 ), .ZN(
        SubCellInst2_LFInst_1_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst2_LFInst_1_LFInst_1_U10  ( .A1(SubCellInput[7]), .A2(
        SubCellInst2_LFInst_1_LFInst_1_n15 ), .ZN(
        SubCellInst2_LFInst_1_LFInst_1_n16 ) );
  AND2_X1 SubCellInst2_LFInst_1_LFInst_1_U9  ( .A1(SubCellInput[4]), .A2(
        SubCellInput[6]), .ZN(SubCellInst2_LFInst_1_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_1_U8  ( .A1(SubCellInput[7]), .A2(
        SubCellInst2_LFInst_1_LFInst_1_n14 ), .ZN(
        SubCellInst2_LFInst_1_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_1_U7  ( .A1(
        SubCellInst2_LFInst_1_LFInst_1_n13 ), .A2(
        SubCellInst2_LFInst_1_LFInst_1_n12 ), .ZN(
        SubCellInst2_LFInst_1_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_1_U6  ( .A1(SubCellInput[4]), .A2(
        SubCellInput[6]), .ZN(SubCellInst2_LFInst_1_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_1_U5  ( .A1(
        SubCellInst2_LFInst_1_LFInst_1_n11 ), .A2(
        SubCellInst2_LFInst_1_LFInst_1_n10 ), .ZN(
        SubCellInst2_LFInst_1_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_1_U4  ( .A1(SubCellInput[4]), .A2(
        SubCellInput[5]), .ZN(SubCellInst2_LFInst_1_LFInst_1_n10 ) );
  INV_X1 SubCellInst2_LFInst_1_LFInst_1_U3  ( .A(SubCellInput[6]), .ZN(
        SubCellInst2_LFInst_1_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_2_U11  ( .A1(
        SubCellInst2_LFInst_1_LFInst_2_n22 ), .A2(
        SubCellInst2_LFInst_1_LFInst_2_n21 ), .ZN(Red_MCInst2_MC3_v3_1[0] )
         );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_2_U10  ( .A1(SubCellInput[6]), .A2(
        SubCellInst2_LFInst_1_LFInst_2_n20 ), .ZN(
        SubCellInst2_LFInst_1_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst2_LFInst_1_LFInst_2_U9  ( .A1(SubCellInput[5]), .A2(
        SubCellInst2_LFInst_1_LFInst_2_n19 ), .ZN(
        SubCellInst2_LFInst_1_LFInst_2_n20 ) );
  INV_X1 SubCellInst2_LFInst_1_LFInst_2_U8  ( .A(SubCellInput[7]), .ZN(
        SubCellInst2_LFInst_1_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_2_U7  ( .A1(
        SubCellInst2_LFInst_1_LFInst_2_n18 ), .A2(
        SubCellInst2_LFInst_1_LFInst_2_n17 ), .ZN(
        SubCellInst2_LFInst_1_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst2_LFInst_1_LFInst_2_U6  ( .A(
        SubCellInst2_LFInst_1_LFInst_2_n16 ), .B(SubCellInput[6]), .Z(
        SubCellInst2_LFInst_1_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_2_U5  ( .A1(SubCellInput[4]), .A2(
        SubCellInput[5]), .ZN(SubCellInst2_LFInst_1_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_2_U4  ( .A1(
        SubCellInst2_LFInst_1_LFInst_2_n15 ), .A2(SubCellInput[7]), .ZN(
        SubCellInst2_LFInst_1_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst2_LFInst_1_LFInst_2_U3  ( .A(SubCellInput[4]), .B(
        SubCellInput[5]), .ZN(SubCellInst2_LFInst_1_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_3_U9  ( .A1(
        SubCellInst2_LFInst_1_LFInst_3_n16 ), .A2(
        SubCellInst2_LFInst_1_LFInst_3_n15 ), .ZN(MCInst2_MC3_v3_2 [2]) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_3_U8  ( .A1(SubCellInput[5]), .A2(
        SubCellInst2_LFInst_1_LFInst_3_n14 ), .ZN(
        SubCellInst2_LFInst_1_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst2_LFInst_1_LFInst_3_U7  ( .A(SubCellInput[7]), .B(
        SubCellInput[6]), .Z(SubCellInst2_LFInst_1_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_3_U6  ( .A1(
        SubCellInst2_LFInst_1_LFInst_3_n13 ), .A2(
        SubCellInst2_LFInst_1_LFInst_3_n12 ), .ZN(
        SubCellInst2_LFInst_1_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_1_LFInst_3_U5  ( .A1(SubCellInput[4]), .A2(
        SubCellInput[6]), .ZN(SubCellInst2_LFInst_1_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst2_LFInst_1_LFInst_3_U4  ( .A(SubCellInput[4]), .B(
        SubCellInst2_LFInst_1_LFInst_3_n11 ), .ZN(
        SubCellInst2_LFInst_1_LFInst_3_n13 ) );
  OR2_X1 SubCellInst2_LFInst_1_LFInst_3_U3  ( .A1(SubCellInput[7]), .A2(
        SubCellInput[5]), .ZN(SubCellInst2_LFInst_1_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_0_U6  ( .A1(SubCellInput[10]), .A2(
        SubCellInst2_LFInst_2_LFInst_0_n4 ), .ZN(
        SubCellInst2_LFInst_2_LFInst_0_n5 ) );
  INV_X1 SubCellInst2_LFInst_2_LFInst_0_U5  ( .A(SubCellInput[9]), .ZN(
        SubCellInst2_LFInst_2_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst2_LFInst_2_LFInst_0_U4  ( .A(SubCellInput[8]), .B(
        SubCellInput[11]), .Z(SubCellInst2_LFInst_2_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst2_LFInst_2_LFInst_0_U3  ( .A(
        SubCellInst2_LFInst_2_LFInst_0_n6 ), .B(
        SubCellInst2_LFInst_2_LFInst_0_n5 ), .ZN(MCInst2_MC2_v3_2 [3]) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_1_U12  ( .A1(
        SubCellInst2_LFInst_2_LFInst_1_n18 ), .A2(
        SubCellInst2_LFInst_2_LFInst_1_n17 ), .ZN(MCInst2_MC2_v3_0 [2]) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_1_U11  ( .A1(SubCellInput[9]), .A2(
        SubCellInst2_LFInst_2_LFInst_1_n16 ), .ZN(
        SubCellInst2_LFInst_2_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst2_LFInst_2_LFInst_1_U10  ( .A1(SubCellInput[11]), .A2(
        SubCellInst2_LFInst_2_LFInst_1_n15 ), .ZN(
        SubCellInst2_LFInst_2_LFInst_1_n16 ) );
  AND2_X1 SubCellInst2_LFInst_2_LFInst_1_U9  ( .A1(SubCellInput[8]), .A2(
        SubCellInput[10]), .ZN(SubCellInst2_LFInst_2_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_1_U8  ( .A1(SubCellInput[11]), .A2(
        SubCellInst2_LFInst_2_LFInst_1_n14 ), .ZN(
        SubCellInst2_LFInst_2_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_1_U7  ( .A1(
        SubCellInst2_LFInst_2_LFInst_1_n13 ), .A2(
        SubCellInst2_LFInst_2_LFInst_1_n12 ), .ZN(
        SubCellInst2_LFInst_2_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_1_U6  ( .A1(SubCellInput[8]), .A2(
        SubCellInput[10]), .ZN(SubCellInst2_LFInst_2_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_1_U5  ( .A1(
        SubCellInst2_LFInst_2_LFInst_1_n11 ), .A2(
        SubCellInst2_LFInst_2_LFInst_1_n10 ), .ZN(
        SubCellInst2_LFInst_2_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_1_U4  ( .A1(SubCellInput[8]), .A2(
        SubCellInput[9]), .ZN(SubCellInst2_LFInst_2_LFInst_1_n10 ) );
  INV_X1 SubCellInst2_LFInst_2_LFInst_1_U3  ( .A(SubCellInput[10]), .ZN(
        SubCellInst2_LFInst_2_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_2_U11  ( .A1(
        SubCellInst2_LFInst_2_LFInst_2_n22 ), .A2(
        SubCellInst2_LFInst_2_LFInst_2_n21 ), .ZN(Red_MCInst2_MC2_v3_1[0] )
         );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_2_U10  ( .A1(SubCellInput[10]), .A2(
        SubCellInst2_LFInst_2_LFInst_2_n20 ), .ZN(
        SubCellInst2_LFInst_2_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst2_LFInst_2_LFInst_2_U9  ( .A1(SubCellInput[9]), .A2(
        SubCellInst2_LFInst_2_LFInst_2_n19 ), .ZN(
        SubCellInst2_LFInst_2_LFInst_2_n20 ) );
  INV_X1 SubCellInst2_LFInst_2_LFInst_2_U8  ( .A(SubCellInput[11]), .ZN(
        SubCellInst2_LFInst_2_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_2_U7  ( .A1(
        SubCellInst2_LFInst_2_LFInst_2_n18 ), .A2(
        SubCellInst2_LFInst_2_LFInst_2_n17 ), .ZN(
        SubCellInst2_LFInst_2_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst2_LFInst_2_LFInst_2_U6  ( .A(
        SubCellInst2_LFInst_2_LFInst_2_n16 ), .B(SubCellInput[10]), .Z(
        SubCellInst2_LFInst_2_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_2_U5  ( .A1(SubCellInput[8]), .A2(
        SubCellInput[9]), .ZN(SubCellInst2_LFInst_2_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_2_U4  ( .A1(
        SubCellInst2_LFInst_2_LFInst_2_n15 ), .A2(SubCellInput[11]), .ZN(
        SubCellInst2_LFInst_2_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst2_LFInst_2_LFInst_2_U3  ( .A(SubCellInput[8]), .B(
        SubCellInput[9]), .ZN(SubCellInst2_LFInst_2_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_3_U9  ( .A1(
        SubCellInst2_LFInst_2_LFInst_3_n16 ), .A2(
        SubCellInst2_LFInst_2_LFInst_3_n15 ), .ZN(MCInst2_MC2_v3_2 [2]) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_3_U8  ( .A1(SubCellInput[9]), .A2(
        SubCellInst2_LFInst_2_LFInst_3_n14 ), .ZN(
        SubCellInst2_LFInst_2_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst2_LFInst_2_LFInst_3_U7  ( .A(SubCellInput[11]), .B(
        SubCellInput[10]), .Z(SubCellInst2_LFInst_2_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_3_U6  ( .A1(
        SubCellInst2_LFInst_2_LFInst_3_n13 ), .A2(
        SubCellInst2_LFInst_2_LFInst_3_n12 ), .ZN(
        SubCellInst2_LFInst_2_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_2_LFInst_3_U5  ( .A1(SubCellInput[8]), .A2(
        SubCellInput[10]), .ZN(SubCellInst2_LFInst_2_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst2_LFInst_2_LFInst_3_U4  ( .A(SubCellInput[8]), .B(
        SubCellInst2_LFInst_2_LFInst_3_n11 ), .ZN(
        SubCellInst2_LFInst_2_LFInst_3_n13 ) );
  OR2_X1 SubCellInst2_LFInst_2_LFInst_3_U3  ( .A1(SubCellInput[11]), .A2(
        SubCellInput[9]), .ZN(SubCellInst2_LFInst_2_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_0_U6  ( .A1(SubCellInput[14]), .A2(
        SubCellInst2_LFInst_3_LFInst_0_n4 ), .ZN(
        SubCellInst2_LFInst_3_LFInst_0_n5 ) );
  INV_X1 SubCellInst2_LFInst_3_LFInst_0_U5  ( .A(SubCellInput[13]), .ZN(
        SubCellInst2_LFInst_3_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst2_LFInst_3_LFInst_0_U4  ( .A(SubCellInput[12]), .B(
        SubCellInput[15]), .Z(SubCellInst2_LFInst_3_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst2_LFInst_3_LFInst_0_U3  ( .A(
        SubCellInst2_LFInst_3_LFInst_0_n6 ), .B(
        SubCellInst2_LFInst_3_LFInst_0_n5 ), .ZN(MCInst2_MC1_v3_2 [3]) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_1_U12  ( .A1(
        SubCellInst2_LFInst_3_LFInst_1_n18 ), .A2(
        SubCellInst2_LFInst_3_LFInst_1_n17 ), .ZN(MCInst2_MC1_v3_0 [2]) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_1_U11  ( .A1(SubCellInput[13]), .A2(
        SubCellInst2_LFInst_3_LFInst_1_n16 ), .ZN(
        SubCellInst2_LFInst_3_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst2_LFInst_3_LFInst_1_U10  ( .A1(SubCellInput[15]), .A2(
        SubCellInst2_LFInst_3_LFInst_1_n15 ), .ZN(
        SubCellInst2_LFInst_3_LFInst_1_n16 ) );
  AND2_X1 SubCellInst2_LFInst_3_LFInst_1_U9  ( .A1(SubCellInput[12]), .A2(
        SubCellInput[14]), .ZN(SubCellInst2_LFInst_3_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_1_U8  ( .A1(SubCellInput[15]), .A2(
        SubCellInst2_LFInst_3_LFInst_1_n14 ), .ZN(
        SubCellInst2_LFInst_3_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_1_U7  ( .A1(
        SubCellInst2_LFInst_3_LFInst_1_n13 ), .A2(
        SubCellInst2_LFInst_3_LFInst_1_n12 ), .ZN(
        SubCellInst2_LFInst_3_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_1_U6  ( .A1(SubCellInput[12]), .A2(
        SubCellInput[14]), .ZN(SubCellInst2_LFInst_3_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_1_U5  ( .A1(
        SubCellInst2_LFInst_3_LFInst_1_n11 ), .A2(
        SubCellInst2_LFInst_3_LFInst_1_n10 ), .ZN(
        SubCellInst2_LFInst_3_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_1_U4  ( .A1(SubCellInput[12]), .A2(
        SubCellInput[13]), .ZN(SubCellInst2_LFInst_3_LFInst_1_n10 ) );
  INV_X1 SubCellInst2_LFInst_3_LFInst_1_U3  ( .A(SubCellInput[14]), .ZN(
        SubCellInst2_LFInst_3_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_2_U11  ( .A1(
        SubCellInst2_LFInst_3_LFInst_2_n22 ), .A2(
        SubCellInst2_LFInst_3_LFInst_2_n21 ), .ZN(Red_MCInst2_MC1_v3_1[0] )
         );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_2_U10  ( .A1(SubCellInput[14]), .A2(
        SubCellInst2_LFInst_3_LFInst_2_n20 ), .ZN(
        SubCellInst2_LFInst_3_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst2_LFInst_3_LFInst_2_U9  ( .A1(SubCellInput[13]), .A2(
        SubCellInst2_LFInst_3_LFInst_2_n19 ), .ZN(
        SubCellInst2_LFInst_3_LFInst_2_n20 ) );
  INV_X1 SubCellInst2_LFInst_3_LFInst_2_U8  ( .A(SubCellInput[15]), .ZN(
        SubCellInst2_LFInst_3_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_2_U7  ( .A1(
        SubCellInst2_LFInst_3_LFInst_2_n18 ), .A2(
        SubCellInst2_LFInst_3_LFInst_2_n17 ), .ZN(
        SubCellInst2_LFInst_3_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst2_LFInst_3_LFInst_2_U6  ( .A(
        SubCellInst2_LFInst_3_LFInst_2_n16 ), .B(SubCellInput[14]), .Z(
        SubCellInst2_LFInst_3_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_2_U5  ( .A1(SubCellInput[12]), .A2(
        SubCellInput[13]), .ZN(SubCellInst2_LFInst_3_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_2_U4  ( .A1(
        SubCellInst2_LFInst_3_LFInst_2_n15 ), .A2(SubCellInput[15]), .ZN(
        SubCellInst2_LFInst_3_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst2_LFInst_3_LFInst_2_U3  ( .A(SubCellInput[12]), .B(
        SubCellInput[13]), .ZN(SubCellInst2_LFInst_3_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_3_U9  ( .A1(
        SubCellInst2_LFInst_3_LFInst_3_n16 ), .A2(
        SubCellInst2_LFInst_3_LFInst_3_n15 ), .ZN(MCInst2_MC1_v3_2 [2]) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_3_U8  ( .A1(SubCellInput[13]), .A2(
        SubCellInst2_LFInst_3_LFInst_3_n14 ), .ZN(
        SubCellInst2_LFInst_3_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst2_LFInst_3_LFInst_3_U7  ( .A(SubCellInput[15]), .B(
        SubCellInput[14]), .Z(SubCellInst2_LFInst_3_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_3_U6  ( .A1(
        SubCellInst2_LFInst_3_LFInst_3_n13 ), .A2(
        SubCellInst2_LFInst_3_LFInst_3_n12 ), .ZN(
        SubCellInst2_LFInst_3_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_3_LFInst_3_U5  ( .A1(SubCellInput[12]), .A2(
        SubCellInput[14]), .ZN(SubCellInst2_LFInst_3_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst2_LFInst_3_LFInst_3_U4  ( .A(SubCellInput[12]), .B(
        SubCellInst2_LFInst_3_LFInst_3_n11 ), .ZN(
        SubCellInst2_LFInst_3_LFInst_3_n13 ) );
  OR2_X1 SubCellInst2_LFInst_3_LFInst_3_U3  ( .A1(SubCellInput[15]), .A2(
        SubCellInput[13]), .ZN(SubCellInst2_LFInst_3_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_0_U6  ( .A1(SubCellInput[18]), .A2(
        SubCellInst2_LFInst_4_LFInst_0_n4 ), .ZN(
        SubCellInst2_LFInst_4_LFInst_0_n5 ) );
  INV_X1 SubCellInst2_LFInst_4_LFInst_0_U5  ( .A(SubCellInput[17]), .ZN(
        SubCellInst2_LFInst_4_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst2_LFInst_4_LFInst_0_U4  ( .A(SubCellInput[16]), .B(
        SubCellInput[19]), .Z(SubCellInst2_LFInst_4_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst2_LFInst_4_LFInst_0_U3  ( .A(
        SubCellInst2_LFInst_4_LFInst_0_n6 ), .B(
        SubCellInst2_LFInst_4_LFInst_0_n5 ), .ZN(MCInst2_MC1_v2_3 [1]) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_1_U12  ( .A1(
        SubCellInst2_LFInst_4_LFInst_1_n18 ), .A2(
        SubCellInst2_LFInst_4_LFInst_1_n17 ), .ZN(MCInst2_MC1_v2_0 [2]) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_1_U11  ( .A1(SubCellInput[17]), .A2(
        SubCellInst2_LFInst_4_LFInst_1_n16 ), .ZN(
        SubCellInst2_LFInst_4_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst2_LFInst_4_LFInst_1_U10  ( .A1(SubCellInput[19]), .A2(
        SubCellInst2_LFInst_4_LFInst_1_n15 ), .ZN(
        SubCellInst2_LFInst_4_LFInst_1_n16 ) );
  AND2_X1 SubCellInst2_LFInst_4_LFInst_1_U9  ( .A1(SubCellInput[16]), .A2(
        SubCellInput[18]), .ZN(SubCellInst2_LFInst_4_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_1_U8  ( .A1(SubCellInput[19]), .A2(
        SubCellInst2_LFInst_4_LFInst_1_n14 ), .ZN(
        SubCellInst2_LFInst_4_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_1_U7  ( .A1(
        SubCellInst2_LFInst_4_LFInst_1_n13 ), .A2(
        SubCellInst2_LFInst_4_LFInst_1_n12 ), .ZN(
        SubCellInst2_LFInst_4_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_1_U6  ( .A1(SubCellInput[16]), .A2(
        SubCellInput[18]), .ZN(SubCellInst2_LFInst_4_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_1_U5  ( .A1(
        SubCellInst2_LFInst_4_LFInst_1_n11 ), .A2(
        SubCellInst2_LFInst_4_LFInst_1_n10 ), .ZN(
        SubCellInst2_LFInst_4_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_1_U4  ( .A1(SubCellInput[16]), .A2(
        SubCellInput[17]), .ZN(SubCellInst2_LFInst_4_LFInst_1_n10 ) );
  INV_X1 SubCellInst2_LFInst_4_LFInst_1_U3  ( .A(SubCellInput[18]), .ZN(
        SubCellInst2_LFInst_4_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_2_U11  ( .A1(
        SubCellInst2_LFInst_4_LFInst_2_n22 ), .A2(
        SubCellInst2_LFInst_4_LFInst_2_n21 ), .ZN(MCInst2_MC1_v2_0 [3]) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_2_U10  ( .A1(SubCellInput[18]), .A2(
        SubCellInst2_LFInst_4_LFInst_2_n20 ), .ZN(
        SubCellInst2_LFInst_4_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst2_LFInst_4_LFInst_2_U9  ( .A1(SubCellInput[17]), .A2(
        SubCellInst2_LFInst_4_LFInst_2_n19 ), .ZN(
        SubCellInst2_LFInst_4_LFInst_2_n20 ) );
  INV_X1 SubCellInst2_LFInst_4_LFInst_2_U8  ( .A(SubCellInput[19]), .ZN(
        SubCellInst2_LFInst_4_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_2_U7  ( .A1(
        SubCellInst2_LFInst_4_LFInst_2_n18 ), .A2(
        SubCellInst2_LFInst_4_LFInst_2_n17 ), .ZN(
        SubCellInst2_LFInst_4_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst2_LFInst_4_LFInst_2_U6  ( .A(
        SubCellInst2_LFInst_4_LFInst_2_n16 ), .B(SubCellInput[18]), .Z(
        SubCellInst2_LFInst_4_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_2_U5  ( .A1(SubCellInput[16]), .A2(
        SubCellInput[17]), .ZN(SubCellInst2_LFInst_4_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_2_U4  ( .A1(
        SubCellInst2_LFInst_4_LFInst_2_n15 ), .A2(SubCellInput[19]), .ZN(
        SubCellInst2_LFInst_4_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst2_LFInst_4_LFInst_2_U3  ( .A(SubCellInput[16]), .B(
        SubCellInput[17]), .ZN(SubCellInst2_LFInst_4_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_3_U9  ( .A1(
        SubCellInst2_LFInst_4_LFInst_3_n16 ), .A2(
        SubCellInst2_LFInst_4_LFInst_3_n15 ), .ZN(MCInst2_MC1_v2_0 [0]) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_3_U8  ( .A1(SubCellInput[17]), .A2(
        SubCellInst2_LFInst_4_LFInst_3_n14 ), .ZN(
        SubCellInst2_LFInst_4_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst2_LFInst_4_LFInst_3_U7  ( .A(SubCellInput[19]), .B(
        SubCellInput[18]), .Z(SubCellInst2_LFInst_4_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_3_U6  ( .A1(
        SubCellInst2_LFInst_4_LFInst_3_n13 ), .A2(
        SubCellInst2_LFInst_4_LFInst_3_n12 ), .ZN(
        SubCellInst2_LFInst_4_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_4_LFInst_3_U5  ( .A1(SubCellInput[16]), .A2(
        SubCellInput[18]), .ZN(SubCellInst2_LFInst_4_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst2_LFInst_4_LFInst_3_U4  ( .A(SubCellInput[16]), .B(
        SubCellInst2_LFInst_4_LFInst_3_n11 ), .ZN(
        SubCellInst2_LFInst_4_LFInst_3_n13 ) );
  OR2_X1 SubCellInst2_LFInst_4_LFInst_3_U3  ( .A1(SubCellInput[19]), .A2(
        SubCellInput[17]), .ZN(SubCellInst2_LFInst_4_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_0_U6  ( .A1(SubCellInput[22]), .A2(
        SubCellInst2_LFInst_5_LFInst_0_n4 ), .ZN(
        SubCellInst2_LFInst_5_LFInst_0_n5 ) );
  INV_X1 SubCellInst2_LFInst_5_LFInst_0_U5  ( .A(SubCellInput[21]), .ZN(
        SubCellInst2_LFInst_5_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst2_LFInst_5_LFInst_0_U4  ( .A(SubCellInput[20]), .B(
        SubCellInput[23]), .Z(SubCellInst2_LFInst_5_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst2_LFInst_5_LFInst_0_U3  ( .A(
        SubCellInst2_LFInst_5_LFInst_0_n6 ), .B(
        SubCellInst2_LFInst_5_LFInst_0_n5 ), .ZN(MCInst2_MC0_v2_3 [1]) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_1_U12  ( .A1(
        SubCellInst2_LFInst_5_LFInst_1_n18 ), .A2(
        SubCellInst2_LFInst_5_LFInst_1_n17 ), .ZN(MCInst2_MC0_v2_0 [2]) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_1_U11  ( .A1(SubCellInput[21]), .A2(
        SubCellInst2_LFInst_5_LFInst_1_n16 ), .ZN(
        SubCellInst2_LFInst_5_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst2_LFInst_5_LFInst_1_U10  ( .A1(SubCellInput[23]), .A2(
        SubCellInst2_LFInst_5_LFInst_1_n15 ), .ZN(
        SubCellInst2_LFInst_5_LFInst_1_n16 ) );
  AND2_X1 SubCellInst2_LFInst_5_LFInst_1_U9  ( .A1(SubCellInput[20]), .A2(
        SubCellInput[22]), .ZN(SubCellInst2_LFInst_5_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_1_U8  ( .A1(SubCellInput[23]), .A2(
        SubCellInst2_LFInst_5_LFInst_1_n14 ), .ZN(
        SubCellInst2_LFInst_5_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_1_U7  ( .A1(
        SubCellInst2_LFInst_5_LFInst_1_n13 ), .A2(
        SubCellInst2_LFInst_5_LFInst_1_n12 ), .ZN(
        SubCellInst2_LFInst_5_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_1_U6  ( .A1(SubCellInput[20]), .A2(
        SubCellInput[22]), .ZN(SubCellInst2_LFInst_5_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_1_U5  ( .A1(
        SubCellInst2_LFInst_5_LFInst_1_n11 ), .A2(
        SubCellInst2_LFInst_5_LFInst_1_n10 ), .ZN(
        SubCellInst2_LFInst_5_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_1_U4  ( .A1(SubCellInput[20]), .A2(
        SubCellInput[21]), .ZN(SubCellInst2_LFInst_5_LFInst_1_n10 ) );
  INV_X1 SubCellInst2_LFInst_5_LFInst_1_U3  ( .A(SubCellInput[22]), .ZN(
        SubCellInst2_LFInst_5_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_2_U11  ( .A1(
        SubCellInst2_LFInst_5_LFInst_2_n22 ), .A2(
        SubCellInst2_LFInst_5_LFInst_2_n21 ), .ZN(MCInst2_MC0_v2_0 [3]) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_2_U10  ( .A1(SubCellInput[22]), .A2(
        SubCellInst2_LFInst_5_LFInst_2_n20 ), .ZN(
        SubCellInst2_LFInst_5_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst2_LFInst_5_LFInst_2_U9  ( .A1(SubCellInput[21]), .A2(
        SubCellInst2_LFInst_5_LFInst_2_n19 ), .ZN(
        SubCellInst2_LFInst_5_LFInst_2_n20 ) );
  INV_X1 SubCellInst2_LFInst_5_LFInst_2_U8  ( .A(SubCellInput[23]), .ZN(
        SubCellInst2_LFInst_5_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_2_U7  ( .A1(
        SubCellInst2_LFInst_5_LFInst_2_n18 ), .A2(
        SubCellInst2_LFInst_5_LFInst_2_n17 ), .ZN(
        SubCellInst2_LFInst_5_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst2_LFInst_5_LFInst_2_U6  ( .A(
        SubCellInst2_LFInst_5_LFInst_2_n16 ), .B(SubCellInput[22]), .Z(
        SubCellInst2_LFInst_5_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_2_U5  ( .A1(SubCellInput[20]), .A2(
        SubCellInput[21]), .ZN(SubCellInst2_LFInst_5_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_2_U4  ( .A1(
        SubCellInst2_LFInst_5_LFInst_2_n15 ), .A2(SubCellInput[23]), .ZN(
        SubCellInst2_LFInst_5_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst2_LFInst_5_LFInst_2_U3  ( .A(SubCellInput[20]), .B(
        SubCellInput[21]), .ZN(SubCellInst2_LFInst_5_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_3_U9  ( .A1(
        SubCellInst2_LFInst_5_LFInst_3_n16 ), .A2(
        SubCellInst2_LFInst_5_LFInst_3_n15 ), .ZN(MCInst2_MC0_v2_0 [0]) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_3_U8  ( .A1(SubCellInput[21]), .A2(
        SubCellInst2_LFInst_5_LFInst_3_n14 ), .ZN(
        SubCellInst2_LFInst_5_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst2_LFInst_5_LFInst_3_U7  ( .A(SubCellInput[23]), .B(
        SubCellInput[22]), .Z(SubCellInst2_LFInst_5_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_3_U6  ( .A1(
        SubCellInst2_LFInst_5_LFInst_3_n13 ), .A2(
        SubCellInst2_LFInst_5_LFInst_3_n12 ), .ZN(
        SubCellInst2_LFInst_5_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_5_LFInst_3_U5  ( .A1(SubCellInput[20]), .A2(
        SubCellInput[22]), .ZN(SubCellInst2_LFInst_5_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst2_LFInst_5_LFInst_3_U4  ( .A(SubCellInput[20]), .B(
        SubCellInst2_LFInst_5_LFInst_3_n11 ), .ZN(
        SubCellInst2_LFInst_5_LFInst_3_n13 ) );
  OR2_X1 SubCellInst2_LFInst_5_LFInst_3_U3  ( .A1(SubCellInput[23]), .A2(
        SubCellInput[21]), .ZN(SubCellInst2_LFInst_5_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_0_U6  ( .A1(SubCellInput[26]), .A2(
        SubCellInst2_LFInst_6_LFInst_0_n4 ), .ZN(
        SubCellInst2_LFInst_6_LFInst_0_n5 ) );
  INV_X1 SubCellInst2_LFInst_6_LFInst_0_U5  ( .A(SubCellInput[25]), .ZN(
        SubCellInst2_LFInst_6_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst2_LFInst_6_LFInst_0_U4  ( .A(SubCellInput[24]), .B(
        SubCellInput[27]), .Z(SubCellInst2_LFInst_6_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst2_LFInst_6_LFInst_0_U3  ( .A(
        SubCellInst2_LFInst_6_LFInst_0_n6 ), .B(
        SubCellInst2_LFInst_6_LFInst_0_n5 ), .ZN(MCInst2_MC3_v2_3 [1]) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_1_U12  ( .A1(
        SubCellInst2_LFInst_6_LFInst_1_n18 ), .A2(
        SubCellInst2_LFInst_6_LFInst_1_n17 ), .ZN(MCInst2_MC3_v2_0 [2]) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_1_U11  ( .A1(SubCellInput[25]), .A2(
        SubCellInst2_LFInst_6_LFInst_1_n16 ), .ZN(
        SubCellInst2_LFInst_6_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst2_LFInst_6_LFInst_1_U10  ( .A1(SubCellInput[27]), .A2(
        SubCellInst2_LFInst_6_LFInst_1_n15 ), .ZN(
        SubCellInst2_LFInst_6_LFInst_1_n16 ) );
  AND2_X1 SubCellInst2_LFInst_6_LFInst_1_U9  ( .A1(SubCellInput[24]), .A2(
        SubCellInput[26]), .ZN(SubCellInst2_LFInst_6_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_1_U8  ( .A1(SubCellInput[27]), .A2(
        SubCellInst2_LFInst_6_LFInst_1_n14 ), .ZN(
        SubCellInst2_LFInst_6_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_1_U7  ( .A1(
        SubCellInst2_LFInst_6_LFInst_1_n13 ), .A2(
        SubCellInst2_LFInst_6_LFInst_1_n12 ), .ZN(
        SubCellInst2_LFInst_6_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_1_U6  ( .A1(SubCellInput[24]), .A2(
        SubCellInput[26]), .ZN(SubCellInst2_LFInst_6_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_1_U5  ( .A1(
        SubCellInst2_LFInst_6_LFInst_1_n11 ), .A2(
        SubCellInst2_LFInst_6_LFInst_1_n10 ), .ZN(
        SubCellInst2_LFInst_6_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_1_U4  ( .A1(SubCellInput[24]), .A2(
        SubCellInput[25]), .ZN(SubCellInst2_LFInst_6_LFInst_1_n10 ) );
  INV_X1 SubCellInst2_LFInst_6_LFInst_1_U3  ( .A(SubCellInput[26]), .ZN(
        SubCellInst2_LFInst_6_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_2_U11  ( .A1(
        SubCellInst2_LFInst_6_LFInst_2_n22 ), .A2(
        SubCellInst2_LFInst_6_LFInst_2_n21 ), .ZN(MCInst2_MC3_v2_0 [3]) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_2_U10  ( .A1(SubCellInput[26]), .A2(
        SubCellInst2_LFInst_6_LFInst_2_n20 ), .ZN(
        SubCellInst2_LFInst_6_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst2_LFInst_6_LFInst_2_U9  ( .A1(SubCellInput[25]), .A2(
        SubCellInst2_LFInst_6_LFInst_2_n19 ), .ZN(
        SubCellInst2_LFInst_6_LFInst_2_n20 ) );
  INV_X1 SubCellInst2_LFInst_6_LFInst_2_U8  ( .A(SubCellInput[27]), .ZN(
        SubCellInst2_LFInst_6_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_2_U7  ( .A1(
        SubCellInst2_LFInst_6_LFInst_2_n18 ), .A2(
        SubCellInst2_LFInst_6_LFInst_2_n17 ), .ZN(
        SubCellInst2_LFInst_6_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst2_LFInst_6_LFInst_2_U6  ( .A(
        SubCellInst2_LFInst_6_LFInst_2_n16 ), .B(SubCellInput[26]), .Z(
        SubCellInst2_LFInst_6_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_2_U5  ( .A1(SubCellInput[24]), .A2(
        SubCellInput[25]), .ZN(SubCellInst2_LFInst_6_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_2_U4  ( .A1(
        SubCellInst2_LFInst_6_LFInst_2_n15 ), .A2(SubCellInput[27]), .ZN(
        SubCellInst2_LFInst_6_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst2_LFInst_6_LFInst_2_U3  ( .A(SubCellInput[24]), .B(
        SubCellInput[25]), .ZN(SubCellInst2_LFInst_6_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_3_U9  ( .A1(
        SubCellInst2_LFInst_6_LFInst_3_n16 ), .A2(
        SubCellInst2_LFInst_6_LFInst_3_n15 ), .ZN(MCInst2_MC3_v2_0 [0]) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_3_U8  ( .A1(SubCellInput[25]), .A2(
        SubCellInst2_LFInst_6_LFInst_3_n14 ), .ZN(
        SubCellInst2_LFInst_6_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst2_LFInst_6_LFInst_3_U7  ( .A(SubCellInput[27]), .B(
        SubCellInput[26]), .Z(SubCellInst2_LFInst_6_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_3_U6  ( .A1(
        SubCellInst2_LFInst_6_LFInst_3_n13 ), .A2(
        SubCellInst2_LFInst_6_LFInst_3_n12 ), .ZN(
        SubCellInst2_LFInst_6_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_6_LFInst_3_U5  ( .A1(SubCellInput[24]), .A2(
        SubCellInput[26]), .ZN(SubCellInst2_LFInst_6_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst2_LFInst_6_LFInst_3_U4  ( .A(SubCellInput[24]), .B(
        SubCellInst2_LFInst_6_LFInst_3_n11 ), .ZN(
        SubCellInst2_LFInst_6_LFInst_3_n13 ) );
  OR2_X1 SubCellInst2_LFInst_6_LFInst_3_U3  ( .A1(SubCellInput[27]), .A2(
        SubCellInput[25]), .ZN(SubCellInst2_LFInst_6_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_0_U6  ( .A1(SubCellInput[30]), .A2(
        SubCellInst2_LFInst_7_LFInst_0_n4 ), .ZN(
        SubCellInst2_LFInst_7_LFInst_0_n5 ) );
  INV_X1 SubCellInst2_LFInst_7_LFInst_0_U5  ( .A(SubCellInput[29]), .ZN(
        SubCellInst2_LFInst_7_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst2_LFInst_7_LFInst_0_U4  ( .A(SubCellInput[28]), .B(
        SubCellInput[31]), .Z(SubCellInst2_LFInst_7_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst2_LFInst_7_LFInst_0_U3  ( .A(
        SubCellInst2_LFInst_7_LFInst_0_n6 ), .B(
        SubCellInst2_LFInst_7_LFInst_0_n5 ), .ZN(MCInst2_MC2_v2_3 [1]) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_1_U12  ( .A1(
        SubCellInst2_LFInst_7_LFInst_1_n18 ), .A2(
        SubCellInst2_LFInst_7_LFInst_1_n17 ), .ZN(MCInst2_MC2_v2_0 [2]) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_1_U11  ( .A1(SubCellInput[29]), .A2(
        SubCellInst2_LFInst_7_LFInst_1_n16 ), .ZN(
        SubCellInst2_LFInst_7_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst2_LFInst_7_LFInst_1_U10  ( .A1(SubCellInput[31]), .A2(
        SubCellInst2_LFInst_7_LFInst_1_n15 ), .ZN(
        SubCellInst2_LFInst_7_LFInst_1_n16 ) );
  AND2_X1 SubCellInst2_LFInst_7_LFInst_1_U9  ( .A1(SubCellInput[28]), .A2(
        SubCellInput[30]), .ZN(SubCellInst2_LFInst_7_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_1_U8  ( .A1(SubCellInput[31]), .A2(
        SubCellInst2_LFInst_7_LFInst_1_n14 ), .ZN(
        SubCellInst2_LFInst_7_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_1_U7  ( .A1(
        SubCellInst2_LFInst_7_LFInst_1_n13 ), .A2(
        SubCellInst2_LFInst_7_LFInst_1_n12 ), .ZN(
        SubCellInst2_LFInst_7_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_1_U6  ( .A1(SubCellInput[28]), .A2(
        SubCellInput[30]), .ZN(SubCellInst2_LFInst_7_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_1_U5  ( .A1(
        SubCellInst2_LFInst_7_LFInst_1_n11 ), .A2(
        SubCellInst2_LFInst_7_LFInst_1_n10 ), .ZN(
        SubCellInst2_LFInst_7_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_1_U4  ( .A1(SubCellInput[28]), .A2(
        SubCellInput[29]), .ZN(SubCellInst2_LFInst_7_LFInst_1_n10 ) );
  INV_X1 SubCellInst2_LFInst_7_LFInst_1_U3  ( .A(SubCellInput[30]), .ZN(
        SubCellInst2_LFInst_7_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_2_U11  ( .A1(
        SubCellInst2_LFInst_7_LFInst_2_n22 ), .A2(
        SubCellInst2_LFInst_7_LFInst_2_n21 ), .ZN(MCInst2_MC2_v2_0 [3]) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_2_U10  ( .A1(SubCellInput[30]), .A2(
        SubCellInst2_LFInst_7_LFInst_2_n20 ), .ZN(
        SubCellInst2_LFInst_7_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst2_LFInst_7_LFInst_2_U9  ( .A1(SubCellInput[29]), .A2(
        SubCellInst2_LFInst_7_LFInst_2_n19 ), .ZN(
        SubCellInst2_LFInst_7_LFInst_2_n20 ) );
  INV_X1 SubCellInst2_LFInst_7_LFInst_2_U8  ( .A(SubCellInput[31]), .ZN(
        SubCellInst2_LFInst_7_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_2_U7  ( .A1(
        SubCellInst2_LFInst_7_LFInst_2_n18 ), .A2(
        SubCellInst2_LFInst_7_LFInst_2_n17 ), .ZN(
        SubCellInst2_LFInst_7_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst2_LFInst_7_LFInst_2_U6  ( .A(
        SubCellInst2_LFInst_7_LFInst_2_n16 ), .B(SubCellInput[30]), .Z(
        SubCellInst2_LFInst_7_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_2_U5  ( .A1(SubCellInput[28]), .A2(
        SubCellInput[29]), .ZN(SubCellInst2_LFInst_7_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_2_U4  ( .A1(
        SubCellInst2_LFInst_7_LFInst_2_n15 ), .A2(SubCellInput[31]), .ZN(
        SubCellInst2_LFInst_7_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst2_LFInst_7_LFInst_2_U3  ( .A(SubCellInput[28]), .B(
        SubCellInput[29]), .ZN(SubCellInst2_LFInst_7_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_3_U9  ( .A1(
        SubCellInst2_LFInst_7_LFInst_3_n16 ), .A2(
        SubCellInst2_LFInst_7_LFInst_3_n15 ), .ZN(MCInst2_MC2_v2_0 [0]) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_3_U8  ( .A1(SubCellInput[29]), .A2(
        SubCellInst2_LFInst_7_LFInst_3_n14 ), .ZN(
        SubCellInst2_LFInst_7_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst2_LFInst_7_LFInst_3_U7  ( .A(SubCellInput[31]), .B(
        SubCellInput[30]), .Z(SubCellInst2_LFInst_7_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_3_U6  ( .A1(
        SubCellInst2_LFInst_7_LFInst_3_n13 ), .A2(
        SubCellInst2_LFInst_7_LFInst_3_n12 ), .ZN(
        SubCellInst2_LFInst_7_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_7_LFInst_3_U5  ( .A1(SubCellInput[28]), .A2(
        SubCellInput[30]), .ZN(SubCellInst2_LFInst_7_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst2_LFInst_7_LFInst_3_U4  ( .A(SubCellInput[28]), .B(
        SubCellInst2_LFInst_7_LFInst_3_n11 ), .ZN(
        SubCellInst2_LFInst_7_LFInst_3_n13 ) );
  OR2_X1 SubCellInst2_LFInst_7_LFInst_3_U3  ( .A1(SubCellInput[31]), .A2(
        SubCellInput[29]), .ZN(SubCellInst2_LFInst_7_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_0_U6  ( .A1(SubCellInput[34]), .A2(
        SubCellInst2_LFInst_8_LFInst_0_n4 ), .ZN(
        SubCellInst2_LFInst_8_LFInst_0_n5 ) );
  INV_X1 SubCellInst2_LFInst_8_LFInst_0_U5  ( .A(SubCellInput[33]), .ZN(
        SubCellInst2_LFInst_8_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst2_LFInst_8_LFInst_0_U4  ( .A(SubCellInput[32]), .B(
        SubCellInput[35]), .Z(SubCellInst2_LFInst_8_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst2_LFInst_8_LFInst_0_U3  ( .A(
        SubCellInst2_LFInst_8_LFInst_0_n6 ), .B(
        SubCellInst2_LFInst_8_LFInst_0_n5 ), .ZN(MCInst2_MC2_v1_0 [0]) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_1_U12  ( .A1(
        SubCellInst2_LFInst_8_LFInst_1_n18 ), .A2(
        SubCellInst2_LFInst_8_LFInst_1_n17 ), .ZN(MCInst2_MC2_v1_3 [2]) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_1_U11  ( .A1(SubCellInput[33]), .A2(
        SubCellInst2_LFInst_8_LFInst_1_n16 ), .ZN(
        SubCellInst2_LFInst_8_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst2_LFInst_8_LFInst_1_U10  ( .A1(SubCellInput[35]), .A2(
        SubCellInst2_LFInst_8_LFInst_1_n15 ), .ZN(
        SubCellInst2_LFInst_8_LFInst_1_n16 ) );
  AND2_X1 SubCellInst2_LFInst_8_LFInst_1_U9  ( .A1(SubCellInput[32]), .A2(
        SubCellInput[34]), .ZN(SubCellInst2_LFInst_8_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_1_U8  ( .A1(SubCellInput[35]), .A2(
        SubCellInst2_LFInst_8_LFInst_1_n14 ), .ZN(
        SubCellInst2_LFInst_8_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_1_U7  ( .A1(
        SubCellInst2_LFInst_8_LFInst_1_n13 ), .A2(
        SubCellInst2_LFInst_8_LFInst_1_n12 ), .ZN(
        SubCellInst2_LFInst_8_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_1_U6  ( .A1(SubCellInput[32]), .A2(
        SubCellInput[34]), .ZN(SubCellInst2_LFInst_8_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_1_U5  ( .A1(
        SubCellInst2_LFInst_8_LFInst_1_n11 ), .A2(
        SubCellInst2_LFInst_8_LFInst_1_n10 ), .ZN(
        SubCellInst2_LFInst_8_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_1_U4  ( .A1(SubCellInput[32]), .A2(
        SubCellInput[33]), .ZN(SubCellInst2_LFInst_8_LFInst_1_n10 ) );
  INV_X1 SubCellInst2_LFInst_8_LFInst_1_U3  ( .A(SubCellInput[34]), .ZN(
        SubCellInst2_LFInst_8_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_2_U11  ( .A1(
        SubCellInst2_LFInst_8_LFInst_2_n22 ), .A2(
        SubCellInst2_LFInst_8_LFInst_2_n21 ), .ZN(Red_MCInst2_MC2_v1_1[0] )
         );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_2_U10  ( .A1(SubCellInput[34]), .A2(
        SubCellInst2_LFInst_8_LFInst_2_n20 ), .ZN(
        SubCellInst2_LFInst_8_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst2_LFInst_8_LFInst_2_U9  ( .A1(SubCellInput[33]), .A2(
        SubCellInst2_LFInst_8_LFInst_2_n19 ), .ZN(
        SubCellInst2_LFInst_8_LFInst_2_n20 ) );
  INV_X1 SubCellInst2_LFInst_8_LFInst_2_U8  ( .A(SubCellInput[35]), .ZN(
        SubCellInst2_LFInst_8_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_2_U7  ( .A1(
        SubCellInst2_LFInst_8_LFInst_2_n18 ), .A2(
        SubCellInst2_LFInst_8_LFInst_2_n17 ), .ZN(
        SubCellInst2_LFInst_8_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst2_LFInst_8_LFInst_2_U6  ( .A(
        SubCellInst2_LFInst_8_LFInst_2_n16 ), .B(SubCellInput[34]), .Z(
        SubCellInst2_LFInst_8_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_2_U5  ( .A1(SubCellInput[32]), .A2(
        SubCellInput[33]), .ZN(SubCellInst2_LFInst_8_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_2_U4  ( .A1(
        SubCellInst2_LFInst_8_LFInst_2_n15 ), .A2(SubCellInput[35]), .ZN(
        SubCellInst2_LFInst_8_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst2_LFInst_8_LFInst_2_U3  ( .A(SubCellInput[32]), .B(
        SubCellInput[33]), .ZN(SubCellInst2_LFInst_8_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_3_U9  ( .A1(
        SubCellInst2_LFInst_8_LFInst_3_n16 ), .A2(
        SubCellInst2_LFInst_8_LFInst_3_n15 ), .ZN(MCInst2_MC2_v1_0 [3]) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_3_U8  ( .A1(SubCellInput[33]), .A2(
        SubCellInst2_LFInst_8_LFInst_3_n14 ), .ZN(
        SubCellInst2_LFInst_8_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst2_LFInst_8_LFInst_3_U7  ( .A(SubCellInput[35]), .B(
        SubCellInput[34]), .Z(SubCellInst2_LFInst_8_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_3_U6  ( .A1(
        SubCellInst2_LFInst_8_LFInst_3_n13 ), .A2(
        SubCellInst2_LFInst_8_LFInst_3_n12 ), .ZN(
        SubCellInst2_LFInst_8_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_8_LFInst_3_U5  ( .A1(SubCellInput[32]), .A2(
        SubCellInput[34]), .ZN(SubCellInst2_LFInst_8_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst2_LFInst_8_LFInst_3_U4  ( .A(SubCellInput[32]), .B(
        SubCellInst2_LFInst_8_LFInst_3_n11 ), .ZN(
        SubCellInst2_LFInst_8_LFInst_3_n13 ) );
  OR2_X1 SubCellInst2_LFInst_8_LFInst_3_U3  ( .A1(SubCellInput[35]), .A2(
        SubCellInput[33]), .ZN(SubCellInst2_LFInst_8_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_0_U6  ( .A1(SubCellInput[38]), .A2(
        SubCellInst2_LFInst_9_LFInst_0_n4 ), .ZN(
        SubCellInst2_LFInst_9_LFInst_0_n5 ) );
  INV_X1 SubCellInst2_LFInst_9_LFInst_0_U5  ( .A(SubCellInput[37]), .ZN(
        SubCellInst2_LFInst_9_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst2_LFInst_9_LFInst_0_U4  ( .A(SubCellInput[36]), .B(
        SubCellInput[39]), .Z(SubCellInst2_LFInst_9_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst2_LFInst_9_LFInst_0_U3  ( .A(
        SubCellInst2_LFInst_9_LFInst_0_n6 ), .B(
        SubCellInst2_LFInst_9_LFInst_0_n5 ), .ZN(MCInst2_MC1_v1_0 [0]) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_1_U12  ( .A1(
        SubCellInst2_LFInst_9_LFInst_1_n18 ), .A2(
        SubCellInst2_LFInst_9_LFInst_1_n17 ), .ZN(MCInst2_MC1_v1_3 [2]) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_1_U11  ( .A1(SubCellInput[37]), .A2(
        SubCellInst2_LFInst_9_LFInst_1_n16 ), .ZN(
        SubCellInst2_LFInst_9_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst2_LFInst_9_LFInst_1_U10  ( .A1(SubCellInput[39]), .A2(
        SubCellInst2_LFInst_9_LFInst_1_n15 ), .ZN(
        SubCellInst2_LFInst_9_LFInst_1_n16 ) );
  AND2_X1 SubCellInst2_LFInst_9_LFInst_1_U9  ( .A1(SubCellInput[36]), .A2(
        SubCellInput[38]), .ZN(SubCellInst2_LFInst_9_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_1_U8  ( .A1(SubCellInput[39]), .A2(
        SubCellInst2_LFInst_9_LFInst_1_n14 ), .ZN(
        SubCellInst2_LFInst_9_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_1_U7  ( .A1(
        SubCellInst2_LFInst_9_LFInst_1_n13 ), .A2(
        SubCellInst2_LFInst_9_LFInst_1_n12 ), .ZN(
        SubCellInst2_LFInst_9_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_1_U6  ( .A1(SubCellInput[36]), .A2(
        SubCellInput[38]), .ZN(SubCellInst2_LFInst_9_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_1_U5  ( .A1(
        SubCellInst2_LFInst_9_LFInst_1_n11 ), .A2(
        SubCellInst2_LFInst_9_LFInst_1_n10 ), .ZN(
        SubCellInst2_LFInst_9_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_1_U4  ( .A1(SubCellInput[36]), .A2(
        SubCellInput[37]), .ZN(SubCellInst2_LFInst_9_LFInst_1_n10 ) );
  INV_X1 SubCellInst2_LFInst_9_LFInst_1_U3  ( .A(SubCellInput[38]), .ZN(
        SubCellInst2_LFInst_9_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_2_U11  ( .A1(
        SubCellInst2_LFInst_9_LFInst_2_n22 ), .A2(
        SubCellInst2_LFInst_9_LFInst_2_n21 ), .ZN(Red_MCInst2_MC1_v1_1[0] )
         );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_2_U10  ( .A1(SubCellInput[38]), .A2(
        SubCellInst2_LFInst_9_LFInst_2_n20 ), .ZN(
        SubCellInst2_LFInst_9_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst2_LFInst_9_LFInst_2_U9  ( .A1(SubCellInput[37]), .A2(
        SubCellInst2_LFInst_9_LFInst_2_n19 ), .ZN(
        SubCellInst2_LFInst_9_LFInst_2_n20 ) );
  INV_X1 SubCellInst2_LFInst_9_LFInst_2_U8  ( .A(SubCellInput[39]), .ZN(
        SubCellInst2_LFInst_9_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_2_U7  ( .A1(
        SubCellInst2_LFInst_9_LFInst_2_n18 ), .A2(
        SubCellInst2_LFInst_9_LFInst_2_n17 ), .ZN(
        SubCellInst2_LFInst_9_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst2_LFInst_9_LFInst_2_U6  ( .A(
        SubCellInst2_LFInst_9_LFInst_2_n16 ), .B(SubCellInput[38]), .Z(
        SubCellInst2_LFInst_9_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_2_U5  ( .A1(SubCellInput[36]), .A2(
        SubCellInput[37]), .ZN(SubCellInst2_LFInst_9_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_2_U4  ( .A1(
        SubCellInst2_LFInst_9_LFInst_2_n15 ), .A2(SubCellInput[39]), .ZN(
        SubCellInst2_LFInst_9_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst2_LFInst_9_LFInst_2_U3  ( .A(SubCellInput[36]), .B(
        SubCellInput[37]), .ZN(SubCellInst2_LFInst_9_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_3_U9  ( .A1(
        SubCellInst2_LFInst_9_LFInst_3_n16 ), .A2(
        SubCellInst2_LFInst_9_LFInst_3_n15 ), .ZN(MCInst2_MC1_v1_0 [3]) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_3_U8  ( .A1(SubCellInput[37]), .A2(
        SubCellInst2_LFInst_9_LFInst_3_n14 ), .ZN(
        SubCellInst2_LFInst_9_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst2_LFInst_9_LFInst_3_U7  ( .A(SubCellInput[39]), .B(
        SubCellInput[38]), .Z(SubCellInst2_LFInst_9_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_3_U6  ( .A1(
        SubCellInst2_LFInst_9_LFInst_3_n13 ), .A2(
        SubCellInst2_LFInst_9_LFInst_3_n12 ), .ZN(
        SubCellInst2_LFInst_9_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_9_LFInst_3_U5  ( .A1(SubCellInput[36]), .A2(
        SubCellInput[38]), .ZN(SubCellInst2_LFInst_9_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst2_LFInst_9_LFInst_3_U4  ( .A(SubCellInput[36]), .B(
        SubCellInst2_LFInst_9_LFInst_3_n11 ), .ZN(
        SubCellInst2_LFInst_9_LFInst_3_n13 ) );
  OR2_X1 SubCellInst2_LFInst_9_LFInst_3_U3  ( .A1(SubCellInput[39]), .A2(
        SubCellInput[37]), .ZN(SubCellInst2_LFInst_9_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_0_U6  ( .A1(SubCellInput[42]), .A2(
        SubCellInst2_LFInst_10_LFInst_0_n4 ), .ZN(
        SubCellInst2_LFInst_10_LFInst_0_n5 ) );
  INV_X1 SubCellInst2_LFInst_10_LFInst_0_U5  ( .A(SubCellInput[41]), .ZN(
        SubCellInst2_LFInst_10_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst2_LFInst_10_LFInst_0_U4  ( .A(SubCellInput[40]), .B(
        SubCellInput[43]), .Z(SubCellInst2_LFInst_10_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst2_LFInst_10_LFInst_0_U3  ( .A(
        SubCellInst2_LFInst_10_LFInst_0_n6 ), .B(
        SubCellInst2_LFInst_10_LFInst_0_n5 ), .ZN(MCInst2_MC0_v1_0 [0]) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_1_U12  ( .A1(
        SubCellInst2_LFInst_10_LFInst_1_n18 ), .A2(
        SubCellInst2_LFInst_10_LFInst_1_n17 ), .ZN(MCInst2_MC0_v1_3 [2]) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_1_U11  ( .A1(SubCellInput[41]), .A2(
        SubCellInst2_LFInst_10_LFInst_1_n16 ), .ZN(
        SubCellInst2_LFInst_10_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst2_LFInst_10_LFInst_1_U10  ( .A1(SubCellInput[43]), .A2(
        SubCellInst2_LFInst_10_LFInst_1_n15 ), .ZN(
        SubCellInst2_LFInst_10_LFInst_1_n16 ) );
  AND2_X1 SubCellInst2_LFInst_10_LFInst_1_U9  ( .A1(SubCellInput[40]), .A2(
        SubCellInput[42]), .ZN(SubCellInst2_LFInst_10_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_1_U8  ( .A1(SubCellInput[43]), .A2(
        SubCellInst2_LFInst_10_LFInst_1_n14 ), .ZN(
        SubCellInst2_LFInst_10_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_1_U7  ( .A1(
        SubCellInst2_LFInst_10_LFInst_1_n13 ), .A2(
        SubCellInst2_LFInst_10_LFInst_1_n12 ), .ZN(
        SubCellInst2_LFInst_10_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_1_U6  ( .A1(SubCellInput[40]), .A2(
        SubCellInput[42]), .ZN(SubCellInst2_LFInst_10_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_1_U5  ( .A1(
        SubCellInst2_LFInst_10_LFInst_1_n11 ), .A2(
        SubCellInst2_LFInst_10_LFInst_1_n10 ), .ZN(
        SubCellInst2_LFInst_10_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_1_U4  ( .A1(SubCellInput[40]), .A2(
        SubCellInput[41]), .ZN(SubCellInst2_LFInst_10_LFInst_1_n10 ) );
  INV_X1 SubCellInst2_LFInst_10_LFInst_1_U3  ( .A(SubCellInput[42]), .ZN(
        SubCellInst2_LFInst_10_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_2_U11  ( .A1(
        SubCellInst2_LFInst_10_LFInst_2_n22 ), .A2(
        SubCellInst2_LFInst_10_LFInst_2_n21 ), .ZN(Red_MCInst2_MC0_v1_1[0] )
         );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_2_U10  ( .A1(SubCellInput[42]), .A2(
        SubCellInst2_LFInst_10_LFInst_2_n20 ), .ZN(
        SubCellInst2_LFInst_10_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst2_LFInst_10_LFInst_2_U9  ( .A1(SubCellInput[41]), .A2(
        SubCellInst2_LFInst_10_LFInst_2_n19 ), .ZN(
        SubCellInst2_LFInst_10_LFInst_2_n20 ) );
  INV_X1 SubCellInst2_LFInst_10_LFInst_2_U8  ( .A(SubCellInput[43]), .ZN(
        SubCellInst2_LFInst_10_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_2_U7  ( .A1(
        SubCellInst2_LFInst_10_LFInst_2_n18 ), .A2(
        SubCellInst2_LFInst_10_LFInst_2_n17 ), .ZN(
        SubCellInst2_LFInst_10_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst2_LFInst_10_LFInst_2_U6  ( .A(
        SubCellInst2_LFInst_10_LFInst_2_n16 ), .B(SubCellInput[42]), .Z(
        SubCellInst2_LFInst_10_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_2_U5  ( .A1(SubCellInput[40]), .A2(
        SubCellInput[41]), .ZN(SubCellInst2_LFInst_10_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_2_U4  ( .A1(
        SubCellInst2_LFInst_10_LFInst_2_n15 ), .A2(SubCellInput[43]), .ZN(
        SubCellInst2_LFInst_10_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst2_LFInst_10_LFInst_2_U3  ( .A(SubCellInput[40]), .B(
        SubCellInput[41]), .ZN(SubCellInst2_LFInst_10_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_3_U9  ( .A1(
        SubCellInst2_LFInst_10_LFInst_3_n16 ), .A2(
        SubCellInst2_LFInst_10_LFInst_3_n15 ), .ZN(MCInst2_MC0_v1_0 [3]) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_3_U8  ( .A1(SubCellInput[41]), .A2(
        SubCellInst2_LFInst_10_LFInst_3_n14 ), .ZN(
        SubCellInst2_LFInst_10_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst2_LFInst_10_LFInst_3_U7  ( .A(SubCellInput[43]), .B(
        SubCellInput[42]), .Z(SubCellInst2_LFInst_10_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_3_U6  ( .A1(
        SubCellInst2_LFInst_10_LFInst_3_n13 ), .A2(
        SubCellInst2_LFInst_10_LFInst_3_n12 ), .ZN(
        SubCellInst2_LFInst_10_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_10_LFInst_3_U5  ( .A1(SubCellInput[40]), .A2(
        SubCellInput[42]), .ZN(SubCellInst2_LFInst_10_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst2_LFInst_10_LFInst_3_U4  ( .A(SubCellInput[40]), .B(
        SubCellInst2_LFInst_10_LFInst_3_n11 ), .ZN(
        SubCellInst2_LFInst_10_LFInst_3_n13 ) );
  OR2_X1 SubCellInst2_LFInst_10_LFInst_3_U3  ( .A1(SubCellInput[43]), .A2(
        SubCellInput[41]), .ZN(SubCellInst2_LFInst_10_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_0_U6  ( .A1(SubCellInput[46]), .A2(
        SubCellInst2_LFInst_11_LFInst_0_n4 ), .ZN(
        SubCellInst2_LFInst_11_LFInst_0_n5 ) );
  INV_X1 SubCellInst2_LFInst_11_LFInst_0_U5  ( .A(SubCellInput[45]), .ZN(
        SubCellInst2_LFInst_11_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst2_LFInst_11_LFInst_0_U4  ( .A(SubCellInput[44]), .B(
        SubCellInput[47]), .Z(SubCellInst2_LFInst_11_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst2_LFInst_11_LFInst_0_U3  ( .A(
        SubCellInst2_LFInst_11_LFInst_0_n6 ), .B(
        SubCellInst2_LFInst_11_LFInst_0_n5 ), .ZN(MCInst2_MC3_v1_0 [0]) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_1_U12  ( .A1(
        SubCellInst2_LFInst_11_LFInst_1_n18 ), .A2(
        SubCellInst2_LFInst_11_LFInst_1_n17 ), .ZN(MCInst2_MC3_v1_3 [2]) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_1_U11  ( .A1(SubCellInput[45]), .A2(
        SubCellInst2_LFInst_11_LFInst_1_n16 ), .ZN(
        SubCellInst2_LFInst_11_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst2_LFInst_11_LFInst_1_U10  ( .A1(SubCellInput[47]), .A2(
        SubCellInst2_LFInst_11_LFInst_1_n15 ), .ZN(
        SubCellInst2_LFInst_11_LFInst_1_n16 ) );
  AND2_X1 SubCellInst2_LFInst_11_LFInst_1_U9  ( .A1(SubCellInput[44]), .A2(
        SubCellInput[46]), .ZN(SubCellInst2_LFInst_11_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_1_U8  ( .A1(SubCellInput[47]), .A2(
        SubCellInst2_LFInst_11_LFInst_1_n14 ), .ZN(
        SubCellInst2_LFInst_11_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_1_U7  ( .A1(
        SubCellInst2_LFInst_11_LFInst_1_n13 ), .A2(
        SubCellInst2_LFInst_11_LFInst_1_n12 ), .ZN(
        SubCellInst2_LFInst_11_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_1_U6  ( .A1(SubCellInput[44]), .A2(
        SubCellInput[46]), .ZN(SubCellInst2_LFInst_11_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_1_U5  ( .A1(
        SubCellInst2_LFInst_11_LFInst_1_n11 ), .A2(
        SubCellInst2_LFInst_11_LFInst_1_n10 ), .ZN(
        SubCellInst2_LFInst_11_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_1_U4  ( .A1(SubCellInput[44]), .A2(
        SubCellInput[45]), .ZN(SubCellInst2_LFInst_11_LFInst_1_n10 ) );
  INV_X1 SubCellInst2_LFInst_11_LFInst_1_U3  ( .A(SubCellInput[46]), .ZN(
        SubCellInst2_LFInst_11_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_2_U11  ( .A1(
        SubCellInst2_LFInst_11_LFInst_2_n22 ), .A2(
        SubCellInst2_LFInst_11_LFInst_2_n21 ), .ZN(Red_MCInst2_MC3_v1_1[0] )
         );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_2_U10  ( .A1(SubCellInput[46]), .A2(
        SubCellInst2_LFInst_11_LFInst_2_n20 ), .ZN(
        SubCellInst2_LFInst_11_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst2_LFInst_11_LFInst_2_U9  ( .A1(SubCellInput[45]), .A2(
        SubCellInst2_LFInst_11_LFInst_2_n19 ), .ZN(
        SubCellInst2_LFInst_11_LFInst_2_n20 ) );
  INV_X1 SubCellInst2_LFInst_11_LFInst_2_U8  ( .A(SubCellInput[47]), .ZN(
        SubCellInst2_LFInst_11_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_2_U7  ( .A1(
        SubCellInst2_LFInst_11_LFInst_2_n18 ), .A2(
        SubCellInst2_LFInst_11_LFInst_2_n17 ), .ZN(
        SubCellInst2_LFInst_11_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst2_LFInst_11_LFInst_2_U6  ( .A(
        SubCellInst2_LFInst_11_LFInst_2_n16 ), .B(SubCellInput[46]), .Z(
        SubCellInst2_LFInst_11_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_2_U5  ( .A1(SubCellInput[44]), .A2(
        SubCellInput[45]), .ZN(SubCellInst2_LFInst_11_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_2_U4  ( .A1(
        SubCellInst2_LFInst_11_LFInst_2_n15 ), .A2(SubCellInput[47]), .ZN(
        SubCellInst2_LFInst_11_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst2_LFInst_11_LFInst_2_U3  ( .A(SubCellInput[44]), .B(
        SubCellInput[45]), .ZN(SubCellInst2_LFInst_11_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_3_U9  ( .A1(
        SubCellInst2_LFInst_11_LFInst_3_n16 ), .A2(
        SubCellInst2_LFInst_11_LFInst_3_n15 ), .ZN(MCInst2_MC3_v1_0 [3]) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_3_U8  ( .A1(SubCellInput[45]), .A2(
        SubCellInst2_LFInst_11_LFInst_3_n14 ), .ZN(
        SubCellInst2_LFInst_11_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst2_LFInst_11_LFInst_3_U7  ( .A(SubCellInput[47]), .B(
        SubCellInput[46]), .Z(SubCellInst2_LFInst_11_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_3_U6  ( .A1(
        SubCellInst2_LFInst_11_LFInst_3_n13 ), .A2(
        SubCellInst2_LFInst_11_LFInst_3_n12 ), .ZN(
        SubCellInst2_LFInst_11_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_11_LFInst_3_U5  ( .A1(SubCellInput[44]), .A2(
        SubCellInput[46]), .ZN(SubCellInst2_LFInst_11_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst2_LFInst_11_LFInst_3_U4  ( .A(SubCellInput[44]), .B(
        SubCellInst2_LFInst_11_LFInst_3_n11 ), .ZN(
        SubCellInst2_LFInst_11_LFInst_3_n13 ) );
  OR2_X1 SubCellInst2_LFInst_11_LFInst_3_U3  ( .A1(SubCellInput[47]), .A2(
        SubCellInput[45]), .ZN(SubCellInst2_LFInst_11_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_0_U6  ( .A1(SubCellInput[50]), .A2(
        SubCellInst2_LFInst_12_LFInst_0_n4 ), .ZN(
        SubCellInst2_LFInst_12_LFInst_0_n5 ) );
  INV_X1 SubCellInst2_LFInst_12_LFInst_0_U5  ( .A(SubCellInput[49]), .ZN(
        SubCellInst2_LFInst_12_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst2_LFInst_12_LFInst_0_U4  ( .A(SubCellInput[48]), .B(
        SubCellInput[51]), .Z(SubCellInst2_LFInst_12_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst2_LFInst_12_LFInst_0_U3  ( .A(
        SubCellInst2_LFInst_12_LFInst_0_n6 ), .B(
        SubCellInst2_LFInst_12_LFInst_0_n5 ), .ZN(Red_MCInst2_MC3_v0_1[0] )
         );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_1_U12  ( .A1(
        SubCellInst2_LFInst_12_LFInst_1_n18 ), .A2(
        SubCellInst2_LFInst_12_LFInst_1_n17 ), .ZN(MCInst2_MC3_v0_0 [3]) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_1_U11  ( .A1(SubCellInput[49]), .A2(
        SubCellInst2_LFInst_12_LFInst_1_n16 ), .ZN(
        SubCellInst2_LFInst_12_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst2_LFInst_12_LFInst_1_U10  ( .A1(SubCellInput[51]), .A2(
        SubCellInst2_LFInst_12_LFInst_1_n15 ), .ZN(
        SubCellInst2_LFInst_12_LFInst_1_n16 ) );
  AND2_X1 SubCellInst2_LFInst_12_LFInst_1_U9  ( .A1(SubCellInput[48]), .A2(
        SubCellInput[50]), .ZN(SubCellInst2_LFInst_12_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_1_U8  ( .A1(SubCellInput[51]), .A2(
        SubCellInst2_LFInst_12_LFInst_1_n14 ), .ZN(
        SubCellInst2_LFInst_12_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_1_U7  ( .A1(
        SubCellInst2_LFInst_12_LFInst_1_n13 ), .A2(
        SubCellInst2_LFInst_12_LFInst_1_n12 ), .ZN(
        SubCellInst2_LFInst_12_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_1_U6  ( .A1(SubCellInput[48]), .A2(
        SubCellInput[50]), .ZN(SubCellInst2_LFInst_12_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_1_U5  ( .A1(
        SubCellInst2_LFInst_12_LFInst_1_n11 ), .A2(
        SubCellInst2_LFInst_12_LFInst_1_n10 ), .ZN(
        SubCellInst2_LFInst_12_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_1_U4  ( .A1(SubCellInput[48]), .A2(
        SubCellInput[49]), .ZN(SubCellInst2_LFInst_12_LFInst_1_n10 ) );
  INV_X1 SubCellInst2_LFInst_12_LFInst_1_U3  ( .A(SubCellInput[50]), .ZN(
        SubCellInst2_LFInst_12_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_2_U11  ( .A1(
        SubCellInst2_LFInst_12_LFInst_2_n22 ), .A2(
        SubCellInst2_LFInst_12_LFInst_2_n21 ), .ZN(MCInst2_MC3_v0_3 [3]) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_2_U10  ( .A1(SubCellInput[50]), .A2(
        SubCellInst2_LFInst_12_LFInst_2_n20 ), .ZN(
        SubCellInst2_LFInst_12_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst2_LFInst_12_LFInst_2_U9  ( .A1(SubCellInput[49]), .A2(
        SubCellInst2_LFInst_12_LFInst_2_n19 ), .ZN(
        SubCellInst2_LFInst_12_LFInst_2_n20 ) );
  INV_X1 SubCellInst2_LFInst_12_LFInst_2_U8  ( .A(SubCellInput[51]), .ZN(
        SubCellInst2_LFInst_12_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_2_U7  ( .A1(
        SubCellInst2_LFInst_12_LFInst_2_n18 ), .A2(
        SubCellInst2_LFInst_12_LFInst_2_n17 ), .ZN(
        SubCellInst2_LFInst_12_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst2_LFInst_12_LFInst_2_U6  ( .A(
        SubCellInst2_LFInst_12_LFInst_2_n16 ), .B(SubCellInput[50]), .Z(
        SubCellInst2_LFInst_12_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_2_U5  ( .A1(SubCellInput[48]), .A2(
        SubCellInput[49]), .ZN(SubCellInst2_LFInst_12_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_2_U4  ( .A1(
        SubCellInst2_LFInst_12_LFInst_2_n15 ), .A2(SubCellInput[51]), .ZN(
        SubCellInst2_LFInst_12_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst2_LFInst_12_LFInst_2_U3  ( .A(SubCellInput[48]), .B(
        SubCellInput[49]), .ZN(SubCellInst2_LFInst_12_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_3_U9  ( .A1(
        SubCellInst2_LFInst_12_LFInst_3_n16 ), .A2(
        SubCellInst2_LFInst_12_LFInst_3_n15 ), .ZN(MCInst2_MC3_v0_3 [0]) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_3_U8  ( .A1(SubCellInput[49]), .A2(
        SubCellInst2_LFInst_12_LFInst_3_n14 ), .ZN(
        SubCellInst2_LFInst_12_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst2_LFInst_12_LFInst_3_U7  ( .A(SubCellInput[51]), .B(
        SubCellInput[50]), .Z(SubCellInst2_LFInst_12_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_3_U6  ( .A1(
        SubCellInst2_LFInst_12_LFInst_3_n13 ), .A2(
        SubCellInst2_LFInst_12_LFInst_3_n12 ), .ZN(
        SubCellInst2_LFInst_12_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_12_LFInst_3_U5  ( .A1(SubCellInput[48]), .A2(
        SubCellInput[50]), .ZN(SubCellInst2_LFInst_12_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst2_LFInst_12_LFInst_3_U4  ( .A(SubCellInput[48]), .B(
        SubCellInst2_LFInst_12_LFInst_3_n11 ), .ZN(
        SubCellInst2_LFInst_12_LFInst_3_n13 ) );
  OR2_X1 SubCellInst2_LFInst_12_LFInst_3_U3  ( .A1(SubCellInput[51]), .A2(
        SubCellInput[49]), .ZN(SubCellInst2_LFInst_12_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_0_U6  ( .A1(SubCellInput[54]), .A2(
        SubCellInst2_LFInst_13_LFInst_0_n4 ), .ZN(
        SubCellInst2_LFInst_13_LFInst_0_n5 ) );
  INV_X1 SubCellInst2_LFInst_13_LFInst_0_U5  ( .A(SubCellInput[53]), .ZN(
        SubCellInst2_LFInst_13_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst2_LFInst_13_LFInst_0_U4  ( .A(SubCellInput[52]), .B(
        SubCellInput[55]), .Z(SubCellInst2_LFInst_13_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst2_LFInst_13_LFInst_0_U3  ( .A(
        SubCellInst2_LFInst_13_LFInst_0_n6 ), .B(
        SubCellInst2_LFInst_13_LFInst_0_n5 ), .ZN(Red_MCInst2_MC2_v0_1[0] )
         );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_1_U12  ( .A1(
        SubCellInst2_LFInst_13_LFInst_1_n18 ), .A2(
        SubCellInst2_LFInst_13_LFInst_1_n17 ), .ZN(MCInst2_MC2_v0_0 [3]) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_1_U11  ( .A1(SubCellInput[53]), .A2(
        SubCellInst2_LFInst_13_LFInst_1_n16 ), .ZN(
        SubCellInst2_LFInst_13_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst2_LFInst_13_LFInst_1_U10  ( .A1(SubCellInput[55]), .A2(
        SubCellInst2_LFInst_13_LFInst_1_n15 ), .ZN(
        SubCellInst2_LFInst_13_LFInst_1_n16 ) );
  AND2_X1 SubCellInst2_LFInst_13_LFInst_1_U9  ( .A1(SubCellInput[52]), .A2(
        SubCellInput[54]), .ZN(SubCellInst2_LFInst_13_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_1_U8  ( .A1(SubCellInput[55]), .A2(
        SubCellInst2_LFInst_13_LFInst_1_n14 ), .ZN(
        SubCellInst2_LFInst_13_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_1_U7  ( .A1(
        SubCellInst2_LFInst_13_LFInst_1_n13 ), .A2(
        SubCellInst2_LFInst_13_LFInst_1_n12 ), .ZN(
        SubCellInst2_LFInst_13_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_1_U6  ( .A1(SubCellInput[52]), .A2(
        SubCellInput[54]), .ZN(SubCellInst2_LFInst_13_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_1_U5  ( .A1(
        SubCellInst2_LFInst_13_LFInst_1_n11 ), .A2(
        SubCellInst2_LFInst_13_LFInst_1_n10 ), .ZN(
        SubCellInst2_LFInst_13_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_1_U4  ( .A1(SubCellInput[52]), .A2(
        SubCellInput[53]), .ZN(SubCellInst2_LFInst_13_LFInst_1_n10 ) );
  INV_X1 SubCellInst2_LFInst_13_LFInst_1_U3  ( .A(SubCellInput[54]), .ZN(
        SubCellInst2_LFInst_13_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_2_U11  ( .A1(
        SubCellInst2_LFInst_13_LFInst_2_n22 ), .A2(
        SubCellInst2_LFInst_13_LFInst_2_n21 ), .ZN(MCInst2_MC2_v0_3 [3]) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_2_U10  ( .A1(SubCellInput[54]), .A2(
        SubCellInst2_LFInst_13_LFInst_2_n20 ), .ZN(
        SubCellInst2_LFInst_13_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst2_LFInst_13_LFInst_2_U9  ( .A1(SubCellInput[53]), .A2(
        SubCellInst2_LFInst_13_LFInst_2_n19 ), .ZN(
        SubCellInst2_LFInst_13_LFInst_2_n20 ) );
  INV_X1 SubCellInst2_LFInst_13_LFInst_2_U8  ( .A(SubCellInput[55]), .ZN(
        SubCellInst2_LFInst_13_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_2_U7  ( .A1(
        SubCellInst2_LFInst_13_LFInst_2_n18 ), .A2(
        SubCellInst2_LFInst_13_LFInst_2_n17 ), .ZN(
        SubCellInst2_LFInst_13_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst2_LFInst_13_LFInst_2_U6  ( .A(
        SubCellInst2_LFInst_13_LFInst_2_n16 ), .B(SubCellInput[54]), .Z(
        SubCellInst2_LFInst_13_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_2_U5  ( .A1(SubCellInput[52]), .A2(
        SubCellInput[53]), .ZN(SubCellInst2_LFInst_13_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_2_U4  ( .A1(
        SubCellInst2_LFInst_13_LFInst_2_n15 ), .A2(SubCellInput[55]), .ZN(
        SubCellInst2_LFInst_13_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst2_LFInst_13_LFInst_2_U3  ( .A(SubCellInput[52]), .B(
        SubCellInput[53]), .ZN(SubCellInst2_LFInst_13_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_3_U9  ( .A1(
        SubCellInst2_LFInst_13_LFInst_3_n16 ), .A2(
        SubCellInst2_LFInst_13_LFInst_3_n15 ), .ZN(MCInst2_MC2_v0_3 [0]) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_3_U8  ( .A1(SubCellInput[53]), .A2(
        SubCellInst2_LFInst_13_LFInst_3_n14 ), .ZN(
        SubCellInst2_LFInst_13_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst2_LFInst_13_LFInst_3_U7  ( .A(SubCellInput[55]), .B(
        SubCellInput[54]), .Z(SubCellInst2_LFInst_13_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_3_U6  ( .A1(
        SubCellInst2_LFInst_13_LFInst_3_n13 ), .A2(
        SubCellInst2_LFInst_13_LFInst_3_n12 ), .ZN(
        SubCellInst2_LFInst_13_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_13_LFInst_3_U5  ( .A1(SubCellInput[52]), .A2(
        SubCellInput[54]), .ZN(SubCellInst2_LFInst_13_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst2_LFInst_13_LFInst_3_U4  ( .A(SubCellInput[52]), .B(
        SubCellInst2_LFInst_13_LFInst_3_n11 ), .ZN(
        SubCellInst2_LFInst_13_LFInst_3_n13 ) );
  OR2_X1 SubCellInst2_LFInst_13_LFInst_3_U3  ( .A1(SubCellInput[55]), .A2(
        SubCellInput[53]), .ZN(SubCellInst2_LFInst_13_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_0_U6  ( .A1(SubCellInput[58]), .A2(
        SubCellInst2_LFInst_14_LFInst_0_n4 ), .ZN(
        SubCellInst2_LFInst_14_LFInst_0_n5 ) );
  INV_X1 SubCellInst2_LFInst_14_LFInst_0_U5  ( .A(SubCellInput[57]), .ZN(
        SubCellInst2_LFInst_14_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst2_LFInst_14_LFInst_0_U4  ( .A(SubCellInput[56]), .B(
        SubCellInput[59]), .Z(SubCellInst2_LFInst_14_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst2_LFInst_14_LFInst_0_U3  ( .A(
        SubCellInst2_LFInst_14_LFInst_0_n6 ), .B(
        SubCellInst2_LFInst_14_LFInst_0_n5 ), .ZN(Red_MCInst2_MC1_v0_1[0] )
         );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_1_U12  ( .A1(
        SubCellInst2_LFInst_14_LFInst_1_n18 ), .A2(
        SubCellInst2_LFInst_14_LFInst_1_n17 ), .ZN(MCInst2_MC1_v0_0 [3]) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_1_U11  ( .A1(SubCellInput[57]), .A2(
        SubCellInst2_LFInst_14_LFInst_1_n16 ), .ZN(
        SubCellInst2_LFInst_14_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst2_LFInst_14_LFInst_1_U10  ( .A1(SubCellInput[59]), .A2(
        SubCellInst2_LFInst_14_LFInst_1_n15 ), .ZN(
        SubCellInst2_LFInst_14_LFInst_1_n16 ) );
  AND2_X1 SubCellInst2_LFInst_14_LFInst_1_U9  ( .A1(SubCellInput[56]), .A2(
        SubCellInput[58]), .ZN(SubCellInst2_LFInst_14_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_1_U8  ( .A1(SubCellInput[59]), .A2(
        SubCellInst2_LFInst_14_LFInst_1_n14 ), .ZN(
        SubCellInst2_LFInst_14_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_1_U7  ( .A1(
        SubCellInst2_LFInst_14_LFInst_1_n13 ), .A2(
        SubCellInst2_LFInst_14_LFInst_1_n12 ), .ZN(
        SubCellInst2_LFInst_14_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_1_U6  ( .A1(SubCellInput[56]), .A2(
        SubCellInput[58]), .ZN(SubCellInst2_LFInst_14_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_1_U5  ( .A1(
        SubCellInst2_LFInst_14_LFInst_1_n11 ), .A2(
        SubCellInst2_LFInst_14_LFInst_1_n10 ), .ZN(
        SubCellInst2_LFInst_14_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_1_U4  ( .A1(SubCellInput[56]), .A2(
        SubCellInput[57]), .ZN(SubCellInst2_LFInst_14_LFInst_1_n10 ) );
  INV_X1 SubCellInst2_LFInst_14_LFInst_1_U3  ( .A(SubCellInput[58]), .ZN(
        SubCellInst2_LFInst_14_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_2_U11  ( .A1(
        SubCellInst2_LFInst_14_LFInst_2_n22 ), .A2(
        SubCellInst2_LFInst_14_LFInst_2_n21 ), .ZN(MCInst2_MC1_v0_3 [3]) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_2_U10  ( .A1(SubCellInput[58]), .A2(
        SubCellInst2_LFInst_14_LFInst_2_n20 ), .ZN(
        SubCellInst2_LFInst_14_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst2_LFInst_14_LFInst_2_U9  ( .A1(SubCellInput[57]), .A2(
        SubCellInst2_LFInst_14_LFInst_2_n19 ), .ZN(
        SubCellInst2_LFInst_14_LFInst_2_n20 ) );
  INV_X1 SubCellInst2_LFInst_14_LFInst_2_U8  ( .A(SubCellInput[59]), .ZN(
        SubCellInst2_LFInst_14_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_2_U7  ( .A1(
        SubCellInst2_LFInst_14_LFInst_2_n18 ), .A2(
        SubCellInst2_LFInst_14_LFInst_2_n17 ), .ZN(
        SubCellInst2_LFInst_14_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst2_LFInst_14_LFInst_2_U6  ( .A(
        SubCellInst2_LFInst_14_LFInst_2_n16 ), .B(SubCellInput[58]), .Z(
        SubCellInst2_LFInst_14_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_2_U5  ( .A1(SubCellInput[56]), .A2(
        SubCellInput[57]), .ZN(SubCellInst2_LFInst_14_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_2_U4  ( .A1(
        SubCellInst2_LFInst_14_LFInst_2_n15 ), .A2(SubCellInput[59]), .ZN(
        SubCellInst2_LFInst_14_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst2_LFInst_14_LFInst_2_U3  ( .A(SubCellInput[56]), .B(
        SubCellInput[57]), .ZN(SubCellInst2_LFInst_14_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_3_U9  ( .A1(
        SubCellInst2_LFInst_14_LFInst_3_n16 ), .A2(
        SubCellInst2_LFInst_14_LFInst_3_n15 ), .ZN(MCInst2_MC1_v0_3 [0]) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_3_U8  ( .A1(SubCellInput[57]), .A2(
        SubCellInst2_LFInst_14_LFInst_3_n14 ), .ZN(
        SubCellInst2_LFInst_14_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst2_LFInst_14_LFInst_3_U7  ( .A(SubCellInput[59]), .B(
        SubCellInput[58]), .Z(SubCellInst2_LFInst_14_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_3_U6  ( .A1(
        SubCellInst2_LFInst_14_LFInst_3_n13 ), .A2(
        SubCellInst2_LFInst_14_LFInst_3_n12 ), .ZN(
        SubCellInst2_LFInst_14_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_14_LFInst_3_U5  ( .A1(SubCellInput[56]), .A2(
        SubCellInput[58]), .ZN(SubCellInst2_LFInst_14_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst2_LFInst_14_LFInst_3_U4  ( .A(SubCellInput[56]), .B(
        SubCellInst2_LFInst_14_LFInst_3_n11 ), .ZN(
        SubCellInst2_LFInst_14_LFInst_3_n13 ) );
  OR2_X1 SubCellInst2_LFInst_14_LFInst_3_U3  ( .A1(SubCellInput[59]), .A2(
        SubCellInput[57]), .ZN(SubCellInst2_LFInst_14_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_0_U6  ( .A1(SubCellInput[62]), .A2(
        SubCellInst2_LFInst_15_LFInst_0_n4 ), .ZN(
        SubCellInst2_LFInst_15_LFInst_0_n5 ) );
  INV_X1 SubCellInst2_LFInst_15_LFInst_0_U5  ( .A(SubCellInput[61]), .ZN(
        SubCellInst2_LFInst_15_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst2_LFInst_15_LFInst_0_U4  ( .A(SubCellInput[60]), .B(
        SubCellInput[63]), .Z(SubCellInst2_LFInst_15_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst2_LFInst_15_LFInst_0_U3  ( .A(
        SubCellInst2_LFInst_15_LFInst_0_n6 ), .B(
        SubCellInst2_LFInst_15_LFInst_0_n5 ), .ZN(Red_MCInst2_MC0_v0_1[0] )
         );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_1_U12  ( .A1(
        SubCellInst2_LFInst_15_LFInst_1_n18 ), .A2(
        SubCellInst2_LFInst_15_LFInst_1_n17 ), .ZN(MCInst2_MC0_v0_0 [3]) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_1_U11  ( .A1(SubCellInput[61]), .A2(
        SubCellInst2_LFInst_15_LFInst_1_n16 ), .ZN(
        SubCellInst2_LFInst_15_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst2_LFInst_15_LFInst_1_U10  ( .A1(SubCellInput[63]), .A2(
        SubCellInst2_LFInst_15_LFInst_1_n15 ), .ZN(
        SubCellInst2_LFInst_15_LFInst_1_n16 ) );
  AND2_X1 SubCellInst2_LFInst_15_LFInst_1_U9  ( .A1(SubCellInput[60]), .A2(
        SubCellInput[62]), .ZN(SubCellInst2_LFInst_15_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_1_U8  ( .A1(SubCellInput[63]), .A2(
        SubCellInst2_LFInst_15_LFInst_1_n14 ), .ZN(
        SubCellInst2_LFInst_15_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_1_U7  ( .A1(
        SubCellInst2_LFInst_15_LFInst_1_n13 ), .A2(
        SubCellInst2_LFInst_15_LFInst_1_n12 ), .ZN(
        SubCellInst2_LFInst_15_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_1_U6  ( .A1(SubCellInput[60]), .A2(
        SubCellInput[62]), .ZN(SubCellInst2_LFInst_15_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_1_U5  ( .A1(
        SubCellInst2_LFInst_15_LFInst_1_n11 ), .A2(
        SubCellInst2_LFInst_15_LFInst_1_n10 ), .ZN(
        SubCellInst2_LFInst_15_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_1_U4  ( .A1(SubCellInput[60]), .A2(
        SubCellInput[61]), .ZN(SubCellInst2_LFInst_15_LFInst_1_n10 ) );
  INV_X1 SubCellInst2_LFInst_15_LFInst_1_U3  ( .A(SubCellInput[62]), .ZN(
        SubCellInst2_LFInst_15_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_2_U11  ( .A1(
        SubCellInst2_LFInst_15_LFInst_2_n22 ), .A2(
        SubCellInst2_LFInst_15_LFInst_2_n21 ), .ZN(MCInst2_MC0_v0_3 [3]) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_2_U10  ( .A1(SubCellInput[62]), .A2(
        SubCellInst2_LFInst_15_LFInst_2_n20 ), .ZN(
        SubCellInst2_LFInst_15_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst2_LFInst_15_LFInst_2_U9  ( .A1(SubCellInput[61]), .A2(
        SubCellInst2_LFInst_15_LFInst_2_n19 ), .ZN(
        SubCellInst2_LFInst_15_LFInst_2_n20 ) );
  INV_X1 SubCellInst2_LFInst_15_LFInst_2_U8  ( .A(SubCellInput[63]), .ZN(
        SubCellInst2_LFInst_15_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_2_U7  ( .A1(
        SubCellInst2_LFInst_15_LFInst_2_n18 ), .A2(
        SubCellInst2_LFInst_15_LFInst_2_n17 ), .ZN(
        SubCellInst2_LFInst_15_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst2_LFInst_15_LFInst_2_U6  ( .A(
        SubCellInst2_LFInst_15_LFInst_2_n16 ), .B(SubCellInput[62]), .Z(
        SubCellInst2_LFInst_15_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_2_U5  ( .A1(SubCellInput[60]), .A2(
        SubCellInput[61]), .ZN(SubCellInst2_LFInst_15_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_2_U4  ( .A1(
        SubCellInst2_LFInst_15_LFInst_2_n15 ), .A2(SubCellInput[63]), .ZN(
        SubCellInst2_LFInst_15_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst2_LFInst_15_LFInst_2_U3  ( .A(SubCellInput[60]), .B(
        SubCellInput[61]), .ZN(SubCellInst2_LFInst_15_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_3_U9  ( .A1(
        SubCellInst2_LFInst_15_LFInst_3_n16 ), .A2(
        SubCellInst2_LFInst_15_LFInst_3_n15 ), .ZN(MCInst2_MC0_v0_3 [0]) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_3_U8  ( .A1(SubCellInput[61]), .A2(
        SubCellInst2_LFInst_15_LFInst_3_n14 ), .ZN(
        SubCellInst2_LFInst_15_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst2_LFInst_15_LFInst_3_U7  ( .A(SubCellInput[63]), .B(
        SubCellInput[62]), .Z(SubCellInst2_LFInst_15_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_3_U6  ( .A1(
        SubCellInst2_LFInst_15_LFInst_3_n13 ), .A2(
        SubCellInst2_LFInst_15_LFInst_3_n12 ), .ZN(
        SubCellInst2_LFInst_15_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst2_LFInst_15_LFInst_3_U5  ( .A1(SubCellInput[60]), .A2(
        SubCellInput[62]), .ZN(SubCellInst2_LFInst_15_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst2_LFInst_15_LFInst_3_U4  ( .A(SubCellInput[60]), .B(
        SubCellInst2_LFInst_15_LFInst_3_n11 ), .ZN(
        SubCellInst2_LFInst_15_LFInst_3_n13 ) );
  OR2_X1 SubCellInst2_LFInst_15_LFInst_3_U3  ( .A1(SubCellInput[63]), .A2(
        SubCellInput[61]), .ZN(SubCellInst2_LFInst_15_LFInst_3_n11 ) );
  XNOR2_X1 MCInst2_MC0_v0_2Inst_0_U4  ( .A(MCInst2_MC0_v0_2Inst_0_n2 ), .B(
        MCInst2_MC0_v0_0 [3]), .ZN(MCInst2_MC0_v0_2 [0]) );
  XNOR2_X1 MCInst2_MC0_v0_2Inst_0_U3  ( .A(MCInst2_MC0_v0_3 [0]), .B(
        Red_MCInst2_MC0_v0_1[0] ), .ZN(MCInst2_MC0_v0_2Inst_0_n2 ) );
  XOR2_X1 MCInst2_MC0_v1_1Inst_0_U3  ( .A(Red_MCInst2_MC0_v1_1[0] ), .B(
        MCInst2_MC0_v1_0 [3]), .Z(MCInst2_MC0_v1_1 [0]) );
  XNOR2_X1 MCInst2_MC0_v1_2Inst_0_U4  ( .A(MCInst2_MC0_v1_2Inst_0_n2 ), .B(
        Red_MCInst2_MC0_v1_1[0] ), .ZN(MCInst2_MC0_v1_2 [0]) );
  XNOR2_X1 MCInst2_MC0_v1_2Inst_0_U3  ( .A(MCInst2_MC0_v1_0 [3]), .B(
        MCInst2_MC0_v1_3 [2]), .ZN(MCInst2_MC0_v1_2Inst_0_n2 ) );
  XOR2_X1 MCInst2_MC0_v2_1Inst_0_U3  ( .A(MCInst2_MC0_v2_3 [1]), .B(
        MCInst2_MC0_v2_0 [3]), .Z(MCInst2_MC0_v2_1 [0]) );
  XOR2_X1 MCInst2_MC0_v2_2Inst_0_U3  ( .A(MCInst2_MC0_v2_0 [2]), .B(
        MCInst2_MC0_v2_0 [0]), .Z(MCInst2_MC0_v2_2 [0]) );
  XNOR2_X1 MCInst2_MC0_v2_3Inst_0_U5  ( .A(MCInst2_MC0_v2_3Inst_0_n4 ), .B(
        MCInst2_MC0_v2_3Inst_0_n3 ), .ZN(MCInst2_MC0_v2_3 [0]) );
  XNOR2_X1 MCInst2_MC0_v2_3Inst_0_U4  ( .A(MCInst2_MC0_v2_0 [2]), .B(
        MCInst2_MC0_v2_3 [1]), .ZN(MCInst2_MC0_v2_3Inst_0_n3 ) );
  XOR2_X1 MCInst2_MC0_v2_3Inst_0_U3  ( .A(MCInst2_MC0_v2_0 [3]), .B(
        MCInst2_MC0_v2_0 [0]), .Z(MCInst2_MC0_v2_3Inst_0_n4 ) );
  XOR2_X1 MCInst2_MC0_v3_1Inst_0_U3  ( .A(Red_MCInst2_MC0_v3_1[0] ), .B(
        MCInst2_MC0_v3_2 [2]), .Z(MCInst2_MC0_v3_1 [0]) );
  XOR2_X1 MCInst2_MC0_v3_2Inst_0_U3  ( .A(MCInst2_MC0_v3_2 [3]), .B(
        MCInst2_MC0_v3_0 [2]), .Z(MCInst2_MC0_v3_2 [0]) );
  XNOR2_X1 MCInst2_MC0_v3_3Inst_0_U4  ( .A(MCInst2_MC0_v3_3Inst_0_n2 ), .B(
        MCInst2_MC0_v3_0 [2]), .ZN(MCInst2_MC0_v3_3 [0]) );
  XNOR2_X1 MCInst2_MC0_v3_3Inst_0_U3  ( .A(MCInst2_MC0_v3_2 [2]), .B(
        MCInst2_MC0_v3_2 [3]), .ZN(MCInst2_MC0_v3_3Inst_0_n2 ) );
  XOR2_X1 MCInst2_MC0_v0_0Inst_1_U3  ( .A(MCInst2_MC0_v0_3 [3]), .B(
        MCInst2_MC0_v0_3 [0]), .Z(MCInst2_MC0_v0_0 [1]) );
  XOR2_X1 MCInst2_MC0_v0_1Inst_1_U3  ( .A(MCInst2_MC0_v0_0 [3]), .B(
        MCInst2_MC0_v0_3 [3]), .Z(MCInst2_MC0_v0_1 [1]) );
  XNOR2_X1 MCInst2_MC0_v0_2Inst_1_U4  ( .A(MCInst2_MC0_v0_2Inst_1_n2 ), .B(
        MCInst2_MC0_v0_3 [3]), .ZN(MCInst2_MC0_v0_2 [1]) );
  XNOR2_X1 MCInst2_MC0_v0_2Inst_1_U3  ( .A(MCInst2_MC0_v0_3 [0]), .B(
        Red_MCInst2_MC0_v0_1[0] ), .ZN(MCInst2_MC0_v0_2Inst_1_n2 ) );
  XOR2_X1 MCInst2_MC0_v0_3Inst_1_U3  ( .A(Red_MCInst2_MC0_v0_1[0] ), .B(
        MCInst2_MC0_v0_3 [0]), .Z(MCInst2_MC0_v0_3 [1]) );
  XOR2_X1 MCInst2_MC0_v1_1Inst_1_U3  ( .A(MCInst2_MC0_v1_0 [0]), .B(
        Red_MCInst2_MC0_v1_1[0] ), .Z(MCInst2_MC0_v1_1 [1]) );
  XOR2_X1 MCInst2_MC0_v1_2Inst_1_U3  ( .A(MCInst2_MC0_v1_0 [0]), .B(
        MCInst2_MC0_v1_3 [2]), .Z(MCInst2_MC0_v1_2 [1]) );
  XOR2_X1 MCInst2_MC0_v1_3Inst_1_U3  ( .A(MCInst2_MC0_v1_0 [0]), .B(
        MCInst2_MC0_v1_0 [3]), .Z(MCInst2_MC0_v1_3 [1]) );
  XOR2_X1 MCInst2_MC0_v2_0Inst_1_U3  ( .A(MCInst2_MC0_v2_3 [1]), .B(
        MCInst2_MC0_v2_0 [0]), .Z(MCInst2_MC0_v2_0 [1]) );
  XNOR2_X1 MCInst2_MC0_v2_1Inst_1_U4  ( .A(MCInst2_MC0_v2_1Inst_1_n2 ), .B(
        MCInst2_MC0_v2_0 [3]), .ZN(MCInst2_MC0_v2_1 [1]) );
  XNOR2_X1 MCInst2_MC0_v2_1Inst_1_U3  ( .A(MCInst2_MC0_v2_0 [0]), .B(
        MCInst2_MC0_v2_0 [2]), .ZN(MCInst2_MC0_v2_1Inst_1_n2 ) );
  XNOR2_X1 MCInst2_MC0_v2_2Inst_1_U5  ( .A(MCInst2_MC0_v2_2Inst_1_n4 ), .B(
        MCInst2_MC0_v2_2Inst_1_n3 ), .ZN(MCInst2_MC0_v2_2 [1]) );
  XNOR2_X1 MCInst2_MC0_v2_2Inst_1_U4  ( .A(MCInst2_MC0_v2_0 [2]), .B(
        MCInst2_MC0_v2_3 [1]), .ZN(MCInst2_MC0_v2_2Inst_1_n3 ) );
  XOR2_X1 MCInst2_MC0_v2_2Inst_1_U3  ( .A(MCInst2_MC0_v2_0 [3]), .B(
        MCInst2_MC0_v2_0 [0]), .Z(MCInst2_MC0_v2_2Inst_1_n4 ) );
  XOR2_X1 MCInst2_MC0_v3_0Inst_1_U3  ( .A(MCInst2_MC0_v3_2 [3]), .B(
        MCInst2_MC0_v3_2 [2]), .Z(MCInst2_MC0_v3_0 [1]) );
  XOR2_X1 MCInst2_MC0_v3_1Inst_1_U3  ( .A(MCInst2_MC0_v3_2 [3]), .B(
        Red_MCInst2_MC0_v3_1[0] ), .Z(MCInst2_MC0_v3_1 [1]) );
  XNOR2_X1 MCInst2_MC0_v3_3Inst_1_U4  ( .A(MCInst2_MC0_v3_3Inst_1_n2 ), .B(
        Red_MCInst2_MC0_v3_1[0] ), .ZN(MCInst2_MC0_v3_3 [1]) );
  XNOR2_X1 MCInst2_MC0_v3_3Inst_1_U3  ( .A(MCInst2_MC0_v3_2 [2]), .B(
        MCInst2_MC0_v3_2 [3]), .ZN(MCInst2_MC0_v3_3Inst_1_n2 ) );
  XOR2_X1 MCInst2_MC0_v0_0Inst_2_U3  ( .A(Red_MCInst2_MC0_v0_1[0] ), .B(
        MCInst2_MC0_v0_3 [0]), .Z(MCInst2_MC0_v0_0 [2]) );
  XOR2_X1 MCInst2_MC0_v0_1Inst_2_U3  ( .A(MCInst2_MC0_v0_3 [3]), .B(
        MCInst2_MC0_v0_3 [0]), .Z(MCInst2_MC0_v0_1 [2]) );
  XOR2_X1 MCInst2_MC0_v0_2Inst_2_U3  ( .A(MCInst2_MC0_v0_0 [3]), .B(
        MCInst2_MC0_v0_3 [0]), .Z(MCInst2_MC0_v0_2 [2]) );
  XNOR2_X1 MCInst2_MC0_v1_1Inst_2_U4  ( .A(MCInst2_MC0_v1_1Inst_2_n2 ), .B(
        MCInst2_MC0_v1_3 [2]), .ZN(MCInst2_MC0_v1_1 [2]) );
  XNOR2_X1 MCInst2_MC0_v1_1Inst_2_U3  ( .A(MCInst2_MC0_v1_0 [3]), .B(
        MCInst2_MC0_v1_0 [0]), .ZN(MCInst2_MC0_v1_1Inst_2_n2 ) );
  XNOR2_X1 MCInst2_MC0_v1_2Inst_2_U4  ( .A(MCInst2_MC0_v1_2Inst_2_n2 ), .B(
        MCInst2_MC0_v1_3 [2]), .ZN(MCInst2_MC0_v1_2 [2]) );
  XNOR2_X1 MCInst2_MC0_v1_2Inst_2_U3  ( .A(Red_MCInst2_MC0_v1_1[0] ), .B(
        MCInst2_MC0_v1_0 [0]), .ZN(MCInst2_MC0_v1_2Inst_2_n2 ) );
  XNOR2_X1 MCInst2_MC0_v2_1Inst_2_U4  ( .A(MCInst2_MC0_v2_1Inst_2_n2 ), .B(
        MCInst2_MC0_v2_0 [3]), .ZN(MCInst2_MC0_v2_1 [2]) );
  XNOR2_X1 MCInst2_MC0_v2_1Inst_2_U3  ( .A(MCInst2_MC0_v2_0 [0]), .B(
        MCInst2_MC0_v2_3 [1]), .ZN(MCInst2_MC0_v2_1Inst_2_n2 ) );
  XNOR2_X1 MCInst2_MC0_v2_2Inst_2_U4  ( .A(MCInst2_MC0_v2_2Inst_2_n2 ), .B(
        MCInst2_MC0_v2_0 [3]), .ZN(MCInst2_MC0_v2_2 [2]) );
  XNOR2_X1 MCInst2_MC0_v2_2Inst_2_U3  ( .A(MCInst2_MC0_v2_0 [0]), .B(
        MCInst2_MC0_v2_0 [2]), .ZN(MCInst2_MC0_v2_2Inst_2_n2 ) );
  XOR2_X1 MCInst2_MC0_v2_3Inst_2_U3  ( .A(MCInst2_MC0_v2_3 [1]), .B(
        MCInst2_MC0_v2_0 [2]), .Z(MCInst2_MC0_v2_3 [2]) );
  XNOR2_X1 MCInst2_MC0_v3_1Inst_2_U4  ( .A(MCInst2_MC0_v3_1Inst_2_n2 ), .B(
        MCInst2_MC0_v3_0 [2]), .ZN(MCInst2_MC0_v3_1 [2]) );
  XNOR2_X1 MCInst2_MC0_v3_1Inst_2_U3  ( .A(MCInst2_MC0_v3_2 [2]), .B(
        MCInst2_MC0_v3_2 [3]), .ZN(MCInst2_MC0_v3_1Inst_2_n2 ) );
  XOR2_X1 MCInst2_MC0_v3_3Inst_2_U3  ( .A(MCInst2_MC0_v3_0 [2]), .B(
        MCInst2_MC0_v3_2 [2]), .Z(MCInst2_MC0_v3_3 [2]) );
  XOR2_X1 MCInst2_MC0_v0_1Inst_3_U3  ( .A(Red_MCInst2_MC0_v0_1[0] ), .B(
        MCInst2_MC0_v0_3 [0]), .Z(MCInst2_MC0_v0_1 [3]) );
  XOR2_X1 MCInst2_MC0_v0_2Inst_3_U3  ( .A(Red_MCInst2_MC0_v0_1[0] ), .B(
        MCInst2_MC0_v0_3 [3]), .Z(MCInst2_MC0_v0_2 [3]) );
  XOR2_X1 MCInst2_MC0_v1_1Inst_3_U3  ( .A(MCInst2_MC0_v1_3 [2]), .B(
        Red_MCInst2_MC0_v1_1[0] ), .Z(MCInst2_MC0_v1_1 [3]) );
  XNOR2_X1 MCInst2_MC0_v1_2Inst_3_U5  ( .A(MCInst2_MC0_v1_2Inst_3_n4 ), .B(
        MCInst2_MC0_v1_2Inst_3_n3 ), .ZN(MCInst2_MC0_v1_2 [3]) );
  XNOR2_X1 MCInst2_MC0_v1_2Inst_3_U4  ( .A(MCInst2_MC0_v1_3 [2]), .B(
        MCInst2_MC0_v1_0 [0]), .ZN(MCInst2_MC0_v1_2Inst_3_n3 ) );
  XOR2_X1 MCInst2_MC0_v1_2Inst_3_U3  ( .A(Red_MCInst2_MC0_v1_1[0] ), .B(
        MCInst2_MC0_v1_0 [3]), .Z(MCInst2_MC0_v1_2Inst_3_n4 ) );
  XOR2_X1 MCInst2_MC0_v2_1Inst_3_U3  ( .A(MCInst2_MC0_v2_0 [2]), .B(
        MCInst2_MC0_v2_0 [0]), .Z(MCInst2_MC0_v2_1 [3]) );
  XNOR2_X1 MCInst2_MC0_v2_2Inst_3_U4  ( .A(MCInst2_MC0_v2_2Inst_3_n2 ), .B(
        MCInst2_MC0_v2_0 [3]), .ZN(MCInst2_MC0_v2_2 [3]) );
  XNOR2_X1 MCInst2_MC0_v2_2Inst_3_U3  ( .A(MCInst2_MC0_v2_0 [0]), .B(
        MCInst2_MC0_v2_3 [1]), .ZN(MCInst2_MC0_v2_2Inst_3_n2 ) );
  XNOR2_X1 MCInst2_MC0_v2_3Inst_3_U4  ( .A(MCInst2_MC0_v2_3Inst_3_n2 ), .B(
        MCInst2_MC0_v2_0 [2]), .ZN(MCInst2_MC0_v2_3 [3]) );
  XNOR2_X1 MCInst2_MC0_v2_3Inst_3_U3  ( .A(MCInst2_MC0_v2_0 [3]), .B(
        MCInst2_MC0_v2_3 [1]), .ZN(MCInst2_MC0_v2_3Inst_3_n2 ) );
  XOR2_X1 MCInst2_MC0_v3_1Inst_3_U3  ( .A(MCInst2_MC0_v3_0 [2]), .B(
        Red_MCInst2_MC0_v3_1[0] ), .Z(MCInst2_MC0_v3_1 [3]) );
  XOR2_X1 MCInst2_MC0_v3_3Inst_3_U3  ( .A(MCInst2_MC0_v3_2 [3]), .B(
        Red_MCInst2_MC0_v3_1[0] ), .Z(MCInst2_MC0_v3_3 [3]) );
  XNOR2_X1 MCInst2_MC0_r0Inst_XORInst_0_0_U3  ( .A(
        MCInst2_MC0_r0Inst_XORInst_0_0_n5 ), .B(
        MCInst2_MC0_r0Inst_XORInst_0_0_n4 ), .ZN(Feedback2[60]) );
  XNOR2_X1 MCInst2_MC0_r0Inst_XORInst_0_0_U2  ( .A(MCInst2_MC0_v3_2 [2]), 
        .B(MCInst2_MC0_v2_0 [0]), .ZN(MCInst2_MC0_r0Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst2_MC0_r0Inst_XORInst_0_0_U1  ( .A(MCInst2_MC0_v0_3 [3]), .B(
        MCInst2_MC0_v1_0 [0]), .Z(MCInst2_MC0_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst2_MC0_r0Inst_XORInst_0_1_U3  ( .A(
        MCInst2_MC0_r0Inst_XORInst_0_1_n5 ), .B(
        MCInst2_MC0_r0Inst_XORInst_0_1_n4 ), .ZN(Feedback2[61]) );
  XNOR2_X1 MCInst2_MC0_r0Inst_XORInst_0_1_U2  ( .A(MCInst2_MC0_v3_0 [1]), 
        .B(MCInst2_MC0_v2_0 [1]), .ZN(MCInst2_MC0_r0Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst2_MC0_r0Inst_XORInst_0_1_U1  ( .A(MCInst2_MC0_v0_0 [1]), .B(
        MCInst2_MC0_v1_3 [2]), .Z(MCInst2_MC0_r0Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst2_MC0_r0Inst_XORInst_0_2_U3  ( .A(
        MCInst2_MC0_r0Inst_XORInst_0_2_n5 ), .B(
        MCInst2_MC0_r0Inst_XORInst_0_2_n4 ), .ZN(Feedback2[62]) );
  XNOR2_X1 MCInst2_MC0_r0Inst_XORInst_0_2_U2  ( .A(MCInst2_MC0_v3_0 [2]), 
        .B(MCInst2_MC0_v2_0 [2]), .ZN(MCInst2_MC0_r0Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst2_MC0_r0Inst_XORInst_0_2_U1  ( .A(MCInst2_MC0_v0_0 [2]), .B(
        Red_MCInst2_MC0_v1_1[0] ), .Z(MCInst2_MC0_r0Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst2_MC0_r0Inst_XORInst_0_3_U3  ( .A(
        MCInst2_MC0_r0Inst_XORInst_0_3_n5 ), .B(
        MCInst2_MC0_r0Inst_XORInst_0_3_n4 ), .ZN(Feedback2[63]) );
  XNOR2_X1 MCInst2_MC0_r0Inst_XORInst_0_3_U2  ( .A(Red_MCInst2_MC0_v3_1[0] ), 
        .B(MCInst2_MC0_v2_0 [3]), .ZN(MCInst2_MC0_r0Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst2_MC0_r0Inst_XORInst_0_3_U1  ( .A(MCInst2_MC0_v0_0 [3]), .B(
        MCInst2_MC0_v1_0 [3]), .Z(MCInst2_MC0_r0Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst2_MC0_r1Inst_XORInst_0_0_U3  ( .A(
        MCInst2_MC0_r1Inst_XORInst_0_0_n5 ), .B(
        MCInst2_MC0_r1Inst_XORInst_0_0_n4 ), .ZN(Feedback2[44]) );
  XNOR2_X1 MCInst2_MC0_r1Inst_XORInst_0_0_U2  ( .A(MCInst2_MC0_v3_1 [0]), 
        .B(MCInst2_MC0_v2_1 [0]), .ZN(MCInst2_MC0_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst2_MC0_r1Inst_XORInst_0_0_U1  ( .A(MCInst2_MC0_v0_0 [3]), .B(
        MCInst2_MC0_v1_1 [0]), .Z(MCInst2_MC0_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst2_MC0_r1Inst_XORInst_0_1_U3  ( .A(
        MCInst2_MC0_r1Inst_XORInst_0_1_n5 ), .B(
        MCInst2_MC0_r1Inst_XORInst_0_1_n4 ), .ZN(Feedback2[45]) );
  XNOR2_X1 MCInst2_MC0_r1Inst_XORInst_0_1_U2  ( .A(MCInst2_MC0_v3_1 [1]), 
        .B(MCInst2_MC0_v2_1 [1]), .ZN(MCInst2_MC0_r1Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst2_MC0_r1Inst_XORInst_0_1_U1  ( .A(MCInst2_MC0_v0_1 [1]), .B(
        MCInst2_MC0_v1_1 [1]), .Z(MCInst2_MC0_r1Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst2_MC0_r1Inst_XORInst_0_2_U3  ( .A(
        MCInst2_MC0_r1Inst_XORInst_0_2_n5 ), .B(
        MCInst2_MC0_r1Inst_XORInst_0_2_n4 ), .ZN(Feedback2[46]) );
  XNOR2_X1 MCInst2_MC0_r1Inst_XORInst_0_2_U2  ( .A(MCInst2_MC0_v3_1 [2]), 
        .B(MCInst2_MC0_v2_1 [2]), .ZN(MCInst2_MC0_r1Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst2_MC0_r1Inst_XORInst_0_2_U1  ( .A(MCInst2_MC0_v0_1 [2]), .B(
        MCInst2_MC0_v1_1 [2]), .Z(MCInst2_MC0_r1Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst2_MC0_r1Inst_XORInst_0_3_U3  ( .A(
        MCInst2_MC0_r1Inst_XORInst_0_3_n5 ), .B(
        MCInst2_MC0_r1Inst_XORInst_0_3_n4 ), .ZN(Feedback2[47]) );
  XNOR2_X1 MCInst2_MC0_r1Inst_XORInst_0_3_U2  ( .A(MCInst2_MC0_v3_1 [3]), 
        .B(MCInst2_MC0_v2_1 [3]), .ZN(MCInst2_MC0_r1Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst2_MC0_r1Inst_XORInst_0_3_U1  ( .A(MCInst2_MC0_v0_1 [3]), .B(
        MCInst2_MC0_v1_1 [3]), .Z(MCInst2_MC0_r1Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst2_MC0_r2Inst_XORInst_0_0_U3  ( .A(
        MCInst2_MC0_r2Inst_XORInst_0_0_n5 ), .B(
        MCInst2_MC0_r2Inst_XORInst_0_0_n4 ), .ZN(Feedback2[28]) );
  XNOR2_X1 MCInst2_MC0_r2Inst_XORInst_0_0_U2  ( .A(MCInst2_MC0_v3_2 [0]), 
        .B(MCInst2_MC0_v2_2 [0]), .ZN(MCInst2_MC0_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst2_MC0_r2Inst_XORInst_0_0_U1  ( .A(MCInst2_MC0_v0_2 [0]), .B(
        MCInst2_MC0_v1_2 [0]), .Z(MCInst2_MC0_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst2_MC0_r2Inst_XORInst_0_1_U3  ( .A(
        MCInst2_MC0_r2Inst_XORInst_0_1_n5 ), .B(
        MCInst2_MC0_r2Inst_XORInst_0_1_n4 ), .ZN(Feedback2[29]) );
  XNOR2_X1 MCInst2_MC0_r2Inst_XORInst_0_1_U2  ( .A(Red_MCInst2_MC0_v3_1[0] ), 
        .B(MCInst2_MC0_v2_2 [1]), .ZN(MCInst2_MC0_r2Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst2_MC0_r2Inst_XORInst_0_1_U1  ( .A(MCInst2_MC0_v0_2 [1]), .B(
        MCInst2_MC0_v1_2 [1]), .Z(MCInst2_MC0_r2Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst2_MC0_r2Inst_XORInst_0_2_U3  ( .A(
        MCInst2_MC0_r2Inst_XORInst_0_2_n5 ), .B(
        MCInst2_MC0_r2Inst_XORInst_0_2_n4 ), .ZN(Feedback2[30]) );
  XNOR2_X1 MCInst2_MC0_r2Inst_XORInst_0_2_U2  ( .A(MCInst2_MC0_v3_2 [2]), 
        .B(MCInst2_MC0_v2_2 [2]), .ZN(MCInst2_MC0_r2Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst2_MC0_r2Inst_XORInst_0_2_U1  ( .A(MCInst2_MC0_v0_2 [2]), .B(
        MCInst2_MC0_v1_2 [2]), .Z(MCInst2_MC0_r2Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst2_MC0_r2Inst_XORInst_0_3_U3  ( .A(
        MCInst2_MC0_r2Inst_XORInst_0_3_n5 ), .B(
        MCInst2_MC0_r2Inst_XORInst_0_3_n4 ), .ZN(Feedback2[31]) );
  XNOR2_X1 MCInst2_MC0_r2Inst_XORInst_0_3_U2  ( .A(MCInst2_MC0_v3_2 [3]), 
        .B(MCInst2_MC0_v2_2 [3]), .ZN(MCInst2_MC0_r2Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst2_MC0_r2Inst_XORInst_0_3_U1  ( .A(MCInst2_MC0_v0_2 [3]), .B(
        MCInst2_MC0_v1_2 [3]), .Z(MCInst2_MC0_r2Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst2_MC0_r3Inst_XORInst_0_0_U3  ( .A(
        MCInst2_MC0_r3Inst_XORInst_0_0_n5 ), .B(
        MCInst2_MC0_r3Inst_XORInst_0_0_n4 ), .ZN(Feedback2[12]) );
  XNOR2_X1 MCInst2_MC0_r3Inst_XORInst_0_0_U2  ( .A(MCInst2_MC0_v3_3 [0]), 
        .B(MCInst2_MC0_v2_3 [0]), .ZN(MCInst2_MC0_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst2_MC0_r3Inst_XORInst_0_0_U1  ( .A(MCInst2_MC0_v0_3 [0]), .B(
        MCInst2_MC0_v1_0 [3]), .Z(MCInst2_MC0_r3Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst2_MC0_r3Inst_XORInst_0_1_U3  ( .A(
        MCInst2_MC0_r3Inst_XORInst_0_1_n5 ), .B(
        MCInst2_MC0_r3Inst_XORInst_0_1_n4 ), .ZN(Feedback2[13]) );
  XNOR2_X1 MCInst2_MC0_r3Inst_XORInst_0_1_U2  ( .A(MCInst2_MC0_v3_3 [1]), 
        .B(MCInst2_MC0_v2_3 [1]), .ZN(MCInst2_MC0_r3Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst2_MC0_r3Inst_XORInst_0_1_U1  ( .A(MCInst2_MC0_v0_3 [1]), .B(
        MCInst2_MC0_v1_3 [1]), .Z(MCInst2_MC0_r3Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst2_MC0_r3Inst_XORInst_0_2_U3  ( .A(
        MCInst2_MC0_r3Inst_XORInst_0_2_n5 ), .B(
        MCInst2_MC0_r3Inst_XORInst_0_2_n4 ), .ZN(Feedback2[14]) );
  XNOR2_X1 MCInst2_MC0_r3Inst_XORInst_0_2_U2  ( .A(MCInst2_MC0_v3_3 [2]), 
        .B(MCInst2_MC0_v2_3 [2]), .ZN(MCInst2_MC0_r3Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst2_MC0_r3Inst_XORInst_0_2_U1  ( .A(MCInst2_MC0_v0_0 [3]), .B(
        MCInst2_MC0_v1_3 [2]), .Z(MCInst2_MC0_r3Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst2_MC0_r3Inst_XORInst_0_3_U3  ( .A(
        MCInst2_MC0_r3Inst_XORInst_0_3_n5 ), .B(
        MCInst2_MC0_r3Inst_XORInst_0_3_n4 ), .ZN(Feedback2[15]) );
  XNOR2_X1 MCInst2_MC0_r3Inst_XORInst_0_3_U2  ( .A(MCInst2_MC0_v3_3 [3]), 
        .B(MCInst2_MC0_v2_3 [3]), .ZN(MCInst2_MC0_r3Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst2_MC0_r3Inst_XORInst_0_3_U1  ( .A(MCInst2_MC0_v0_3 [3]), .B(
        Red_MCInst2_MC0_v1_1[0] ), .Z(MCInst2_MC0_r3Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst2_MC1_v0_2Inst_0_U4  ( .A(MCInst2_MC1_v0_2Inst_0_n2 ), .B(
        MCInst2_MC1_v0_0 [3]), .ZN(MCInst2_MC1_v0_2 [0]) );
  XNOR2_X1 MCInst2_MC1_v0_2Inst_0_U3  ( .A(MCInst2_MC1_v0_3 [0]), .B(
        Red_MCInst2_MC1_v0_1[0] ), .ZN(MCInst2_MC1_v0_2Inst_0_n2 ) );
  XOR2_X1 MCInst2_MC1_v1_1Inst_0_U3  ( .A(Red_MCInst2_MC1_v1_1[0] ), .B(
        MCInst2_MC1_v1_0 [3]), .Z(MCInst2_MC1_v1_1 [0]) );
  XNOR2_X1 MCInst2_MC1_v1_2Inst_0_U4  ( .A(MCInst2_MC1_v1_2Inst_0_n2 ), .B(
        Red_MCInst2_MC1_v1_1[0] ), .ZN(MCInst2_MC1_v1_2 [0]) );
  XNOR2_X1 MCInst2_MC1_v1_2Inst_0_U3  ( .A(MCInst2_MC1_v1_0 [3]), .B(
        MCInst2_MC1_v1_3 [2]), .ZN(MCInst2_MC1_v1_2Inst_0_n2 ) );
  XOR2_X1 MCInst2_MC1_v2_1Inst_0_U3  ( .A(MCInst2_MC1_v2_3 [1]), .B(
        MCInst2_MC1_v2_0 [3]), .Z(MCInst2_MC1_v2_1 [0]) );
  XOR2_X1 MCInst2_MC1_v2_2Inst_0_U3  ( .A(MCInst2_MC1_v2_0 [2]), .B(
        MCInst2_MC1_v2_0 [0]), .Z(MCInst2_MC1_v2_2 [0]) );
  XNOR2_X1 MCInst2_MC1_v2_3Inst_0_U5  ( .A(MCInst2_MC1_v2_3Inst_0_n4 ), .B(
        MCInst2_MC1_v2_3Inst_0_n3 ), .ZN(MCInst2_MC1_v2_3 [0]) );
  XNOR2_X1 MCInst2_MC1_v2_3Inst_0_U4  ( .A(MCInst2_MC1_v2_0 [2]), .B(
        MCInst2_MC1_v2_3 [1]), .ZN(MCInst2_MC1_v2_3Inst_0_n3 ) );
  XOR2_X1 MCInst2_MC1_v2_3Inst_0_U3  ( .A(MCInst2_MC1_v2_0 [3]), .B(
        MCInst2_MC1_v2_0 [0]), .Z(MCInst2_MC1_v2_3Inst_0_n4 ) );
  XOR2_X1 MCInst2_MC1_v3_1Inst_0_U3  ( .A(Red_MCInst2_MC1_v3_1[0] ), .B(
        MCInst2_MC1_v3_2 [2]), .Z(MCInst2_MC1_v3_1 [0]) );
  XOR2_X1 MCInst2_MC1_v3_2Inst_0_U3  ( .A(MCInst2_MC1_v3_2 [3]), .B(
        MCInst2_MC1_v3_0 [2]), .Z(MCInst2_MC1_v3_2 [0]) );
  XNOR2_X1 MCInst2_MC1_v3_3Inst_0_U4  ( .A(MCInst2_MC1_v3_3Inst_0_n2 ), .B(
        MCInst2_MC1_v3_0 [2]), .ZN(MCInst2_MC1_v3_3 [0]) );
  XNOR2_X1 MCInst2_MC1_v3_3Inst_0_U3  ( .A(MCInst2_MC1_v3_2 [2]), .B(
        MCInst2_MC1_v3_2 [3]), .ZN(MCInst2_MC1_v3_3Inst_0_n2 ) );
  XOR2_X1 MCInst2_MC1_v0_0Inst_1_U3  ( .A(MCInst2_MC1_v0_3 [3]), .B(
        MCInst2_MC1_v0_3 [0]), .Z(MCInst2_MC1_v0_0 [1]) );
  XOR2_X1 MCInst2_MC1_v0_1Inst_1_U3  ( .A(MCInst2_MC1_v0_0 [3]), .B(
        MCInst2_MC1_v0_3 [3]), .Z(MCInst2_MC1_v0_1 [1]) );
  XNOR2_X1 MCInst2_MC1_v0_2Inst_1_U4  ( .A(MCInst2_MC1_v0_2Inst_1_n2 ), .B(
        MCInst2_MC1_v0_3 [3]), .ZN(MCInst2_MC1_v0_2 [1]) );
  XNOR2_X1 MCInst2_MC1_v0_2Inst_1_U3  ( .A(MCInst2_MC1_v0_3 [0]), .B(
        Red_MCInst2_MC1_v0_1[0] ), .ZN(MCInst2_MC1_v0_2Inst_1_n2 ) );
  XOR2_X1 MCInst2_MC1_v0_3Inst_1_U3  ( .A(Red_MCInst2_MC1_v0_1[0] ), .B(
        MCInst2_MC1_v0_3 [0]), .Z(MCInst2_MC1_v0_3 [1]) );
  XOR2_X1 MCInst2_MC1_v1_1Inst_1_U3  ( .A(MCInst2_MC1_v1_0 [0]), .B(
        Red_MCInst2_MC1_v1_1[0] ), .Z(MCInst2_MC1_v1_1 [1]) );
  XOR2_X1 MCInst2_MC1_v1_2Inst_1_U3  ( .A(MCInst2_MC1_v1_0 [0]), .B(
        MCInst2_MC1_v1_3 [2]), .Z(MCInst2_MC1_v1_2 [1]) );
  XOR2_X1 MCInst2_MC1_v1_3Inst_1_U3  ( .A(MCInst2_MC1_v1_0 [0]), .B(
        MCInst2_MC1_v1_0 [3]), .Z(MCInst2_MC1_v1_3 [1]) );
  XOR2_X1 MCInst2_MC1_v2_0Inst_1_U3  ( .A(MCInst2_MC1_v2_3 [1]), .B(
        MCInst2_MC1_v2_0 [0]), .Z(MCInst2_MC1_v2_0 [1]) );
  XNOR2_X1 MCInst2_MC1_v2_1Inst_1_U4  ( .A(MCInst2_MC1_v2_1Inst_1_n2 ), .B(
        MCInst2_MC1_v2_0 [3]), .ZN(MCInst2_MC1_v2_1 [1]) );
  XNOR2_X1 MCInst2_MC1_v2_1Inst_1_U3  ( .A(MCInst2_MC1_v2_0 [0]), .B(
        MCInst2_MC1_v2_0 [2]), .ZN(MCInst2_MC1_v2_1Inst_1_n2 ) );
  XNOR2_X1 MCInst2_MC1_v2_2Inst_1_U5  ( .A(MCInst2_MC1_v2_2Inst_1_n4 ), .B(
        MCInst2_MC1_v2_2Inst_1_n3 ), .ZN(MCInst2_MC1_v2_2 [1]) );
  XNOR2_X1 MCInst2_MC1_v2_2Inst_1_U4  ( .A(MCInst2_MC1_v2_0 [2]), .B(
        MCInst2_MC1_v2_3 [1]), .ZN(MCInst2_MC1_v2_2Inst_1_n3 ) );
  XOR2_X1 MCInst2_MC1_v2_2Inst_1_U3  ( .A(MCInst2_MC1_v2_0 [3]), .B(
        MCInst2_MC1_v2_0 [0]), .Z(MCInst2_MC1_v2_2Inst_1_n4 ) );
  XOR2_X1 MCInst2_MC1_v3_0Inst_1_U3  ( .A(MCInst2_MC1_v3_2 [3]), .B(
        MCInst2_MC1_v3_2 [2]), .Z(MCInst2_MC1_v3_0 [1]) );
  XOR2_X1 MCInst2_MC1_v3_1Inst_1_U3  ( .A(MCInst2_MC1_v3_2 [3]), .B(
        Red_MCInst2_MC1_v3_1[0] ), .Z(MCInst2_MC1_v3_1 [1]) );
  XNOR2_X1 MCInst2_MC1_v3_3Inst_1_U4  ( .A(MCInst2_MC1_v3_3Inst_1_n2 ), .B(
        Red_MCInst2_MC1_v3_1[0] ), .ZN(MCInst2_MC1_v3_3 [1]) );
  XNOR2_X1 MCInst2_MC1_v3_3Inst_1_U3  ( .A(MCInst2_MC1_v3_2 [2]), .B(
        MCInst2_MC1_v3_2 [3]), .ZN(MCInst2_MC1_v3_3Inst_1_n2 ) );
  XOR2_X1 MCInst2_MC1_v0_0Inst_2_U3  ( .A(Red_MCInst2_MC1_v0_1[0] ), .B(
        MCInst2_MC1_v0_3 [0]), .Z(MCInst2_MC1_v0_0 [2]) );
  XOR2_X1 MCInst2_MC1_v0_1Inst_2_U3  ( .A(MCInst2_MC1_v0_3 [3]), .B(
        MCInst2_MC1_v0_3 [0]), .Z(MCInst2_MC1_v0_1 [2]) );
  XOR2_X1 MCInst2_MC1_v0_2Inst_2_U3  ( .A(MCInst2_MC1_v0_0 [3]), .B(
        MCInst2_MC1_v0_3 [0]), .Z(MCInst2_MC1_v0_2 [2]) );
  XNOR2_X1 MCInst2_MC1_v1_1Inst_2_U4  ( .A(MCInst2_MC1_v1_1Inst_2_n2 ), .B(
        MCInst2_MC1_v1_3 [2]), .ZN(MCInst2_MC1_v1_1 [2]) );
  XNOR2_X1 MCInst2_MC1_v1_1Inst_2_U3  ( .A(MCInst2_MC1_v1_0 [3]), .B(
        MCInst2_MC1_v1_0 [0]), .ZN(MCInst2_MC1_v1_1Inst_2_n2 ) );
  XNOR2_X1 MCInst2_MC1_v1_2Inst_2_U4  ( .A(MCInst2_MC1_v1_2Inst_2_n2 ), .B(
        MCInst2_MC1_v1_3 [2]), .ZN(MCInst2_MC1_v1_2 [2]) );
  XNOR2_X1 MCInst2_MC1_v1_2Inst_2_U3  ( .A(Red_MCInst2_MC1_v1_1[0] ), .B(
        MCInst2_MC1_v1_0 [0]), .ZN(MCInst2_MC1_v1_2Inst_2_n2 ) );
  XNOR2_X1 MCInst2_MC1_v2_1Inst_2_U4  ( .A(MCInst2_MC1_v2_1Inst_2_n2 ), .B(
        MCInst2_MC1_v2_0 [3]), .ZN(MCInst2_MC1_v2_1 [2]) );
  XNOR2_X1 MCInst2_MC1_v2_1Inst_2_U3  ( .A(MCInst2_MC1_v2_0 [0]), .B(
        MCInst2_MC1_v2_3 [1]), .ZN(MCInst2_MC1_v2_1Inst_2_n2 ) );
  XNOR2_X1 MCInst2_MC1_v2_2Inst_2_U4  ( .A(MCInst2_MC1_v2_2Inst_2_n2 ), .B(
        MCInst2_MC1_v2_0 [3]), .ZN(MCInst2_MC1_v2_2 [2]) );
  XNOR2_X1 MCInst2_MC1_v2_2Inst_2_U3  ( .A(MCInst2_MC1_v2_0 [0]), .B(
        MCInst2_MC1_v2_0 [2]), .ZN(MCInst2_MC1_v2_2Inst_2_n2 ) );
  XOR2_X1 MCInst2_MC1_v2_3Inst_2_U3  ( .A(MCInst2_MC1_v2_3 [1]), .B(
        MCInst2_MC1_v2_0 [2]), .Z(MCInst2_MC1_v2_3 [2]) );
  XNOR2_X1 MCInst2_MC1_v3_1Inst_2_U4  ( .A(MCInst2_MC1_v3_1Inst_2_n2 ), .B(
        MCInst2_MC1_v3_0 [2]), .ZN(MCInst2_MC1_v3_1 [2]) );
  XNOR2_X1 MCInst2_MC1_v3_1Inst_2_U3  ( .A(MCInst2_MC1_v3_2 [2]), .B(
        MCInst2_MC1_v3_2 [3]), .ZN(MCInst2_MC1_v3_1Inst_2_n2 ) );
  XOR2_X1 MCInst2_MC1_v3_3Inst_2_U3  ( .A(MCInst2_MC1_v3_0 [2]), .B(
        MCInst2_MC1_v3_2 [2]), .Z(MCInst2_MC1_v3_3 [2]) );
  XOR2_X1 MCInst2_MC1_v0_1Inst_3_U3  ( .A(Red_MCInst2_MC1_v0_1[0] ), .B(
        MCInst2_MC1_v0_3 [0]), .Z(MCInst2_MC1_v0_1 [3]) );
  XOR2_X1 MCInst2_MC1_v0_2Inst_3_U3  ( .A(Red_MCInst2_MC1_v0_1[0] ), .B(
        MCInst2_MC1_v0_3 [3]), .Z(MCInst2_MC1_v0_2 [3]) );
  XOR2_X1 MCInst2_MC1_v1_1Inst_3_U3  ( .A(MCInst2_MC1_v1_3 [2]), .B(
        Red_MCInst2_MC1_v1_1[0] ), .Z(MCInst2_MC1_v1_1 [3]) );
  XNOR2_X1 MCInst2_MC1_v1_2Inst_3_U5  ( .A(MCInst2_MC1_v1_2Inst_3_n4 ), .B(
        MCInst2_MC1_v1_2Inst_3_n3 ), .ZN(MCInst2_MC1_v1_2 [3]) );
  XNOR2_X1 MCInst2_MC1_v1_2Inst_3_U4  ( .A(MCInst2_MC1_v1_3 [2]), .B(
        MCInst2_MC1_v1_0 [0]), .ZN(MCInst2_MC1_v1_2Inst_3_n3 ) );
  XOR2_X1 MCInst2_MC1_v1_2Inst_3_U3  ( .A(Red_MCInst2_MC1_v1_1[0] ), .B(
        MCInst2_MC1_v1_0 [3]), .Z(MCInst2_MC1_v1_2Inst_3_n4 ) );
  XOR2_X1 MCInst2_MC1_v2_1Inst_3_U3  ( .A(MCInst2_MC1_v2_0 [2]), .B(
        MCInst2_MC1_v2_0 [0]), .Z(MCInst2_MC1_v2_1 [3]) );
  XNOR2_X1 MCInst2_MC1_v2_2Inst_3_U4  ( .A(MCInst2_MC1_v2_2Inst_3_n2 ), .B(
        MCInst2_MC1_v2_0 [3]), .ZN(MCInst2_MC1_v2_2 [3]) );
  XNOR2_X1 MCInst2_MC1_v2_2Inst_3_U3  ( .A(MCInst2_MC1_v2_0 [0]), .B(
        MCInst2_MC1_v2_3 [1]), .ZN(MCInst2_MC1_v2_2Inst_3_n2 ) );
  XNOR2_X1 MCInst2_MC1_v2_3Inst_3_U4  ( .A(MCInst2_MC1_v2_3Inst_3_n2 ), .B(
        MCInst2_MC1_v2_0 [2]), .ZN(MCInst2_MC1_v2_3 [3]) );
  XNOR2_X1 MCInst2_MC1_v2_3Inst_3_U3  ( .A(MCInst2_MC1_v2_0 [3]), .B(
        MCInst2_MC1_v2_3 [1]), .ZN(MCInst2_MC1_v2_3Inst_3_n2 ) );
  XOR2_X1 MCInst2_MC1_v3_1Inst_3_U3  ( .A(MCInst2_MC1_v3_0 [2]), .B(
        Red_MCInst2_MC1_v3_1[0] ), .Z(MCInst2_MC1_v3_1 [3]) );
  XOR2_X1 MCInst2_MC1_v3_3Inst_3_U3  ( .A(MCInst2_MC1_v3_2 [3]), .B(
        Red_MCInst2_MC1_v3_1[0] ), .Z(MCInst2_MC1_v3_3 [3]) );
  XNOR2_X1 MCInst2_MC1_r0Inst_XORInst_0_0_U3  ( .A(
        MCInst2_MC1_r0Inst_XORInst_0_0_n5 ), .B(
        MCInst2_MC1_r0Inst_XORInst_0_0_n4 ), .ZN(Feedback2[56]) );
  XNOR2_X1 MCInst2_MC1_r0Inst_XORInst_0_0_U2  ( .A(MCInst2_MC1_v3_2 [2]), 
        .B(MCInst2_MC1_v2_0 [0]), .ZN(MCInst2_MC1_r0Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst2_MC1_r0Inst_XORInst_0_0_U1  ( .A(MCInst2_MC1_v0_3 [3]), .B(
        MCInst2_MC1_v1_0 [0]), .Z(MCInst2_MC1_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst2_MC1_r0Inst_XORInst_0_1_U3  ( .A(
        MCInst2_MC1_r0Inst_XORInst_0_1_n5 ), .B(
        MCInst2_MC1_r0Inst_XORInst_0_1_n4 ), .ZN(Feedback2[57]) );
  XNOR2_X1 MCInst2_MC1_r0Inst_XORInst_0_1_U2  ( .A(MCInst2_MC1_v3_0 [1]), 
        .B(MCInst2_MC1_v2_0 [1]), .ZN(MCInst2_MC1_r0Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst2_MC1_r0Inst_XORInst_0_1_U1  ( .A(MCInst2_MC1_v0_0 [1]), .B(
        MCInst2_MC1_v1_3 [2]), .Z(MCInst2_MC1_r0Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst2_MC1_r0Inst_XORInst_0_2_U3  ( .A(
        MCInst2_MC1_r0Inst_XORInst_0_2_n5 ), .B(
        MCInst2_MC1_r0Inst_XORInst_0_2_n4 ), .ZN(Feedback2[58]) );
  XNOR2_X1 MCInst2_MC1_r0Inst_XORInst_0_2_U2  ( .A(MCInst2_MC1_v3_0 [2]), 
        .B(MCInst2_MC1_v2_0 [2]), .ZN(MCInst2_MC1_r0Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst2_MC1_r0Inst_XORInst_0_2_U1  ( .A(MCInst2_MC1_v0_0 [2]), .B(
        Red_MCInst2_MC1_v1_1[0] ), .Z(MCInst2_MC1_r0Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst2_MC1_r0Inst_XORInst_0_3_U3  ( .A(
        MCInst2_MC1_r0Inst_XORInst_0_3_n5 ), .B(
        MCInst2_MC1_r0Inst_XORInst_0_3_n4 ), .ZN(Feedback2[59]) );
  XNOR2_X1 MCInst2_MC1_r0Inst_XORInst_0_3_U2  ( .A(Red_MCInst2_MC1_v3_1[0] ), 
        .B(MCInst2_MC1_v2_0 [3]), .ZN(MCInst2_MC1_r0Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst2_MC1_r0Inst_XORInst_0_3_U1  ( .A(MCInst2_MC1_v0_0 [3]), .B(
        MCInst2_MC1_v1_0 [3]), .Z(MCInst2_MC1_r0Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst2_MC1_r1Inst_XORInst_0_0_U3  ( .A(
        MCInst2_MC1_r1Inst_XORInst_0_0_n5 ), .B(
        MCInst2_MC1_r1Inst_XORInst_0_0_n4 ), .ZN(Feedback2[40]) );
  XNOR2_X1 MCInst2_MC1_r1Inst_XORInst_0_0_U2  ( .A(MCInst2_MC1_v3_1 [0]), 
        .B(MCInst2_MC1_v2_1 [0]), .ZN(MCInst2_MC1_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst2_MC1_r1Inst_XORInst_0_0_U1  ( .A(MCInst2_MC1_v0_0 [3]), .B(
        MCInst2_MC1_v1_1 [0]), .Z(MCInst2_MC1_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst2_MC1_r1Inst_XORInst_0_1_U3  ( .A(
        MCInst2_MC1_r1Inst_XORInst_0_1_n5 ), .B(
        MCInst2_MC1_r1Inst_XORInst_0_1_n4 ), .ZN(Feedback2[41]) );
  XNOR2_X1 MCInst2_MC1_r1Inst_XORInst_0_1_U2  ( .A(MCInst2_MC1_v3_1 [1]), 
        .B(MCInst2_MC1_v2_1 [1]), .ZN(MCInst2_MC1_r1Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst2_MC1_r1Inst_XORInst_0_1_U1  ( .A(MCInst2_MC1_v0_1 [1]), .B(
        MCInst2_MC1_v1_1 [1]), .Z(MCInst2_MC1_r1Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst2_MC1_r1Inst_XORInst_0_2_U3  ( .A(
        MCInst2_MC1_r1Inst_XORInst_0_2_n5 ), .B(
        MCInst2_MC1_r1Inst_XORInst_0_2_n4 ), .ZN(Feedback2[42]) );
  XNOR2_X1 MCInst2_MC1_r1Inst_XORInst_0_2_U2  ( .A(MCInst2_MC1_v3_1 [2]), 
        .B(MCInst2_MC1_v2_1 [2]), .ZN(MCInst2_MC1_r1Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst2_MC1_r1Inst_XORInst_0_2_U1  ( .A(MCInst2_MC1_v0_1 [2]), .B(
        MCInst2_MC1_v1_1 [2]), .Z(MCInst2_MC1_r1Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst2_MC1_r1Inst_XORInst_0_3_U3  ( .A(
        MCInst2_MC1_r1Inst_XORInst_0_3_n5 ), .B(
        MCInst2_MC1_r1Inst_XORInst_0_3_n4 ), .ZN(Feedback2[43]) );
  XNOR2_X1 MCInst2_MC1_r1Inst_XORInst_0_3_U2  ( .A(MCInst2_MC1_v3_1 [3]), 
        .B(MCInst2_MC1_v2_1 [3]), .ZN(MCInst2_MC1_r1Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst2_MC1_r1Inst_XORInst_0_3_U1  ( .A(MCInst2_MC1_v0_1 [3]), .B(
        MCInst2_MC1_v1_1 [3]), .Z(MCInst2_MC1_r1Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst2_MC1_r2Inst_XORInst_0_0_U3  ( .A(
        MCInst2_MC1_r2Inst_XORInst_0_0_n5 ), .B(
        MCInst2_MC1_r2Inst_XORInst_0_0_n4 ), .ZN(Feedback2[24]) );
  XNOR2_X1 MCInst2_MC1_r2Inst_XORInst_0_0_U2  ( .A(MCInst2_MC1_v3_2 [0]), 
        .B(MCInst2_MC1_v2_2 [0]), .ZN(MCInst2_MC1_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst2_MC1_r2Inst_XORInst_0_0_U1  ( .A(MCInst2_MC1_v0_2 [0]), .B(
        MCInst2_MC1_v1_2 [0]), .Z(MCInst2_MC1_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst2_MC1_r2Inst_XORInst_0_1_U3  ( .A(
        MCInst2_MC1_r2Inst_XORInst_0_1_n5 ), .B(
        MCInst2_MC1_r2Inst_XORInst_0_1_n4 ), .ZN(Feedback2[25]) );
  XNOR2_X1 MCInst2_MC1_r2Inst_XORInst_0_1_U2  ( .A(Red_MCInst2_MC1_v3_1[0] ), 
        .B(MCInst2_MC1_v2_2 [1]), .ZN(MCInst2_MC1_r2Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst2_MC1_r2Inst_XORInst_0_1_U1  ( .A(MCInst2_MC1_v0_2 [1]), .B(
        MCInst2_MC1_v1_2 [1]), .Z(MCInst2_MC1_r2Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst2_MC1_r2Inst_XORInst_0_2_U3  ( .A(
        MCInst2_MC1_r2Inst_XORInst_0_2_n5 ), .B(
        MCInst2_MC1_r2Inst_XORInst_0_2_n4 ), .ZN(Feedback2[26]) );
  XNOR2_X1 MCInst2_MC1_r2Inst_XORInst_0_2_U2  ( .A(MCInst2_MC1_v3_2 [2]), 
        .B(MCInst2_MC1_v2_2 [2]), .ZN(MCInst2_MC1_r2Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst2_MC1_r2Inst_XORInst_0_2_U1  ( .A(MCInst2_MC1_v0_2 [2]), .B(
        MCInst2_MC1_v1_2 [2]), .Z(MCInst2_MC1_r2Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst2_MC1_r2Inst_XORInst_0_3_U3  ( .A(
        MCInst2_MC1_r2Inst_XORInst_0_3_n5 ), .B(
        MCInst2_MC1_r2Inst_XORInst_0_3_n4 ), .ZN(Feedback2[27]) );
  XNOR2_X1 MCInst2_MC1_r2Inst_XORInst_0_3_U2  ( .A(MCInst2_MC1_v3_2 [3]), 
        .B(MCInst2_MC1_v2_2 [3]), .ZN(MCInst2_MC1_r2Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst2_MC1_r2Inst_XORInst_0_3_U1  ( .A(MCInst2_MC1_v0_2 [3]), .B(
        MCInst2_MC1_v1_2 [3]), .Z(MCInst2_MC1_r2Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst2_MC1_r3Inst_XORInst_0_0_U3  ( .A(
        MCInst2_MC1_r3Inst_XORInst_0_0_n5 ), .B(
        MCInst2_MC1_r3Inst_XORInst_0_0_n4 ), .ZN(Feedback2[8]) );
  XNOR2_X1 MCInst2_MC1_r3Inst_XORInst_0_0_U2  ( .A(MCInst2_MC1_v3_3 [0]), 
        .B(MCInst2_MC1_v2_3 [0]), .ZN(MCInst2_MC1_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst2_MC1_r3Inst_XORInst_0_0_U1  ( .A(MCInst2_MC1_v0_3 [0]), .B(
        MCInst2_MC1_v1_0 [3]), .Z(MCInst2_MC1_r3Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst2_MC1_r3Inst_XORInst_0_1_U3  ( .A(
        MCInst2_MC1_r3Inst_XORInst_0_1_n5 ), .B(
        MCInst2_MC1_r3Inst_XORInst_0_1_n4 ), .ZN(Feedback2[9]) );
  XNOR2_X1 MCInst2_MC1_r3Inst_XORInst_0_1_U2  ( .A(MCInst2_MC1_v3_3 [1]), 
        .B(MCInst2_MC1_v2_3 [1]), .ZN(MCInst2_MC1_r3Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst2_MC1_r3Inst_XORInst_0_1_U1  ( .A(MCInst2_MC1_v0_3 [1]), .B(
        MCInst2_MC1_v1_3 [1]), .Z(MCInst2_MC1_r3Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst2_MC1_r3Inst_XORInst_0_2_U3  ( .A(
        MCInst2_MC1_r3Inst_XORInst_0_2_n5 ), .B(
        MCInst2_MC1_r3Inst_XORInst_0_2_n4 ), .ZN(Feedback2[10]) );
  XNOR2_X1 MCInst2_MC1_r3Inst_XORInst_0_2_U2  ( .A(MCInst2_MC1_v3_3 [2]), 
        .B(MCInst2_MC1_v2_3 [2]), .ZN(MCInst2_MC1_r3Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst2_MC1_r3Inst_XORInst_0_2_U1  ( .A(MCInst2_MC1_v0_0 [3]), .B(
        MCInst2_MC1_v1_3 [2]), .Z(MCInst2_MC1_r3Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst2_MC1_r3Inst_XORInst_0_3_U3  ( .A(
        MCInst2_MC1_r3Inst_XORInst_0_3_n5 ), .B(
        MCInst2_MC1_r3Inst_XORInst_0_3_n4 ), .ZN(Feedback2[11]) );
  XNOR2_X1 MCInst2_MC1_r3Inst_XORInst_0_3_U2  ( .A(MCInst2_MC1_v3_3 [3]), 
        .B(MCInst2_MC1_v2_3 [3]), .ZN(MCInst2_MC1_r3Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst2_MC1_r3Inst_XORInst_0_3_U1  ( .A(MCInst2_MC1_v0_3 [3]), .B(
        Red_MCInst2_MC1_v1_1[0] ), .Z(MCInst2_MC1_r3Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst2_MC2_v0_2Inst_0_U4  ( .A(MCInst2_MC2_v0_2Inst_0_n2 ), .B(
        MCInst2_MC2_v0_0 [3]), .ZN(MCInst2_MC2_v0_2 [0]) );
  XNOR2_X1 MCInst2_MC2_v0_2Inst_0_U3  ( .A(MCInst2_MC2_v0_3 [0]), .B(
        Red_MCInst2_MC2_v0_1[0] ), .ZN(MCInst2_MC2_v0_2Inst_0_n2 ) );
  XOR2_X1 MCInst2_MC2_v1_1Inst_0_U3  ( .A(Red_MCInst2_MC2_v1_1[0] ), .B(
        MCInst2_MC2_v1_0 [3]), .Z(MCInst2_MC2_v1_1 [0]) );
  XNOR2_X1 MCInst2_MC2_v1_2Inst_0_U4  ( .A(MCInst2_MC2_v1_2Inst_0_n2 ), .B(
        Red_MCInst2_MC2_v1_1[0] ), .ZN(MCInst2_MC2_v1_2 [0]) );
  XNOR2_X1 MCInst2_MC2_v1_2Inst_0_U3  ( .A(MCInst2_MC2_v1_0 [3]), .B(
        MCInst2_MC2_v1_3 [2]), .ZN(MCInst2_MC2_v1_2Inst_0_n2 ) );
  XOR2_X1 MCInst2_MC2_v2_1Inst_0_U3  ( .A(MCInst2_MC2_v2_3 [1]), .B(
        MCInst2_MC2_v2_0 [3]), .Z(MCInst2_MC2_v2_1 [0]) );
  XOR2_X1 MCInst2_MC2_v2_2Inst_0_U3  ( .A(MCInst2_MC2_v2_0 [2]), .B(
        MCInst2_MC2_v2_0 [0]), .Z(MCInst2_MC2_v2_2 [0]) );
  XNOR2_X1 MCInst2_MC2_v2_3Inst_0_U5  ( .A(MCInst2_MC2_v2_3Inst_0_n4 ), .B(
        MCInst2_MC2_v2_3Inst_0_n3 ), .ZN(MCInst2_MC2_v2_3 [0]) );
  XNOR2_X1 MCInst2_MC2_v2_3Inst_0_U4  ( .A(MCInst2_MC2_v2_0 [2]), .B(
        MCInst2_MC2_v2_3 [1]), .ZN(MCInst2_MC2_v2_3Inst_0_n3 ) );
  XOR2_X1 MCInst2_MC2_v2_3Inst_0_U3  ( .A(MCInst2_MC2_v2_0 [3]), .B(
        MCInst2_MC2_v2_0 [0]), .Z(MCInst2_MC2_v2_3Inst_0_n4 ) );
  XOR2_X1 MCInst2_MC2_v3_1Inst_0_U3  ( .A(Red_MCInst2_MC2_v3_1[0] ), .B(
        MCInst2_MC2_v3_2 [2]), .Z(MCInst2_MC2_v3_1 [0]) );
  XOR2_X1 MCInst2_MC2_v3_2Inst_0_U3  ( .A(MCInst2_MC2_v3_2 [3]), .B(
        MCInst2_MC2_v3_0 [2]), .Z(MCInst2_MC2_v3_2 [0]) );
  XNOR2_X1 MCInst2_MC2_v3_3Inst_0_U4  ( .A(MCInst2_MC2_v3_3Inst_0_n2 ), .B(
        MCInst2_MC2_v3_0 [2]), .ZN(MCInst2_MC2_v3_3 [0]) );
  XNOR2_X1 MCInst2_MC2_v3_3Inst_0_U3  ( .A(MCInst2_MC2_v3_2 [2]), .B(
        MCInst2_MC2_v3_2 [3]), .ZN(MCInst2_MC2_v3_3Inst_0_n2 ) );
  XOR2_X1 MCInst2_MC2_v0_0Inst_1_U3  ( .A(MCInst2_MC2_v0_3 [3]), .B(
        MCInst2_MC2_v0_3 [0]), .Z(MCInst2_MC2_v0_0 [1]) );
  XOR2_X1 MCInst2_MC2_v0_1Inst_1_U3  ( .A(MCInst2_MC2_v0_0 [3]), .B(
        MCInst2_MC2_v0_3 [3]), .Z(MCInst2_MC2_v0_1 [1]) );
  XNOR2_X1 MCInst2_MC2_v0_2Inst_1_U4  ( .A(MCInst2_MC2_v0_2Inst_1_n2 ), .B(
        MCInst2_MC2_v0_3 [3]), .ZN(MCInst2_MC2_v0_2 [1]) );
  XNOR2_X1 MCInst2_MC2_v0_2Inst_1_U3  ( .A(MCInst2_MC2_v0_3 [0]), .B(
        Red_MCInst2_MC2_v0_1[0] ), .ZN(MCInst2_MC2_v0_2Inst_1_n2 ) );
  XOR2_X1 MCInst2_MC2_v0_3Inst_1_U3  ( .A(Red_MCInst2_MC2_v0_1[0] ), .B(
        MCInst2_MC2_v0_3 [0]), .Z(MCInst2_MC2_v0_3 [1]) );
  XOR2_X1 MCInst2_MC2_v1_1Inst_1_U3  ( .A(MCInst2_MC2_v1_0 [0]), .B(
        Red_MCInst2_MC2_v1_1[0] ), .Z(MCInst2_MC2_v1_1 [1]) );
  XOR2_X1 MCInst2_MC2_v1_2Inst_1_U3  ( .A(MCInst2_MC2_v1_0 [0]), .B(
        MCInst2_MC2_v1_3 [2]), .Z(MCInst2_MC2_v1_2 [1]) );
  XOR2_X1 MCInst2_MC2_v1_3Inst_1_U3  ( .A(MCInst2_MC2_v1_0 [0]), .B(
        MCInst2_MC2_v1_0 [3]), .Z(MCInst2_MC2_v1_3 [1]) );
  XOR2_X1 MCInst2_MC2_v2_0Inst_1_U3  ( .A(MCInst2_MC2_v2_3 [1]), .B(
        MCInst2_MC2_v2_0 [0]), .Z(MCInst2_MC2_v2_0 [1]) );
  XNOR2_X1 MCInst2_MC2_v2_1Inst_1_U4  ( .A(MCInst2_MC2_v2_1Inst_1_n2 ), .B(
        MCInst2_MC2_v2_0 [3]), .ZN(MCInst2_MC2_v2_1 [1]) );
  XNOR2_X1 MCInst2_MC2_v2_1Inst_1_U3  ( .A(MCInst2_MC2_v2_0 [0]), .B(
        MCInst2_MC2_v2_0 [2]), .ZN(MCInst2_MC2_v2_1Inst_1_n2 ) );
  XNOR2_X1 MCInst2_MC2_v2_2Inst_1_U5  ( .A(MCInst2_MC2_v2_2Inst_1_n4 ), .B(
        MCInst2_MC2_v2_2Inst_1_n3 ), .ZN(MCInst2_MC2_v2_2 [1]) );
  XNOR2_X1 MCInst2_MC2_v2_2Inst_1_U4  ( .A(MCInst2_MC2_v2_0 [2]), .B(
        MCInst2_MC2_v2_3 [1]), .ZN(MCInst2_MC2_v2_2Inst_1_n3 ) );
  XOR2_X1 MCInst2_MC2_v2_2Inst_1_U3  ( .A(MCInst2_MC2_v2_0 [3]), .B(
        MCInst2_MC2_v2_0 [0]), .Z(MCInst2_MC2_v2_2Inst_1_n4 ) );
  XOR2_X1 MCInst2_MC2_v3_0Inst_1_U3  ( .A(MCInst2_MC2_v3_2 [3]), .B(
        MCInst2_MC2_v3_2 [2]), .Z(MCInst2_MC2_v3_0 [1]) );
  XOR2_X1 MCInst2_MC2_v3_1Inst_1_U3  ( .A(MCInst2_MC2_v3_2 [3]), .B(
        Red_MCInst2_MC2_v3_1[0] ), .Z(MCInst2_MC2_v3_1 [1]) );
  XNOR2_X1 MCInst2_MC2_v3_3Inst_1_U4  ( .A(MCInst2_MC2_v3_3Inst_1_n2 ), .B(
        Red_MCInst2_MC2_v3_1[0] ), .ZN(MCInst2_MC2_v3_3 [1]) );
  XNOR2_X1 MCInst2_MC2_v3_3Inst_1_U3  ( .A(MCInst2_MC2_v3_2 [2]), .B(
        MCInst2_MC2_v3_2 [3]), .ZN(MCInst2_MC2_v3_3Inst_1_n2 ) );
  XOR2_X1 MCInst2_MC2_v0_0Inst_2_U3  ( .A(Red_MCInst2_MC2_v0_1[0] ), .B(
        MCInst2_MC2_v0_3 [0]), .Z(MCInst2_MC2_v0_0 [2]) );
  XOR2_X1 MCInst2_MC2_v0_1Inst_2_U3  ( .A(MCInst2_MC2_v0_3 [3]), .B(
        MCInst2_MC2_v0_3 [0]), .Z(MCInst2_MC2_v0_1 [2]) );
  XOR2_X1 MCInst2_MC2_v0_2Inst_2_U3  ( .A(MCInst2_MC2_v0_0 [3]), .B(
        MCInst2_MC2_v0_3 [0]), .Z(MCInst2_MC2_v0_2 [2]) );
  XNOR2_X1 MCInst2_MC2_v1_1Inst_2_U4  ( .A(MCInst2_MC2_v1_1Inst_2_n2 ), .B(
        MCInst2_MC2_v1_3 [2]), .ZN(MCInst2_MC2_v1_1 [2]) );
  XNOR2_X1 MCInst2_MC2_v1_1Inst_2_U3  ( .A(MCInst2_MC2_v1_0 [3]), .B(
        MCInst2_MC2_v1_0 [0]), .ZN(MCInst2_MC2_v1_1Inst_2_n2 ) );
  XNOR2_X1 MCInst2_MC2_v1_2Inst_2_U4  ( .A(MCInst2_MC2_v1_2Inst_2_n2 ), .B(
        MCInst2_MC2_v1_3 [2]), .ZN(MCInst2_MC2_v1_2 [2]) );
  XNOR2_X1 MCInst2_MC2_v1_2Inst_2_U3  ( .A(Red_MCInst2_MC2_v1_1[0] ), .B(
        MCInst2_MC2_v1_0 [0]), .ZN(MCInst2_MC2_v1_2Inst_2_n2 ) );
  XNOR2_X1 MCInst2_MC2_v2_1Inst_2_U4  ( .A(MCInst2_MC2_v2_1Inst_2_n2 ), .B(
        MCInst2_MC2_v2_0 [3]), .ZN(MCInst2_MC2_v2_1 [2]) );
  XNOR2_X1 MCInst2_MC2_v2_1Inst_2_U3  ( .A(MCInst2_MC2_v2_0 [0]), .B(
        MCInst2_MC2_v2_3 [1]), .ZN(MCInst2_MC2_v2_1Inst_2_n2 ) );
  XNOR2_X1 MCInst2_MC2_v2_2Inst_2_U4  ( .A(MCInst2_MC2_v2_2Inst_2_n2 ), .B(
        MCInst2_MC2_v2_0 [3]), .ZN(MCInst2_MC2_v2_2 [2]) );
  XNOR2_X1 MCInst2_MC2_v2_2Inst_2_U3  ( .A(MCInst2_MC2_v2_0 [0]), .B(
        MCInst2_MC2_v2_0 [2]), .ZN(MCInst2_MC2_v2_2Inst_2_n2 ) );
  XOR2_X1 MCInst2_MC2_v2_3Inst_2_U3  ( .A(MCInst2_MC2_v2_3 [1]), .B(
        MCInst2_MC2_v2_0 [2]), .Z(MCInst2_MC2_v2_3 [2]) );
  XNOR2_X1 MCInst2_MC2_v3_1Inst_2_U4  ( .A(MCInst2_MC2_v3_1Inst_2_n2 ), .B(
        MCInst2_MC2_v3_0 [2]), .ZN(MCInst2_MC2_v3_1 [2]) );
  XNOR2_X1 MCInst2_MC2_v3_1Inst_2_U3  ( .A(MCInst2_MC2_v3_2 [2]), .B(
        MCInst2_MC2_v3_2 [3]), .ZN(MCInst2_MC2_v3_1Inst_2_n2 ) );
  XOR2_X1 MCInst2_MC2_v3_3Inst_2_U3  ( .A(MCInst2_MC2_v3_0 [2]), .B(
        MCInst2_MC2_v3_2 [2]), .Z(MCInst2_MC2_v3_3 [2]) );
  XOR2_X1 MCInst2_MC2_v0_1Inst_3_U3  ( .A(Red_MCInst2_MC2_v0_1[0] ), .B(
        MCInst2_MC2_v0_3 [0]), .Z(MCInst2_MC2_v0_1 [3]) );
  XOR2_X1 MCInst2_MC2_v0_2Inst_3_U3  ( .A(Red_MCInst2_MC2_v0_1[0] ), .B(
        MCInst2_MC2_v0_3 [3]), .Z(MCInst2_MC2_v0_2 [3]) );
  XOR2_X1 MCInst2_MC2_v1_1Inst_3_U3  ( .A(MCInst2_MC2_v1_3 [2]), .B(
        Red_MCInst2_MC2_v1_1[0] ), .Z(MCInst2_MC2_v1_1 [3]) );
  XNOR2_X1 MCInst2_MC2_v1_2Inst_3_U5  ( .A(MCInst2_MC2_v1_2Inst_3_n4 ), .B(
        MCInst2_MC2_v1_2Inst_3_n3 ), .ZN(MCInst2_MC2_v1_2 [3]) );
  XNOR2_X1 MCInst2_MC2_v1_2Inst_3_U4  ( .A(MCInst2_MC2_v1_3 [2]), .B(
        MCInst2_MC2_v1_0 [0]), .ZN(MCInst2_MC2_v1_2Inst_3_n3 ) );
  XOR2_X1 MCInst2_MC2_v1_2Inst_3_U3  ( .A(Red_MCInst2_MC2_v1_1[0] ), .B(
        MCInst2_MC2_v1_0 [3]), .Z(MCInst2_MC2_v1_2Inst_3_n4 ) );
  XOR2_X1 MCInst2_MC2_v2_1Inst_3_U3  ( .A(MCInst2_MC2_v2_0 [2]), .B(
        MCInst2_MC2_v2_0 [0]), .Z(MCInst2_MC2_v2_1 [3]) );
  XNOR2_X1 MCInst2_MC2_v2_2Inst_3_U4  ( .A(MCInst2_MC2_v2_2Inst_3_n2 ), .B(
        MCInst2_MC2_v2_0 [3]), .ZN(MCInst2_MC2_v2_2 [3]) );
  XNOR2_X1 MCInst2_MC2_v2_2Inst_3_U3  ( .A(MCInst2_MC2_v2_0 [0]), .B(
        MCInst2_MC2_v2_3 [1]), .ZN(MCInst2_MC2_v2_2Inst_3_n2 ) );
  XNOR2_X1 MCInst2_MC2_v2_3Inst_3_U4  ( .A(MCInst2_MC2_v2_3Inst_3_n2 ), .B(
        MCInst2_MC2_v2_0 [2]), .ZN(MCInst2_MC2_v2_3 [3]) );
  XNOR2_X1 MCInst2_MC2_v2_3Inst_3_U3  ( .A(MCInst2_MC2_v2_0 [3]), .B(
        MCInst2_MC2_v2_3 [1]), .ZN(MCInst2_MC2_v2_3Inst_3_n2 ) );
  XOR2_X1 MCInst2_MC2_v3_1Inst_3_U3  ( .A(MCInst2_MC2_v3_0 [2]), .B(
        Red_MCInst2_MC2_v3_1[0] ), .Z(MCInst2_MC2_v3_1 [3]) );
  XOR2_X1 MCInst2_MC2_v3_3Inst_3_U3  ( .A(MCInst2_MC2_v3_2 [3]), .B(
        Red_MCInst2_MC2_v3_1[0] ), .Z(MCInst2_MC2_v3_3 [3]) );
  XNOR2_X1 MCInst2_MC2_r0Inst_XORInst_0_0_U3  ( .A(
        MCInst2_MC2_r0Inst_XORInst_0_0_n5 ), .B(
        MCInst2_MC2_r0Inst_XORInst_0_0_n4 ), .ZN(Feedback2[52]) );
  XNOR2_X1 MCInst2_MC2_r0Inst_XORInst_0_0_U2  ( .A(MCInst2_MC2_v3_2 [2]), 
        .B(MCInst2_MC2_v2_0 [0]), .ZN(MCInst2_MC2_r0Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst2_MC2_r0Inst_XORInst_0_0_U1  ( .A(MCInst2_MC2_v0_3 [3]), .B(
        MCInst2_MC2_v1_0 [0]), .Z(MCInst2_MC2_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst2_MC2_r0Inst_XORInst_0_1_U3  ( .A(
        MCInst2_MC2_r0Inst_XORInst_0_1_n5 ), .B(
        MCInst2_MC2_r0Inst_XORInst_0_1_n4 ), .ZN(Feedback2[53]) );
  XNOR2_X1 MCInst2_MC2_r0Inst_XORInst_0_1_U2  ( .A(MCInst2_MC2_v3_0 [1]), 
        .B(MCInst2_MC2_v2_0 [1]), .ZN(MCInst2_MC2_r0Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst2_MC2_r0Inst_XORInst_0_1_U1  ( .A(MCInst2_MC2_v0_0 [1]), .B(
        MCInst2_MC2_v1_3 [2]), .Z(MCInst2_MC2_r0Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst2_MC2_r0Inst_XORInst_0_2_U3  ( .A(
        MCInst2_MC2_r0Inst_XORInst_0_2_n5 ), .B(
        MCInst2_MC2_r0Inst_XORInst_0_2_n4 ), .ZN(Feedback2[54]) );
  XNOR2_X1 MCInst2_MC2_r0Inst_XORInst_0_2_U2  ( .A(MCInst2_MC2_v3_0 [2]), 
        .B(MCInst2_MC2_v2_0 [2]), .ZN(MCInst2_MC2_r0Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst2_MC2_r0Inst_XORInst_0_2_U1  ( .A(MCInst2_MC2_v0_0 [2]), .B(
        Red_MCInst2_MC2_v1_1[0] ), .Z(MCInst2_MC2_r0Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst2_MC2_r0Inst_XORInst_0_3_U3  ( .A(
        MCInst2_MC2_r0Inst_XORInst_0_3_n5 ), .B(
        MCInst2_MC2_r0Inst_XORInst_0_3_n4 ), .ZN(Feedback2[55]) );
  XNOR2_X1 MCInst2_MC2_r0Inst_XORInst_0_3_U2  ( .A(Red_MCInst2_MC2_v3_1[0] ), 
        .B(MCInst2_MC2_v2_0 [3]), .ZN(MCInst2_MC2_r0Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst2_MC2_r0Inst_XORInst_0_3_U1  ( .A(MCInst2_MC2_v0_0 [3]), .B(
        MCInst2_MC2_v1_0 [3]), .Z(MCInst2_MC2_r0Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst2_MC2_r1Inst_XORInst_0_0_U3  ( .A(
        MCInst2_MC2_r1Inst_XORInst_0_0_n5 ), .B(
        MCInst2_MC2_r1Inst_XORInst_0_0_n4 ), .ZN(Feedback2[36]) );
  XNOR2_X1 MCInst2_MC2_r1Inst_XORInst_0_0_U2  ( .A(MCInst2_MC2_v3_1 [0]), 
        .B(MCInst2_MC2_v2_1 [0]), .ZN(MCInst2_MC2_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst2_MC2_r1Inst_XORInst_0_0_U1  ( .A(MCInst2_MC2_v0_0 [3]), .B(
        MCInst2_MC2_v1_1 [0]), .Z(MCInst2_MC2_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst2_MC2_r1Inst_XORInst_0_1_U3  ( .A(
        MCInst2_MC2_r1Inst_XORInst_0_1_n5 ), .B(
        MCInst2_MC2_r1Inst_XORInst_0_1_n4 ), .ZN(Feedback2[37]) );
  XNOR2_X1 MCInst2_MC2_r1Inst_XORInst_0_1_U2  ( .A(MCInst2_MC2_v3_1 [1]), 
        .B(MCInst2_MC2_v2_1 [1]), .ZN(MCInst2_MC2_r1Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst2_MC2_r1Inst_XORInst_0_1_U1  ( .A(MCInst2_MC2_v0_1 [1]), .B(
        MCInst2_MC2_v1_1 [1]), .Z(MCInst2_MC2_r1Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst2_MC2_r1Inst_XORInst_0_2_U3  ( .A(
        MCInst2_MC2_r1Inst_XORInst_0_2_n5 ), .B(
        MCInst2_MC2_r1Inst_XORInst_0_2_n4 ), .ZN(Feedback2[38]) );
  XNOR2_X1 MCInst2_MC2_r1Inst_XORInst_0_2_U2  ( .A(MCInst2_MC2_v3_1 [2]), 
        .B(MCInst2_MC2_v2_1 [2]), .ZN(MCInst2_MC2_r1Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst2_MC2_r1Inst_XORInst_0_2_U1  ( .A(MCInst2_MC2_v0_1 [2]), .B(
        MCInst2_MC2_v1_1 [2]), .Z(MCInst2_MC2_r1Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst2_MC2_r1Inst_XORInst_0_3_U3  ( .A(
        MCInst2_MC2_r1Inst_XORInst_0_3_n5 ), .B(
        MCInst2_MC2_r1Inst_XORInst_0_3_n4 ), .ZN(Feedback2[39]) );
  XNOR2_X1 MCInst2_MC2_r1Inst_XORInst_0_3_U2  ( .A(MCInst2_MC2_v3_1 [3]), 
        .B(MCInst2_MC2_v2_1 [3]), .ZN(MCInst2_MC2_r1Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst2_MC2_r1Inst_XORInst_0_3_U1  ( .A(MCInst2_MC2_v0_1 [3]), .B(
        MCInst2_MC2_v1_1 [3]), .Z(MCInst2_MC2_r1Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst2_MC2_r2Inst_XORInst_0_0_U3  ( .A(
        MCInst2_MC2_r2Inst_XORInst_0_0_n5 ), .B(
        MCInst2_MC2_r2Inst_XORInst_0_0_n4 ), .ZN(Feedback2[20]) );
  XNOR2_X1 MCInst2_MC2_r2Inst_XORInst_0_0_U2  ( .A(MCInst2_MC2_v3_2 [0]), 
        .B(MCInst2_MC2_v2_2 [0]), .ZN(MCInst2_MC2_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst2_MC2_r2Inst_XORInst_0_0_U1  ( .A(MCInst2_MC2_v0_2 [0]), .B(
        MCInst2_MC2_v1_2 [0]), .Z(MCInst2_MC2_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst2_MC2_r2Inst_XORInst_0_1_U3  ( .A(
        MCInst2_MC2_r2Inst_XORInst_0_1_n5 ), .B(
        MCInst2_MC2_r2Inst_XORInst_0_1_n4 ), .ZN(Feedback2[21]) );
  XNOR2_X1 MCInst2_MC2_r2Inst_XORInst_0_1_U2  ( .A(Red_MCInst2_MC2_v3_1[0] ), 
        .B(MCInst2_MC2_v2_2 [1]), .ZN(MCInst2_MC2_r2Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst2_MC2_r2Inst_XORInst_0_1_U1  ( .A(MCInst2_MC2_v0_2 [1]), .B(
        MCInst2_MC2_v1_2 [1]), .Z(MCInst2_MC2_r2Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst2_MC2_r2Inst_XORInst_0_2_U3  ( .A(
        MCInst2_MC2_r2Inst_XORInst_0_2_n5 ), .B(
        MCInst2_MC2_r2Inst_XORInst_0_2_n4 ), .ZN(Feedback2[22]) );
  XNOR2_X1 MCInst2_MC2_r2Inst_XORInst_0_2_U2  ( .A(MCInst2_MC2_v3_2 [2]), 
        .B(MCInst2_MC2_v2_2 [2]), .ZN(MCInst2_MC2_r2Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst2_MC2_r2Inst_XORInst_0_2_U1  ( .A(MCInst2_MC2_v0_2 [2]), .B(
        MCInst2_MC2_v1_2 [2]), .Z(MCInst2_MC2_r2Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst2_MC2_r2Inst_XORInst_0_3_U3  ( .A(
        MCInst2_MC2_r2Inst_XORInst_0_3_n5 ), .B(
        MCInst2_MC2_r2Inst_XORInst_0_3_n4 ), .ZN(Feedback2[23]) );
  XNOR2_X1 MCInst2_MC2_r2Inst_XORInst_0_3_U2  ( .A(MCInst2_MC2_v3_2 [3]), 
        .B(MCInst2_MC2_v2_2 [3]), .ZN(MCInst2_MC2_r2Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst2_MC2_r2Inst_XORInst_0_3_U1  ( .A(MCInst2_MC2_v0_2 [3]), .B(
        MCInst2_MC2_v1_2 [3]), .Z(MCInst2_MC2_r2Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst2_MC2_r3Inst_XORInst_0_0_U3  ( .A(
        MCInst2_MC2_r3Inst_XORInst_0_0_n5 ), .B(
        MCInst2_MC2_r3Inst_XORInst_0_0_n4 ), .ZN(Feedback2[4]) );
  XNOR2_X1 MCInst2_MC2_r3Inst_XORInst_0_0_U2  ( .A(MCInst2_MC2_v3_3 [0]), 
        .B(MCInst2_MC2_v2_3 [0]), .ZN(MCInst2_MC2_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst2_MC2_r3Inst_XORInst_0_0_U1  ( .A(MCInst2_MC2_v0_3 [0]), .B(
        MCInst2_MC2_v1_0 [3]), .Z(MCInst2_MC2_r3Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst2_MC2_r3Inst_XORInst_0_1_U3  ( .A(
        MCInst2_MC2_r3Inst_XORInst_0_1_n5 ), .B(
        MCInst2_MC2_r3Inst_XORInst_0_1_n4 ), .ZN(Feedback2[5]) );
  XNOR2_X1 MCInst2_MC2_r3Inst_XORInst_0_1_U2  ( .A(MCInst2_MC2_v3_3 [1]), 
        .B(MCInst2_MC2_v2_3 [1]), .ZN(MCInst2_MC2_r3Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst2_MC2_r3Inst_XORInst_0_1_U1  ( .A(MCInst2_MC2_v0_3 [1]), .B(
        MCInst2_MC2_v1_3 [1]), .Z(MCInst2_MC2_r3Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst2_MC2_r3Inst_XORInst_0_2_U3  ( .A(
        MCInst2_MC2_r3Inst_XORInst_0_2_n5 ), .B(
        MCInst2_MC2_r3Inst_XORInst_0_2_n4 ), .ZN(Feedback2[6]) );
  XNOR2_X1 MCInst2_MC2_r3Inst_XORInst_0_2_U2  ( .A(MCInst2_MC2_v3_3 [2]), 
        .B(MCInst2_MC2_v2_3 [2]), .ZN(MCInst2_MC2_r3Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst2_MC2_r3Inst_XORInst_0_2_U1  ( .A(MCInst2_MC2_v0_0 [3]), .B(
        MCInst2_MC2_v1_3 [2]), .Z(MCInst2_MC2_r3Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst2_MC2_r3Inst_XORInst_0_3_U3  ( .A(
        MCInst2_MC2_r3Inst_XORInst_0_3_n5 ), .B(
        MCInst2_MC2_r3Inst_XORInst_0_3_n4 ), .ZN(Feedback2[7]) );
  XNOR2_X1 MCInst2_MC2_r3Inst_XORInst_0_3_U2  ( .A(MCInst2_MC2_v3_3 [3]), 
        .B(MCInst2_MC2_v2_3 [3]), .ZN(MCInst2_MC2_r3Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst2_MC2_r3Inst_XORInst_0_3_U1  ( .A(MCInst2_MC2_v0_3 [3]), .B(
        Red_MCInst2_MC2_v1_1[0] ), .Z(MCInst2_MC2_r3Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst2_MC3_v0_2Inst_0_U4  ( .A(MCInst2_MC3_v0_2Inst_0_n2 ), .B(
        MCInst2_MC3_v0_0 [3]), .ZN(MCInst2_MC3_v0_2 [0]) );
  XNOR2_X1 MCInst2_MC3_v0_2Inst_0_U3  ( .A(MCInst2_MC3_v0_3 [0]), .B(
        Red_MCInst2_MC3_v0_1[0] ), .ZN(MCInst2_MC3_v0_2Inst_0_n2 ) );
  XOR2_X1 MCInst2_MC3_v1_1Inst_0_U3  ( .A(Red_MCInst2_MC3_v1_1[0] ), .B(
        MCInst2_MC3_v1_0 [3]), .Z(MCInst2_MC3_v1_1 [0]) );
  XNOR2_X1 MCInst2_MC3_v1_2Inst_0_U4  ( .A(MCInst2_MC3_v1_2Inst_0_n2 ), .B(
        Red_MCInst2_MC3_v1_1[0] ), .ZN(MCInst2_MC3_v1_2 [0]) );
  XNOR2_X1 MCInst2_MC3_v1_2Inst_0_U3  ( .A(MCInst2_MC3_v1_0 [3]), .B(
        MCInst2_MC3_v1_3 [2]), .ZN(MCInst2_MC3_v1_2Inst_0_n2 ) );
  XOR2_X1 MCInst2_MC3_v2_1Inst_0_U3  ( .A(MCInst2_MC3_v2_3 [1]), .B(
        MCInst2_MC3_v2_0 [3]), .Z(MCInst2_MC3_v2_1 [0]) );
  XOR2_X1 MCInst2_MC3_v2_2Inst_0_U3  ( .A(MCInst2_MC3_v2_0 [2]), .B(
        MCInst2_MC3_v2_0 [0]), .Z(MCInst2_MC3_v2_2 [0]) );
  XNOR2_X1 MCInst2_MC3_v2_3Inst_0_U5  ( .A(MCInst2_MC3_v2_3Inst_0_n4 ), .B(
        MCInst2_MC3_v2_3Inst_0_n3 ), .ZN(MCInst2_MC3_v2_3 [0]) );
  XNOR2_X1 MCInst2_MC3_v2_3Inst_0_U4  ( .A(MCInst2_MC3_v2_0 [2]), .B(
        MCInst2_MC3_v2_3 [1]), .ZN(MCInst2_MC3_v2_3Inst_0_n3 ) );
  XOR2_X1 MCInst2_MC3_v2_3Inst_0_U3  ( .A(MCInst2_MC3_v2_0 [3]), .B(
        MCInst2_MC3_v2_0 [0]), .Z(MCInst2_MC3_v2_3Inst_0_n4 ) );
  XOR2_X1 MCInst2_MC3_v3_1Inst_0_U3  ( .A(Red_MCInst2_MC3_v3_1[0] ), .B(
        MCInst2_MC3_v3_2 [2]), .Z(MCInst2_MC3_v3_1 [0]) );
  XOR2_X1 MCInst2_MC3_v3_2Inst_0_U3  ( .A(MCInst2_MC3_v3_2 [3]), .B(
        MCInst2_MC3_v3_0 [2]), .Z(MCInst2_MC3_v3_2 [0]) );
  XNOR2_X1 MCInst2_MC3_v3_3Inst_0_U4  ( .A(MCInst2_MC3_v3_3Inst_0_n2 ), .B(
        MCInst2_MC3_v3_0 [2]), .ZN(MCInst2_MC3_v3_3 [0]) );
  XNOR2_X1 MCInst2_MC3_v3_3Inst_0_U3  ( .A(MCInst2_MC3_v3_2 [2]), .B(
        MCInst2_MC3_v3_2 [3]), .ZN(MCInst2_MC3_v3_3Inst_0_n2 ) );
  XOR2_X1 MCInst2_MC3_v0_0Inst_1_U3  ( .A(MCInst2_MC3_v0_3 [3]), .B(
        MCInst2_MC3_v0_3 [0]), .Z(MCInst2_MC3_v0_0 [1]) );
  XOR2_X1 MCInst2_MC3_v0_1Inst_1_U3  ( .A(MCInst2_MC3_v0_0 [3]), .B(
        MCInst2_MC3_v0_3 [3]), .Z(MCInst2_MC3_v0_1 [1]) );
  XNOR2_X1 MCInst2_MC3_v0_2Inst_1_U4  ( .A(MCInst2_MC3_v0_2Inst_1_n2 ), .B(
        MCInst2_MC3_v0_3 [3]), .ZN(MCInst2_MC3_v0_2 [1]) );
  XNOR2_X1 MCInst2_MC3_v0_2Inst_1_U3  ( .A(MCInst2_MC3_v0_3 [0]), .B(
        Red_MCInst2_MC3_v0_1[0] ), .ZN(MCInst2_MC3_v0_2Inst_1_n2 ) );
  XOR2_X1 MCInst2_MC3_v0_3Inst_1_U3  ( .A(Red_MCInst2_MC3_v0_1[0] ), .B(
        MCInst2_MC3_v0_3 [0]), .Z(MCInst2_MC3_v0_3 [1]) );
  XOR2_X1 MCInst2_MC3_v1_1Inst_1_U3  ( .A(MCInst2_MC3_v1_0 [0]), .B(
        Red_MCInst2_MC3_v1_1[0] ), .Z(MCInst2_MC3_v1_1 [1]) );
  XOR2_X1 MCInst2_MC3_v1_2Inst_1_U3  ( .A(MCInst2_MC3_v1_0 [0]), .B(
        MCInst2_MC3_v1_3 [2]), .Z(MCInst2_MC3_v1_2 [1]) );
  XOR2_X1 MCInst2_MC3_v1_3Inst_1_U3  ( .A(MCInst2_MC3_v1_0 [0]), .B(
        MCInst2_MC3_v1_0 [3]), .Z(MCInst2_MC3_v1_3 [1]) );
  XOR2_X1 MCInst2_MC3_v2_0Inst_1_U3  ( .A(MCInst2_MC3_v2_3 [1]), .B(
        MCInst2_MC3_v2_0 [0]), .Z(MCInst2_MC3_v2_0 [1]) );
  XNOR2_X1 MCInst2_MC3_v2_1Inst_1_U4  ( .A(MCInst2_MC3_v2_1Inst_1_n2 ), .B(
        MCInst2_MC3_v2_0 [3]), .ZN(MCInst2_MC3_v2_1 [1]) );
  XNOR2_X1 MCInst2_MC3_v2_1Inst_1_U3  ( .A(MCInst2_MC3_v2_0 [0]), .B(
        MCInst2_MC3_v2_0 [2]), .ZN(MCInst2_MC3_v2_1Inst_1_n2 ) );
  XNOR2_X1 MCInst2_MC3_v2_2Inst_1_U5  ( .A(MCInst2_MC3_v2_2Inst_1_n4 ), .B(
        MCInst2_MC3_v2_2Inst_1_n3 ), .ZN(MCInst2_MC3_v2_2 [1]) );
  XNOR2_X1 MCInst2_MC3_v2_2Inst_1_U4  ( .A(MCInst2_MC3_v2_0 [2]), .B(
        MCInst2_MC3_v2_3 [1]), .ZN(MCInst2_MC3_v2_2Inst_1_n3 ) );
  XOR2_X1 MCInst2_MC3_v2_2Inst_1_U3  ( .A(MCInst2_MC3_v2_0 [3]), .B(
        MCInst2_MC3_v2_0 [0]), .Z(MCInst2_MC3_v2_2Inst_1_n4 ) );
  XOR2_X1 MCInst2_MC3_v3_0Inst_1_U3  ( .A(MCInst2_MC3_v3_2 [3]), .B(
        MCInst2_MC3_v3_2 [2]), .Z(MCInst2_MC3_v3_0 [1]) );
  XOR2_X1 MCInst2_MC3_v3_1Inst_1_U3  ( .A(MCInst2_MC3_v3_2 [3]), .B(
        Red_MCInst2_MC3_v3_1[0] ), .Z(MCInst2_MC3_v3_1 [1]) );
  XNOR2_X1 MCInst2_MC3_v3_3Inst_1_U4  ( .A(MCInst2_MC3_v3_3Inst_1_n2 ), .B(
        Red_MCInst2_MC3_v3_1[0] ), .ZN(MCInst2_MC3_v3_3 [1]) );
  XNOR2_X1 MCInst2_MC3_v3_3Inst_1_U3  ( .A(MCInst2_MC3_v3_2 [2]), .B(
        MCInst2_MC3_v3_2 [3]), .ZN(MCInst2_MC3_v3_3Inst_1_n2 ) );
  XOR2_X1 MCInst2_MC3_v0_0Inst_2_U3  ( .A(Red_MCInst2_MC3_v0_1[0] ), .B(
        MCInst2_MC3_v0_3 [0]), .Z(MCInst2_MC3_v0_0 [2]) );
  XOR2_X1 MCInst2_MC3_v0_1Inst_2_U3  ( .A(MCInst2_MC3_v0_3 [3]), .B(
        MCInst2_MC3_v0_3 [0]), .Z(MCInst2_MC3_v0_1 [2]) );
  XOR2_X1 MCInst2_MC3_v0_2Inst_2_U3  ( .A(MCInst2_MC3_v0_0 [3]), .B(
        MCInst2_MC3_v0_3 [0]), .Z(MCInst2_MC3_v0_2 [2]) );
  XNOR2_X1 MCInst2_MC3_v1_1Inst_2_U4  ( .A(MCInst2_MC3_v1_1Inst_2_n2 ), .B(
        MCInst2_MC3_v1_3 [2]), .ZN(MCInst2_MC3_v1_1 [2]) );
  XNOR2_X1 MCInst2_MC3_v1_1Inst_2_U3  ( .A(MCInst2_MC3_v1_0 [3]), .B(
        MCInst2_MC3_v1_0 [0]), .ZN(MCInst2_MC3_v1_1Inst_2_n2 ) );
  XNOR2_X1 MCInst2_MC3_v1_2Inst_2_U4  ( .A(MCInst2_MC3_v1_2Inst_2_n2 ), .B(
        MCInst2_MC3_v1_3 [2]), .ZN(MCInst2_MC3_v1_2 [2]) );
  XNOR2_X1 MCInst2_MC3_v1_2Inst_2_U3  ( .A(Red_MCInst2_MC3_v1_1[0] ), .B(
        MCInst2_MC3_v1_0 [0]), .ZN(MCInst2_MC3_v1_2Inst_2_n2 ) );
  XNOR2_X1 MCInst2_MC3_v2_1Inst_2_U4  ( .A(MCInst2_MC3_v2_1Inst_2_n2 ), .B(
        MCInst2_MC3_v2_0 [3]), .ZN(MCInst2_MC3_v2_1 [2]) );
  XNOR2_X1 MCInst2_MC3_v2_1Inst_2_U3  ( .A(MCInst2_MC3_v2_0 [0]), .B(
        MCInst2_MC3_v2_3 [1]), .ZN(MCInst2_MC3_v2_1Inst_2_n2 ) );
  XNOR2_X1 MCInst2_MC3_v2_2Inst_2_U4  ( .A(MCInst2_MC3_v2_2Inst_2_n2 ), .B(
        MCInst2_MC3_v2_0 [3]), .ZN(MCInst2_MC3_v2_2 [2]) );
  XNOR2_X1 MCInst2_MC3_v2_2Inst_2_U3  ( .A(MCInst2_MC3_v2_0 [0]), .B(
        MCInst2_MC3_v2_0 [2]), .ZN(MCInst2_MC3_v2_2Inst_2_n2 ) );
  XOR2_X1 MCInst2_MC3_v2_3Inst_2_U3  ( .A(MCInst2_MC3_v2_3 [1]), .B(
        MCInst2_MC3_v2_0 [2]), .Z(MCInst2_MC3_v2_3 [2]) );
  XNOR2_X1 MCInst2_MC3_v3_1Inst_2_U4  ( .A(MCInst2_MC3_v3_1Inst_2_n2 ), .B(
        MCInst2_MC3_v3_0 [2]), .ZN(MCInst2_MC3_v3_1 [2]) );
  XNOR2_X1 MCInst2_MC3_v3_1Inst_2_U3  ( .A(MCInst2_MC3_v3_2 [2]), .B(
        MCInst2_MC3_v3_2 [3]), .ZN(MCInst2_MC3_v3_1Inst_2_n2 ) );
  XOR2_X1 MCInst2_MC3_v3_3Inst_2_U3  ( .A(MCInst2_MC3_v3_0 [2]), .B(
        MCInst2_MC3_v3_2 [2]), .Z(MCInst2_MC3_v3_3 [2]) );
  XOR2_X1 MCInst2_MC3_v0_1Inst_3_U3  ( .A(Red_MCInst2_MC3_v0_1[0] ), .B(
        MCInst2_MC3_v0_3 [0]), .Z(MCInst2_MC3_v0_1 [3]) );
  XOR2_X1 MCInst2_MC3_v0_2Inst_3_U3  ( .A(Red_MCInst2_MC3_v0_1[0] ), .B(
        MCInst2_MC3_v0_3 [3]), .Z(MCInst2_MC3_v0_2 [3]) );
  XOR2_X1 MCInst2_MC3_v1_1Inst_3_U3  ( .A(MCInst2_MC3_v1_3 [2]), .B(
        Red_MCInst2_MC3_v1_1[0] ), .Z(MCInst2_MC3_v1_1 [3]) );
  XNOR2_X1 MCInst2_MC3_v1_2Inst_3_U5  ( .A(MCInst2_MC3_v1_2Inst_3_n4 ), .B(
        MCInst2_MC3_v1_2Inst_3_n3 ), .ZN(MCInst2_MC3_v1_2 [3]) );
  XNOR2_X1 MCInst2_MC3_v1_2Inst_3_U4  ( .A(MCInst2_MC3_v1_3 [2]), .B(
        MCInst2_MC3_v1_0 [0]), .ZN(MCInst2_MC3_v1_2Inst_3_n3 ) );
  XOR2_X1 MCInst2_MC3_v1_2Inst_3_U3  ( .A(Red_MCInst2_MC3_v1_1[0] ), .B(
        MCInst2_MC3_v1_0 [3]), .Z(MCInst2_MC3_v1_2Inst_3_n4 ) );
  XOR2_X1 MCInst2_MC3_v2_1Inst_3_U3  ( .A(MCInst2_MC3_v2_0 [2]), .B(
        MCInst2_MC3_v2_0 [0]), .Z(MCInst2_MC3_v2_1 [3]) );
  XNOR2_X1 MCInst2_MC3_v2_2Inst_3_U4  ( .A(MCInst2_MC3_v2_2Inst_3_n2 ), .B(
        MCInst2_MC3_v2_0 [3]), .ZN(MCInst2_MC3_v2_2 [3]) );
  XNOR2_X1 MCInst2_MC3_v2_2Inst_3_U3  ( .A(MCInst2_MC3_v2_0 [0]), .B(
        MCInst2_MC3_v2_3 [1]), .ZN(MCInst2_MC3_v2_2Inst_3_n2 ) );
  XNOR2_X1 MCInst2_MC3_v2_3Inst_3_U4  ( .A(MCInst2_MC3_v2_3Inst_3_n2 ), .B(
        MCInst2_MC3_v2_0 [2]), .ZN(MCInst2_MC3_v2_3 [3]) );
  XNOR2_X1 MCInst2_MC3_v2_3Inst_3_U3  ( .A(MCInst2_MC3_v2_0 [3]), .B(
        MCInst2_MC3_v2_3 [1]), .ZN(MCInst2_MC3_v2_3Inst_3_n2 ) );
  XOR2_X1 MCInst2_MC3_v3_1Inst_3_U3  ( .A(MCInst2_MC3_v3_0 [2]), .B(
        Red_MCInst2_MC3_v3_1[0] ), .Z(MCInst2_MC3_v3_1 [3]) );
  XOR2_X1 MCInst2_MC3_v3_3Inst_3_U3  ( .A(MCInst2_MC3_v3_2 [3]), .B(
        Red_MCInst2_MC3_v3_1[0] ), .Z(MCInst2_MC3_v3_3 [3]) );
  XNOR2_X1 MCInst2_MC3_r0Inst_XORInst_0_0_U3  ( .A(
        MCInst2_MC3_r0Inst_XORInst_0_0_n5 ), .B(
        MCInst2_MC3_r0Inst_XORInst_0_0_n4 ), .ZN(Feedback2[48]) );
  XNOR2_X1 MCInst2_MC3_r0Inst_XORInst_0_0_U2  ( .A(MCInst2_MC3_v3_2 [2]), 
        .B(MCInst2_MC3_v2_0 [0]), .ZN(MCInst2_MC3_r0Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst2_MC3_r0Inst_XORInst_0_0_U1  ( .A(MCInst2_MC3_v0_3 [3]), .B(
        MCInst2_MC3_v1_0 [0]), .Z(MCInst2_MC3_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst2_MC3_r0Inst_XORInst_0_1_U3  ( .A(
        MCInst2_MC3_r0Inst_XORInst_0_1_n5 ), .B(
        MCInst2_MC3_r0Inst_XORInst_0_1_n4 ), .ZN(Feedback2[49]) );
  XNOR2_X1 MCInst2_MC3_r0Inst_XORInst_0_1_U2  ( .A(MCInst2_MC3_v3_0 [1]), 
        .B(MCInst2_MC3_v2_0 [1]), .ZN(MCInst2_MC3_r0Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst2_MC3_r0Inst_XORInst_0_1_U1  ( .A(MCInst2_MC3_v0_0 [1]), .B(
        MCInst2_MC3_v1_3 [2]), .Z(MCInst2_MC3_r0Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst2_MC3_r0Inst_XORInst_0_2_U3  ( .A(
        MCInst2_MC3_r0Inst_XORInst_0_2_n5 ), .B(
        MCInst2_MC3_r0Inst_XORInst_0_2_n4 ), .ZN(Feedback2[50]) );
  XNOR2_X1 MCInst2_MC3_r0Inst_XORInst_0_2_U2  ( .A(MCInst2_MC3_v3_0 [2]), 
        .B(MCInst2_MC3_v2_0 [2]), .ZN(MCInst2_MC3_r0Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst2_MC3_r0Inst_XORInst_0_2_U1  ( .A(MCInst2_MC3_v0_0 [2]), .B(
        Red_MCInst2_MC3_v1_1[0] ), .Z(MCInst2_MC3_r0Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst2_MC3_r0Inst_XORInst_0_3_U3  ( .A(
        MCInst2_MC3_r0Inst_XORInst_0_3_n5 ), .B(
        MCInst2_MC3_r0Inst_XORInst_0_3_n4 ), .ZN(Feedback2[51]) );
  XNOR2_X1 MCInst2_MC3_r0Inst_XORInst_0_3_U2  ( .A(Red_MCInst2_MC3_v3_1[0] ), 
        .B(MCInst2_MC3_v2_0 [3]), .ZN(MCInst2_MC3_r0Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst2_MC3_r0Inst_XORInst_0_3_U1  ( .A(MCInst2_MC3_v0_0 [3]), .B(
        MCInst2_MC3_v1_0 [3]), .Z(MCInst2_MC3_r0Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst2_MC3_r1Inst_XORInst_0_0_U3  ( .A(
        MCInst2_MC3_r1Inst_XORInst_0_0_n5 ), .B(
        MCInst2_MC3_r1Inst_XORInst_0_0_n4 ), .ZN(Feedback2[32]) );
  XNOR2_X1 MCInst2_MC3_r1Inst_XORInst_0_0_U2  ( .A(MCInst2_MC3_v3_1 [0]), 
        .B(MCInst2_MC3_v2_1 [0]), .ZN(MCInst2_MC3_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst2_MC3_r1Inst_XORInst_0_0_U1  ( .A(MCInst2_MC3_v0_0 [3]), .B(
        MCInst2_MC3_v1_1 [0]), .Z(MCInst2_MC3_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst2_MC3_r1Inst_XORInst_0_1_U3  ( .A(
        MCInst2_MC3_r1Inst_XORInst_0_1_n5 ), .B(
        MCInst2_MC3_r1Inst_XORInst_0_1_n4 ), .ZN(Feedback2[33]) );
  XNOR2_X1 MCInst2_MC3_r1Inst_XORInst_0_1_U2  ( .A(MCInst2_MC3_v3_1 [1]), 
        .B(MCInst2_MC3_v2_1 [1]), .ZN(MCInst2_MC3_r1Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst2_MC3_r1Inst_XORInst_0_1_U1  ( .A(MCInst2_MC3_v0_1 [1]), .B(
        MCInst2_MC3_v1_1 [1]), .Z(MCInst2_MC3_r1Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst2_MC3_r1Inst_XORInst_0_2_U3  ( .A(
        MCInst2_MC3_r1Inst_XORInst_0_2_n5 ), .B(
        MCInst2_MC3_r1Inst_XORInst_0_2_n4 ), .ZN(Feedback2[34]) );
  XNOR2_X1 MCInst2_MC3_r1Inst_XORInst_0_2_U2  ( .A(MCInst2_MC3_v3_1 [2]), 
        .B(MCInst2_MC3_v2_1 [2]), .ZN(MCInst2_MC3_r1Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst2_MC3_r1Inst_XORInst_0_2_U1  ( .A(MCInst2_MC3_v0_1 [2]), .B(
        MCInst2_MC3_v1_1 [2]), .Z(MCInst2_MC3_r1Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst2_MC3_r1Inst_XORInst_0_3_U3  ( .A(
        MCInst2_MC3_r1Inst_XORInst_0_3_n5 ), .B(
        MCInst2_MC3_r1Inst_XORInst_0_3_n4 ), .ZN(Feedback2[35]) );
  XNOR2_X1 MCInst2_MC3_r1Inst_XORInst_0_3_U2  ( .A(MCInst2_MC3_v3_1 [3]), 
        .B(MCInst2_MC3_v2_1 [3]), .ZN(MCInst2_MC3_r1Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst2_MC3_r1Inst_XORInst_0_3_U1  ( .A(MCInst2_MC3_v0_1 [3]), .B(
        MCInst2_MC3_v1_1 [3]), .Z(MCInst2_MC3_r1Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst2_MC3_r2Inst_XORInst_0_0_U3  ( .A(
        MCInst2_MC3_r2Inst_XORInst_0_0_n5 ), .B(
        MCInst2_MC3_r2Inst_XORInst_0_0_n4 ), .ZN(Feedback2[16]) );
  XNOR2_X1 MCInst2_MC3_r2Inst_XORInst_0_0_U2  ( .A(MCInst2_MC3_v3_2 [0]), 
        .B(MCInst2_MC3_v2_2 [0]), .ZN(MCInst2_MC3_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst2_MC3_r2Inst_XORInst_0_0_U1  ( .A(MCInst2_MC3_v0_2 [0]), .B(
        MCInst2_MC3_v1_2 [0]), .Z(MCInst2_MC3_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst2_MC3_r2Inst_XORInst_0_1_U3  ( .A(
        MCInst2_MC3_r2Inst_XORInst_0_1_n5 ), .B(
        MCInst2_MC3_r2Inst_XORInst_0_1_n4 ), .ZN(Feedback2[17]) );
  XNOR2_X1 MCInst2_MC3_r2Inst_XORInst_0_1_U2  ( .A(Red_MCInst2_MC3_v3_1[0] ), 
        .B(MCInst2_MC3_v2_2 [1]), .ZN(MCInst2_MC3_r2Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst2_MC3_r2Inst_XORInst_0_1_U1  ( .A(MCInst2_MC3_v0_2 [1]), .B(
        MCInst2_MC3_v1_2 [1]), .Z(MCInst2_MC3_r2Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst2_MC3_r2Inst_XORInst_0_2_U3  ( .A(
        MCInst2_MC3_r2Inst_XORInst_0_2_n5 ), .B(
        MCInst2_MC3_r2Inst_XORInst_0_2_n4 ), .ZN(Feedback2[18]) );
  XNOR2_X1 MCInst2_MC3_r2Inst_XORInst_0_2_U2  ( .A(MCInst2_MC3_v3_2 [2]), 
        .B(MCInst2_MC3_v2_2 [2]), .ZN(MCInst2_MC3_r2Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst2_MC3_r2Inst_XORInst_0_2_U1  ( .A(MCInst2_MC3_v0_2 [2]), .B(
        MCInst2_MC3_v1_2 [2]), .Z(MCInst2_MC3_r2Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst2_MC3_r2Inst_XORInst_0_3_U3  ( .A(
        MCInst2_MC3_r2Inst_XORInst_0_3_n5 ), .B(
        MCInst2_MC3_r2Inst_XORInst_0_3_n4 ), .ZN(Feedback2[19]) );
  XNOR2_X1 MCInst2_MC3_r2Inst_XORInst_0_3_U2  ( .A(MCInst2_MC3_v3_2 [3]), 
        .B(MCInst2_MC3_v2_2 [3]), .ZN(MCInst2_MC3_r2Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst2_MC3_r2Inst_XORInst_0_3_U1  ( .A(MCInst2_MC3_v0_2 [3]), .B(
        MCInst2_MC3_v1_2 [3]), .Z(MCInst2_MC3_r2Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst2_MC3_r3Inst_XORInst_0_0_U3  ( .A(
        MCInst2_MC3_r3Inst_XORInst_0_0_n5 ), .B(
        MCInst2_MC3_r3Inst_XORInst_0_0_n4 ), .ZN(Feedback2[0]) );
  XNOR2_X1 MCInst2_MC3_r3Inst_XORInst_0_0_U2  ( .A(MCInst2_MC3_v3_3 [0]), 
        .B(MCInst2_MC3_v2_3 [0]), .ZN(MCInst2_MC3_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst2_MC3_r3Inst_XORInst_0_0_U1  ( .A(MCInst2_MC3_v0_3 [0]), .B(
        MCInst2_MC3_v1_0 [3]), .Z(MCInst2_MC3_r3Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst2_MC3_r3Inst_XORInst_0_1_U3  ( .A(
        MCInst2_MC3_r3Inst_XORInst_0_1_n5 ), .B(
        MCInst2_MC3_r3Inst_XORInst_0_1_n4 ), .ZN(Feedback2[1]) );
  XNOR2_X1 MCInst2_MC3_r3Inst_XORInst_0_1_U2  ( .A(MCInst2_MC3_v3_3 [1]), 
        .B(MCInst2_MC3_v2_3 [1]), .ZN(MCInst2_MC3_r3Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst2_MC3_r3Inst_XORInst_0_1_U1  ( .A(MCInst2_MC3_v0_3 [1]), .B(
        MCInst2_MC3_v1_3 [1]), .Z(MCInst2_MC3_r3Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst2_MC3_r3Inst_XORInst_0_2_U3  ( .A(
        MCInst2_MC3_r3Inst_XORInst_0_2_n5 ), .B(
        MCInst2_MC3_r3Inst_XORInst_0_2_n4 ), .ZN(Feedback2[2]) );
  XNOR2_X1 MCInst2_MC3_r3Inst_XORInst_0_2_U2  ( .A(MCInst2_MC3_v3_3 [2]), 
        .B(MCInst2_MC3_v2_3 [2]), .ZN(MCInst2_MC3_r3Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst2_MC3_r3Inst_XORInst_0_2_U1  ( .A(MCInst2_MC3_v0_0 [3]), .B(
        MCInst2_MC3_v1_3 [2]), .Z(MCInst2_MC3_r3Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst2_MC3_r3Inst_XORInst_0_3_U3  ( .A(
        MCInst2_MC3_r3Inst_XORInst_0_3_n5 ), .B(
        MCInst2_MC3_r3Inst_XORInst_0_3_n4 ), .ZN(Feedback2[3]) );
  XNOR2_X1 MCInst2_MC3_r3Inst_XORInst_0_3_U2  ( .A(MCInst2_MC3_v3_3 [3]), 
        .B(MCInst2_MC3_v2_3 [3]), .ZN(MCInst2_MC3_r3Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst2_MC3_r3Inst_XORInst_0_3_U1  ( .A(MCInst2_MC3_v0_3 [3]), .B(
        Red_MCInst2_MC3_v1_1[0] ), .Z(MCInst2_MC3_r3Inst_XORInst_0_3_n5 ) );
  DFF_X1 StateReg2_s_current_state_reg[0]  ( .D(Feedback2[0]), .CK(clk), .Q(
        SubCellInput2[0]) );
  DFF_X1 StateReg2_s_current_state_reg[1]  ( .D(Feedback2[1]), .CK(clk), .Q(
        SubCellInput2[1]) );
  DFF_X1 StateReg2_s_current_state_reg[2]  ( .D(Feedback2[2]), .CK(clk), .Q(
        SubCellInput2[2]) );
  DFF_X1 StateReg2_s_current_state_reg[3]  ( .D(Feedback2[3]), .CK(clk), .Q(
        SubCellInput2[3]) );
  DFF_X1 StateReg2_s_current_state_reg[4]  ( .D(Feedback2[4]), .CK(clk), .Q(
        SubCellInput2[4]) );
  DFF_X1 StateReg2_s_current_state_reg[5]  ( .D(Feedback2[5]), .CK(clk), .Q(
        SubCellInput2[5]) );
  DFF_X1 StateReg2_s_current_state_reg[6]  ( .D(Feedback2[6]), .CK(clk), .Q(
        SubCellInput2[6]) );
  DFF_X1 StateReg2_s_current_state_reg[7]  ( .D(Feedback2[7]), .CK(clk), .Q(
        SubCellInput2[7]) );
  DFF_X1 StateReg2_s_current_state_reg[8]  ( .D(Feedback2[8]), .CK(clk), .Q(
        SubCellInput2[8]) );
  DFF_X1 StateReg2_s_current_state_reg[9]  ( .D(Feedback2[9]), .CK(clk), .Q(
        SubCellInput2[9]) );
  DFF_X1 StateReg2_s_current_state_reg[10]  ( .D(Feedback2[10]), .CK(clk), 
        .Q(SubCellInput2[10]) );
  DFF_X1 StateReg2_s_current_state_reg[11]  ( .D(Feedback2[11]), .CK(clk), 
        .Q(SubCellInput2[11]) );
  DFF_X1 StateReg2_s_current_state_reg[12]  ( .D(Feedback2[12]), .CK(clk), 
        .Q(SubCellInput2[12]) );
  DFF_X1 StateReg2_s_current_state_reg[13]  ( .D(Feedback2[13]), .CK(clk), 
        .Q(SubCellInput2[13]) );
  DFF_X1 StateReg2_s_current_state_reg[14]  ( .D(Feedback2[14]), .CK(clk), 
        .Q(SubCellInput2[14]) );
  DFF_X1 StateReg2_s_current_state_reg[15]  ( .D(Feedback2[15]), .CK(clk), 
        .Q(SubCellInput2[15]) );
  DFF_X1 StateReg2_s_current_state_reg[16]  ( .D(Feedback2[16]), .CK(clk), 
        .Q(SubCellInput2[16]) );
  DFF_X1 StateReg2_s_current_state_reg[17]  ( .D(Feedback2[17]), .CK(clk), 
        .Q(SubCellInput2[17]) );
  DFF_X1 StateReg2_s_current_state_reg[18]  ( .D(Feedback2[18]), .CK(clk), 
        .Q(SubCellInput2[18]) );
  DFF_X1 StateReg2_s_current_state_reg[19]  ( .D(Feedback2[19]), .CK(clk), 
        .Q(SubCellInput2[19]) );
  DFF_X1 StateReg2_s_current_state_reg[20]  ( .D(Feedback2[20]), .CK(clk), 
        .Q(SubCellInput2[20]) );
  DFF_X1 StateReg2_s_current_state_reg[21]  ( .D(Feedback2[21]), .CK(clk), 
        .Q(SubCellInput2[21]) );
  DFF_X1 StateReg2_s_current_state_reg[22]  ( .D(Feedback2[22]), .CK(clk), 
        .Q(SubCellInput2[22]) );
  DFF_X1 StateReg2_s_current_state_reg[23]  ( .D(Feedback2[23]), .CK(clk), 
        .Q(SubCellInput2[23]) );
  DFF_X1 StateReg2_s_current_state_reg[24]  ( .D(Feedback2[24]), .CK(clk), 
        .Q(SubCellInput2[24]) );
  DFF_X1 StateReg2_s_current_state_reg[25]  ( .D(Feedback2[25]), .CK(clk), 
        .Q(SubCellInput2[25]) );
  DFF_X1 StateReg2_s_current_state_reg[26]  ( .D(Feedback2[26]), .CK(clk), 
        .Q(SubCellInput2[26]) );
  DFF_X1 StateReg2_s_current_state_reg[27]  ( .D(Feedback2[27]), .CK(clk), 
        .Q(SubCellInput2[27]) );
  DFF_X1 StateReg2_s_current_state_reg[28]  ( .D(Feedback2[28]), .CK(clk), 
        .Q(SubCellInput2[28]) );
  DFF_X1 StateReg2_s_current_state_reg[29]  ( .D(Feedback2[29]), .CK(clk), 
        .Q(SubCellInput2[29]) );
  DFF_X1 StateReg2_s_current_state_reg[30]  ( .D(Feedback2[30]), .CK(clk), 
        .Q(SubCellInput2[30]) );
  DFF_X1 StateReg2_s_current_state_reg[31]  ( .D(Feedback2[31]), .CK(clk), 
        .Q(SubCellInput2[31]) );
  DFF_X1 StateReg2_s_current_state_reg[32]  ( .D(Feedback2[32]), .CK(clk), 
        .Q(SubCellInput2[32]) );
  DFF_X1 StateReg2_s_current_state_reg[33]  ( .D(Feedback2[33]), .CK(clk), 
        .Q(SubCellInput2[33]) );
  DFF_X1 StateReg2_s_current_state_reg[34]  ( .D(Feedback2[34]), .CK(clk), 
        .Q(SubCellInput2[34]) );
  DFF_X1 StateReg2_s_current_state_reg[35]  ( .D(Feedback2[35]), .CK(clk), 
        .Q(SubCellInput2[35]) );
  DFF_X1 StateReg2_s_current_state_reg[36]  ( .D(Feedback2[36]), .CK(clk), 
        .Q(SubCellInput2[36]) );
  DFF_X1 StateReg2_s_current_state_reg[37]  ( .D(Feedback2[37]), .CK(clk), 
        .Q(SubCellInput2[37]) );
  DFF_X1 StateReg2_s_current_state_reg[38]  ( .D(Feedback2[38]), .CK(clk), 
        .Q(SubCellInput2[38]) );
  DFF_X1 StateReg2_s_current_state_reg[39]  ( .D(Feedback2[39]), .CK(clk), 
        .Q(SubCellInput2[39]) );
  DFF_X1 StateReg2_s_current_state_reg[40]  ( .D(Feedback2[40]), .CK(clk), 
        .Q(SubCellInput2[40]) );
  DFF_X1 StateReg2_s_current_state_reg[41]  ( .D(Feedback2[41]), .CK(clk), 
        .Q(SubCellInput2[41]) );
  DFF_X1 StateReg2_s_current_state_reg[42]  ( .D(Feedback2[42]), .CK(clk), 
        .Q(SubCellInput2[42]) );
  DFF_X1 StateReg2_s_current_state_reg[43]  ( .D(Feedback2[43]), .CK(clk), 
        .Q(SubCellInput2[43]) );
  DFF_X1 StateReg2_s_current_state_reg[44]  ( .D(Feedback2[44]), .CK(clk), 
        .Q(SubCellInput2[44]) );
  DFF_X1 StateReg2_s_current_state_reg[45]  ( .D(Feedback2[45]), .CK(clk), 
        .Q(SubCellInput2[45]) );
  DFF_X1 StateReg2_s_current_state_reg[46]  ( .D(Feedback2[46]), .CK(clk), 
        .Q(SubCellInput2[46]) );
  DFF_X1 StateReg2_s_current_state_reg[47]  ( .D(Feedback2[47]), .CK(clk), 
        .Q(SubCellInput2[47]) );
  DFF_X1 StateReg2_s_current_state_reg[48]  ( .D(Feedback2[48]), .CK(clk), 
        .Q(SubCellInput2[48]) );
  DFF_X1 StateReg2_s_current_state_reg[49]  ( .D(Feedback2[49]), .CK(clk), 
        .Q(SubCellInput2[49]) );
  DFF_X1 StateReg2_s_current_state_reg[50]  ( .D(Feedback2[50]), .CK(clk), 
        .Q(SubCellInput2[50]) );
  DFF_X1 StateReg2_s_current_state_reg[51]  ( .D(Feedback2[51]), .CK(clk), 
        .Q(SubCellInput2[51]) );
  DFF_X1 StateReg2_s_current_state_reg[52]  ( .D(Feedback2[52]), .CK(clk), 
        .Q(SubCellInput2[52]) );
  DFF_X1 StateReg2_s_current_state_reg[53]  ( .D(Feedback2[53]), .CK(clk), 
        .Q(SubCellInput2[53]) );
  DFF_X1 StateReg2_s_current_state_reg[54]  ( .D(Feedback2[54]), .CK(clk), 
        .Q(SubCellInput2[54]) );
  DFF_X1 StateReg2_s_current_state_reg[55]  ( .D(Feedback2[55]), .CK(clk), 
        .Q(SubCellInput2[55]) );
  DFF_X1 StateReg2_s_current_state_reg[56]  ( .D(Feedback2[56]), .CK(clk), 
        .Q(SubCellInput2[56]) );
  DFF_X1 StateReg2_s_current_state_reg[57]  ( .D(Feedback2[57]), .CK(clk), 
        .Q(SubCellInput2[57]) );
  DFF_X1 StateReg2_s_current_state_reg[58]  ( .D(Feedback2[58]), .CK(clk), 
        .Q(SubCellInput2[58]) );
  DFF_X1 StateReg2_s_current_state_reg[59]  ( .D(Feedback2[59]), .CK(clk), 
        .Q(SubCellInput2[59]) );
  DFF_X1 StateReg2_s_current_state_reg[60]  ( .D(Feedback2[60]), .CK(clk), 
        .Q(SubCellInput2[60]) );
  DFF_X1 StateReg2_s_current_state_reg[61]  ( .D(Feedback2[61]), .CK(clk), 
        .Q(SubCellInput2[61]) );
  DFF_X1 StateReg2_s_current_state_reg[62]  ( .D(Feedback2[62]), .CK(clk), 
        .Q(SubCellInput2[62]) );
  DFF_X1 StateReg2_s_current_state_reg[63]  ( .D(Feedback2[63]), .CK(clk), 
        .Q(SubCellInput2[63]) );
  NAND2_X1 SubCellInst3_LFInst_0_LFInst_0_U6  ( .A1(SubCellInput2[2]), .A2(
        SubCellInst3_LFInst_0_LFInst_0_n4 ), .ZN(
        SubCellInst3_LFInst_0_LFInst_0_n5 ) );
  INV_X1 SubCellInst3_LFInst_0_LFInst_0_U5  ( .A(SubCellInput2[1]), .ZN(
        SubCellInst3_LFInst_0_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst3_LFInst_0_LFInst_0_U4  ( .A(SubCellInput2[0]), .B(
        SubCellInput2[3]), .Z(SubCellInst3_LFInst_0_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst3_LFInst_0_LFInst_0_U3  ( .A(
        SubCellInst3_LFInst_0_LFInst_0_n6 ), .B(
        SubCellInst3_LFInst_0_LFInst_0_n5 ), .ZN(MCInst3_MC0_v3_2 [3]) );
  NAND2_X1 SubCellInst3_LFInst_0_LFInst_1_U12  ( .A1(
        SubCellInst3_LFInst_0_LFInst_1_n18 ), .A2(
        SubCellInst3_LFInst_0_LFInst_1_n17 ), .ZN(MCInst3_MC0_v3_0 [2]) );
  NAND2_X1 SubCellInst3_LFInst_0_LFInst_1_U11  ( .A1(SubCellInput2[1]), .A2(
        SubCellInst3_LFInst_0_LFInst_1_n16 ), .ZN(
        SubCellInst3_LFInst_0_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst3_LFInst_0_LFInst_1_U10  ( .A1(SubCellInput2[3]), .A2(
        SubCellInst3_LFInst_0_LFInst_1_n15 ), .ZN(
        SubCellInst3_LFInst_0_LFInst_1_n16 ) );
  AND2_X1 SubCellInst3_LFInst_0_LFInst_1_U9  ( .A1(SubCellInput2[0]), .A2(
        SubCellInput2[2]), .ZN(SubCellInst3_LFInst_0_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst3_LFInst_0_LFInst_1_U8  ( .A1(SubCellInput2[3]), .A2(
        SubCellInst3_LFInst_0_LFInst_1_n14 ), .ZN(
        SubCellInst3_LFInst_0_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst3_LFInst_0_LFInst_1_U7  ( .A1(
        SubCellInst3_LFInst_0_LFInst_1_n13 ), .A2(
        SubCellInst3_LFInst_0_LFInst_1_n12 ), .ZN(
        SubCellInst3_LFInst_0_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst3_LFInst_0_LFInst_1_U6  ( .A1(SubCellInput2[0]), .A2(
        SubCellInput2[2]), .ZN(SubCellInst3_LFInst_0_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst3_LFInst_0_LFInst_1_U5  ( .A1(
        SubCellInst3_LFInst_0_LFInst_1_n11 ), .A2(
        SubCellInst3_LFInst_0_LFInst_1_n10 ), .ZN(
        SubCellInst3_LFInst_0_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst3_LFInst_0_LFInst_1_U4  ( .A1(SubCellInput2[0]), .A2(
        SubCellInput2[1]), .ZN(SubCellInst3_LFInst_0_LFInst_1_n10 ) );
  INV_X1 SubCellInst3_LFInst_0_LFInst_1_U3  ( .A(SubCellInput2[2]), .ZN(
        SubCellInst3_LFInst_0_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst3_LFInst_0_LFInst_2_U11  ( .A1(
        SubCellInst3_LFInst_0_LFInst_2_n22 ), .A2(
        SubCellInst3_LFInst_0_LFInst_2_n21 ), .ZN(Red_MCInst3_MC0_v3_1[0] )
         );
  NAND2_X1 SubCellInst3_LFInst_0_LFInst_2_U10  ( .A1(SubCellInput2[2]), .A2(
        SubCellInst3_LFInst_0_LFInst_2_n20 ), .ZN(
        SubCellInst3_LFInst_0_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst3_LFInst_0_LFInst_2_U9  ( .A1(SubCellInput2[1]), .A2(
        SubCellInst3_LFInst_0_LFInst_2_n19 ), .ZN(
        SubCellInst3_LFInst_0_LFInst_2_n20 ) );
  INV_X1 SubCellInst3_LFInst_0_LFInst_2_U8  ( .A(SubCellInput2[3]), .ZN(
        SubCellInst3_LFInst_0_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst3_LFInst_0_LFInst_2_U7  ( .A1(
        SubCellInst3_LFInst_0_LFInst_2_n18 ), .A2(
        SubCellInst3_LFInst_0_LFInst_2_n17 ), .ZN(
        SubCellInst3_LFInst_0_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst3_LFInst_0_LFInst_2_U6  ( .A(
        SubCellInst3_LFInst_0_LFInst_2_n16 ), .B(SubCellInput2[2]), .Z(
        SubCellInst3_LFInst_0_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst3_LFInst_0_LFInst_2_U5  ( .A1(SubCellInput2[0]), .A2(
        SubCellInput2[1]), .ZN(SubCellInst3_LFInst_0_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst3_LFInst_0_LFInst_2_U4  ( .A1(
        SubCellInst3_LFInst_0_LFInst_2_n15 ), .A2(SubCellInput2[3]), .ZN(
        SubCellInst3_LFInst_0_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst3_LFInst_0_LFInst_2_U3  ( .A(SubCellInput2[0]), .B(
        SubCellInput2[1]), .ZN(SubCellInst3_LFInst_0_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst3_LFInst_0_LFInst_3_U9  ( .A1(
        SubCellInst3_LFInst_0_LFInst_3_n16 ), .A2(
        SubCellInst3_LFInst_0_LFInst_3_n15 ), .ZN(MCInst3_MC0_v3_2 [2]) );
  NAND2_X1 SubCellInst3_LFInst_0_LFInst_3_U8  ( .A1(SubCellInput2[1]), .A2(
        SubCellInst3_LFInst_0_LFInst_3_n14 ), .ZN(
        SubCellInst3_LFInst_0_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst3_LFInst_0_LFInst_3_U7  ( .A(SubCellInput2[3]), .B(
        SubCellInput2[2]), .Z(SubCellInst3_LFInst_0_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst3_LFInst_0_LFInst_3_U6  ( .A1(
        SubCellInst3_LFInst_0_LFInst_3_n13 ), .A2(
        SubCellInst3_LFInst_0_LFInst_3_n12 ), .ZN(
        SubCellInst3_LFInst_0_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst3_LFInst_0_LFInst_3_U5  ( .A1(SubCellInput2[0]), .A2(
        SubCellInput2[2]), .ZN(SubCellInst3_LFInst_0_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst3_LFInst_0_LFInst_3_U4  ( .A(SubCellInput2[0]), .B(
        SubCellInst3_LFInst_0_LFInst_3_n11 ), .ZN(
        SubCellInst3_LFInst_0_LFInst_3_n13 ) );
  OR2_X1 SubCellInst3_LFInst_0_LFInst_3_U3  ( .A1(SubCellInput2[3]), .A2(
        SubCellInput2[1]), .ZN(SubCellInst3_LFInst_0_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst3_LFInst_1_LFInst_0_U6  ( .A1(SubCellInput2[6]), .A2(
        SubCellInst3_LFInst_1_LFInst_0_n4 ), .ZN(
        SubCellInst3_LFInst_1_LFInst_0_n5 ) );
  INV_X1 SubCellInst3_LFInst_1_LFInst_0_U5  ( .A(SubCellInput2[5]), .ZN(
        SubCellInst3_LFInst_1_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst3_LFInst_1_LFInst_0_U4  ( .A(SubCellInput2[4]), .B(
        SubCellInput2[7]), .Z(SubCellInst3_LFInst_1_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst3_LFInst_1_LFInst_0_U3  ( .A(
        SubCellInst3_LFInst_1_LFInst_0_n6 ), .B(
        SubCellInst3_LFInst_1_LFInst_0_n5 ), .ZN(MCInst3_MC3_v3_2 [3]) );
  NAND2_X1 SubCellInst3_LFInst_1_LFInst_1_U12  ( .A1(
        SubCellInst3_LFInst_1_LFInst_1_n18 ), .A2(
        SubCellInst3_LFInst_1_LFInst_1_n17 ), .ZN(MCInst3_MC3_v3_0 [2]) );
  NAND2_X1 SubCellInst3_LFInst_1_LFInst_1_U11  ( .A1(SubCellInput2[5]), .A2(
        SubCellInst3_LFInst_1_LFInst_1_n16 ), .ZN(
        SubCellInst3_LFInst_1_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst3_LFInst_1_LFInst_1_U10  ( .A1(SubCellInput2[7]), .A2(
        SubCellInst3_LFInst_1_LFInst_1_n15 ), .ZN(
        SubCellInst3_LFInst_1_LFInst_1_n16 ) );
  AND2_X1 SubCellInst3_LFInst_1_LFInst_1_U9  ( .A1(SubCellInput2[4]), .A2(
        SubCellInput2[6]), .ZN(SubCellInst3_LFInst_1_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst3_LFInst_1_LFInst_1_U8  ( .A1(SubCellInput2[7]), .A2(
        SubCellInst3_LFInst_1_LFInst_1_n14 ), .ZN(
        SubCellInst3_LFInst_1_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst3_LFInst_1_LFInst_1_U7  ( .A1(
        SubCellInst3_LFInst_1_LFInst_1_n13 ), .A2(
        SubCellInst3_LFInst_1_LFInst_1_n12 ), .ZN(
        SubCellInst3_LFInst_1_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst3_LFInst_1_LFInst_1_U6  ( .A1(SubCellInput2[4]), .A2(
        SubCellInput2[6]), .ZN(SubCellInst3_LFInst_1_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst3_LFInst_1_LFInst_1_U5  ( .A1(
        SubCellInst3_LFInst_1_LFInst_1_n11 ), .A2(
        SubCellInst3_LFInst_1_LFInst_1_n10 ), .ZN(
        SubCellInst3_LFInst_1_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst3_LFInst_1_LFInst_1_U4  ( .A1(SubCellInput2[4]), .A2(
        SubCellInput2[5]), .ZN(SubCellInst3_LFInst_1_LFInst_1_n10 ) );
  INV_X1 SubCellInst3_LFInst_1_LFInst_1_U3  ( .A(SubCellInput2[6]), .ZN(
        SubCellInst3_LFInst_1_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst3_LFInst_1_LFInst_2_U11  ( .A1(
        SubCellInst3_LFInst_1_LFInst_2_n22 ), .A2(
        SubCellInst3_LFInst_1_LFInst_2_n21 ), .ZN(Red_MCInst3_MC3_v3_1[0] )
         );
  NAND2_X1 SubCellInst3_LFInst_1_LFInst_2_U10  ( .A1(SubCellInput2[6]), .A2(
        SubCellInst3_LFInst_1_LFInst_2_n20 ), .ZN(
        SubCellInst3_LFInst_1_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst3_LFInst_1_LFInst_2_U9  ( .A1(SubCellInput2[5]), .A2(
        SubCellInst3_LFInst_1_LFInst_2_n19 ), .ZN(
        SubCellInst3_LFInst_1_LFInst_2_n20 ) );
  INV_X1 SubCellInst3_LFInst_1_LFInst_2_U8  ( .A(SubCellInput2[7]), .ZN(
        SubCellInst3_LFInst_1_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst3_LFInst_1_LFInst_2_U7  ( .A1(
        SubCellInst3_LFInst_1_LFInst_2_n18 ), .A2(
        SubCellInst3_LFInst_1_LFInst_2_n17 ), .ZN(
        SubCellInst3_LFInst_1_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst3_LFInst_1_LFInst_2_U6  ( .A(
        SubCellInst3_LFInst_1_LFInst_2_n16 ), .B(SubCellInput2[6]), .Z(
        SubCellInst3_LFInst_1_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst3_LFInst_1_LFInst_2_U5  ( .A1(SubCellInput2[4]), .A2(
        SubCellInput2[5]), .ZN(SubCellInst3_LFInst_1_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst3_LFInst_1_LFInst_2_U4  ( .A1(
        SubCellInst3_LFInst_1_LFInst_2_n15 ), .A2(SubCellInput2[7]), .ZN(
        SubCellInst3_LFInst_1_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst3_LFInst_1_LFInst_2_U3  ( .A(SubCellInput2[4]), .B(
        SubCellInput2[5]), .ZN(SubCellInst3_LFInst_1_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst3_LFInst_1_LFInst_3_U9  ( .A1(
        SubCellInst3_LFInst_1_LFInst_3_n16 ), .A2(
        SubCellInst3_LFInst_1_LFInst_3_n15 ), .ZN(MCInst3_MC3_v3_2 [2]) );
  NAND2_X1 SubCellInst3_LFInst_1_LFInst_3_U8  ( .A1(SubCellInput2[5]), .A2(
        SubCellInst3_LFInst_1_LFInst_3_n14 ), .ZN(
        SubCellInst3_LFInst_1_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst3_LFInst_1_LFInst_3_U7  ( .A(SubCellInput2[7]), .B(
        SubCellInput2[6]), .Z(SubCellInst3_LFInst_1_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst3_LFInst_1_LFInst_3_U6  ( .A1(
        SubCellInst3_LFInst_1_LFInst_3_n13 ), .A2(
        SubCellInst3_LFInst_1_LFInst_3_n12 ), .ZN(
        SubCellInst3_LFInst_1_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst3_LFInst_1_LFInst_3_U5  ( .A1(SubCellInput2[4]), .A2(
        SubCellInput2[6]), .ZN(SubCellInst3_LFInst_1_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst3_LFInst_1_LFInst_3_U4  ( .A(SubCellInput2[4]), .B(
        SubCellInst3_LFInst_1_LFInst_3_n11 ), .ZN(
        SubCellInst3_LFInst_1_LFInst_3_n13 ) );
  OR2_X1 SubCellInst3_LFInst_1_LFInst_3_U3  ( .A1(SubCellInput2[7]), .A2(
        SubCellInput2[5]), .ZN(SubCellInst3_LFInst_1_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst3_LFInst_2_LFInst_0_U6  ( .A1(SubCellInput2[10]), .A2(
        SubCellInst3_LFInst_2_LFInst_0_n4 ), .ZN(
        SubCellInst3_LFInst_2_LFInst_0_n5 ) );
  INV_X1 SubCellInst3_LFInst_2_LFInst_0_U5  ( .A(SubCellInput2[9]), .ZN(
        SubCellInst3_LFInst_2_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst3_LFInst_2_LFInst_0_U4  ( .A(SubCellInput2[8]), .B(
        SubCellInput2[11]), .Z(SubCellInst3_LFInst_2_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst3_LFInst_2_LFInst_0_U3  ( .A(
        SubCellInst3_LFInst_2_LFInst_0_n6 ), .B(
        SubCellInst3_LFInst_2_LFInst_0_n5 ), .ZN(MCInst3_MC2_v3_2 [3]) );
  NAND2_X1 SubCellInst3_LFInst_2_LFInst_1_U12  ( .A1(
        SubCellInst3_LFInst_2_LFInst_1_n18 ), .A2(
        SubCellInst3_LFInst_2_LFInst_1_n17 ), .ZN(MCInst3_MC2_v3_0 [2]) );
  NAND2_X1 SubCellInst3_LFInst_2_LFInst_1_U11  ( .A1(SubCellInput2[9]), .A2(
        SubCellInst3_LFInst_2_LFInst_1_n16 ), .ZN(
        SubCellInst3_LFInst_2_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst3_LFInst_2_LFInst_1_U10  ( .A1(SubCellInput2[11]), .A2(
        SubCellInst3_LFInst_2_LFInst_1_n15 ), .ZN(
        SubCellInst3_LFInst_2_LFInst_1_n16 ) );
  AND2_X1 SubCellInst3_LFInst_2_LFInst_1_U9  ( .A1(SubCellInput2[8]), .A2(
        SubCellInput2[10]), .ZN(SubCellInst3_LFInst_2_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst3_LFInst_2_LFInst_1_U8  ( .A1(SubCellInput2[11]), .A2(
        SubCellInst3_LFInst_2_LFInst_1_n14 ), .ZN(
        SubCellInst3_LFInst_2_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst3_LFInst_2_LFInst_1_U7  ( .A1(
        SubCellInst3_LFInst_2_LFInst_1_n13 ), .A2(
        SubCellInst3_LFInst_2_LFInst_1_n12 ), .ZN(
        SubCellInst3_LFInst_2_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst3_LFInst_2_LFInst_1_U6  ( .A1(SubCellInput2[8]), .A2(
        SubCellInput2[10]), .ZN(SubCellInst3_LFInst_2_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst3_LFInst_2_LFInst_1_U5  ( .A1(
        SubCellInst3_LFInst_2_LFInst_1_n11 ), .A2(
        SubCellInst3_LFInst_2_LFInst_1_n10 ), .ZN(
        SubCellInst3_LFInst_2_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst3_LFInst_2_LFInst_1_U4  ( .A1(SubCellInput2[8]), .A2(
        SubCellInput2[9]), .ZN(SubCellInst3_LFInst_2_LFInst_1_n10 ) );
  INV_X1 SubCellInst3_LFInst_2_LFInst_1_U3  ( .A(SubCellInput2[10]), .ZN(
        SubCellInst3_LFInst_2_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst3_LFInst_2_LFInst_2_U11  ( .A1(
        SubCellInst3_LFInst_2_LFInst_2_n22 ), .A2(
        SubCellInst3_LFInst_2_LFInst_2_n21 ), .ZN(Red_MCInst3_MC2_v3_1[0] )
         );
  NAND2_X1 SubCellInst3_LFInst_2_LFInst_2_U10  ( .A1(SubCellInput2[10]), .A2(
        SubCellInst3_LFInst_2_LFInst_2_n20 ), .ZN(
        SubCellInst3_LFInst_2_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst3_LFInst_2_LFInst_2_U9  ( .A1(SubCellInput2[9]), .A2(
        SubCellInst3_LFInst_2_LFInst_2_n19 ), .ZN(
        SubCellInst3_LFInst_2_LFInst_2_n20 ) );
  INV_X1 SubCellInst3_LFInst_2_LFInst_2_U8  ( .A(SubCellInput2[11]), .ZN(
        SubCellInst3_LFInst_2_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst3_LFInst_2_LFInst_2_U7  ( .A1(
        SubCellInst3_LFInst_2_LFInst_2_n18 ), .A2(
        SubCellInst3_LFInst_2_LFInst_2_n17 ), .ZN(
        SubCellInst3_LFInst_2_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst3_LFInst_2_LFInst_2_U6  ( .A(
        SubCellInst3_LFInst_2_LFInst_2_n16 ), .B(SubCellInput2[10]), .Z(
        SubCellInst3_LFInst_2_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst3_LFInst_2_LFInst_2_U5  ( .A1(SubCellInput2[8]), .A2(
        SubCellInput2[9]), .ZN(SubCellInst3_LFInst_2_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst3_LFInst_2_LFInst_2_U4  ( .A1(
        SubCellInst3_LFInst_2_LFInst_2_n15 ), .A2(SubCellInput2[11]), .ZN(
        SubCellInst3_LFInst_2_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst3_LFInst_2_LFInst_2_U3  ( .A(SubCellInput2[8]), .B(
        SubCellInput2[9]), .ZN(SubCellInst3_LFInst_2_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst3_LFInst_2_LFInst_3_U9  ( .A1(
        SubCellInst3_LFInst_2_LFInst_3_n16 ), .A2(
        SubCellInst3_LFInst_2_LFInst_3_n15 ), .ZN(MCInst3_MC2_v3_2 [2]) );
  NAND2_X1 SubCellInst3_LFInst_2_LFInst_3_U8  ( .A1(SubCellInput2[9]), .A2(
        SubCellInst3_LFInst_2_LFInst_3_n14 ), .ZN(
        SubCellInst3_LFInst_2_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst3_LFInst_2_LFInst_3_U7  ( .A(SubCellInput2[11]), .B(
        SubCellInput2[10]), .Z(SubCellInst3_LFInst_2_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst3_LFInst_2_LFInst_3_U6  ( .A1(
        SubCellInst3_LFInst_2_LFInst_3_n13 ), .A2(
        SubCellInst3_LFInst_2_LFInst_3_n12 ), .ZN(
        SubCellInst3_LFInst_2_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst3_LFInst_2_LFInst_3_U5  ( .A1(SubCellInput2[8]), .A2(
        SubCellInput2[10]), .ZN(SubCellInst3_LFInst_2_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst3_LFInst_2_LFInst_3_U4  ( .A(SubCellInput2[8]), .B(
        SubCellInst3_LFInst_2_LFInst_3_n11 ), .ZN(
        SubCellInst3_LFInst_2_LFInst_3_n13 ) );
  OR2_X1 SubCellInst3_LFInst_2_LFInst_3_U3  ( .A1(SubCellInput2[11]), .A2(
        SubCellInput2[9]), .ZN(SubCellInst3_LFInst_2_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst3_LFInst_3_LFInst_0_U6  ( .A1(SubCellInput2[14]), .A2(
        SubCellInst3_LFInst_3_LFInst_0_n4 ), .ZN(
        SubCellInst3_LFInst_3_LFInst_0_n5 ) );
  INV_X1 SubCellInst3_LFInst_3_LFInst_0_U5  ( .A(SubCellInput2[13]), .ZN(
        SubCellInst3_LFInst_3_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst3_LFInst_3_LFInst_0_U4  ( .A(SubCellInput2[12]), .B(
        SubCellInput2[15]), .Z(SubCellInst3_LFInst_3_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst3_LFInst_3_LFInst_0_U3  ( .A(
        SubCellInst3_LFInst_3_LFInst_0_n6 ), .B(
        SubCellInst3_LFInst_3_LFInst_0_n5 ), .ZN(MCInst3_MC1_v3_2 [3]) );
  NAND2_X1 SubCellInst3_LFInst_3_LFInst_1_U12  ( .A1(
        SubCellInst3_LFInst_3_LFInst_1_n18 ), .A2(
        SubCellInst3_LFInst_3_LFInst_1_n17 ), .ZN(MCInst3_MC1_v3_0 [2]) );
  NAND2_X1 SubCellInst3_LFInst_3_LFInst_1_U11  ( .A1(SubCellInput2[13]), .A2(
        SubCellInst3_LFInst_3_LFInst_1_n16 ), .ZN(
        SubCellInst3_LFInst_3_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst3_LFInst_3_LFInst_1_U10  ( .A1(SubCellInput2[15]), .A2(
        SubCellInst3_LFInst_3_LFInst_1_n15 ), .ZN(
        SubCellInst3_LFInst_3_LFInst_1_n16 ) );
  AND2_X1 SubCellInst3_LFInst_3_LFInst_1_U9  ( .A1(SubCellInput2[12]), .A2(
        SubCellInput2[14]), .ZN(SubCellInst3_LFInst_3_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst3_LFInst_3_LFInst_1_U8  ( .A1(SubCellInput2[15]), .A2(
        SubCellInst3_LFInst_3_LFInst_1_n14 ), .ZN(
        SubCellInst3_LFInst_3_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst3_LFInst_3_LFInst_1_U7  ( .A1(
        SubCellInst3_LFInst_3_LFInst_1_n13 ), .A2(
        SubCellInst3_LFInst_3_LFInst_1_n12 ), .ZN(
        SubCellInst3_LFInst_3_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst3_LFInst_3_LFInst_1_U6  ( .A1(SubCellInput2[12]), .A2(
        SubCellInput2[14]), .ZN(SubCellInst3_LFInst_3_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst3_LFInst_3_LFInst_1_U5  ( .A1(
        SubCellInst3_LFInst_3_LFInst_1_n11 ), .A2(
        SubCellInst3_LFInst_3_LFInst_1_n10 ), .ZN(
        SubCellInst3_LFInst_3_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst3_LFInst_3_LFInst_1_U4  ( .A1(SubCellInput2[12]), .A2(
        SubCellInput2[13]), .ZN(SubCellInst3_LFInst_3_LFInst_1_n10 ) );
  INV_X1 SubCellInst3_LFInst_3_LFInst_1_U3  ( .A(SubCellInput2[14]), .ZN(
        SubCellInst3_LFInst_3_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst3_LFInst_3_LFInst_2_U11  ( .A1(
        SubCellInst3_LFInst_3_LFInst_2_n22 ), .A2(
        SubCellInst3_LFInst_3_LFInst_2_n21 ), .ZN(Red_MCInst3_MC1_v3_1[0] )
         );
  NAND2_X1 SubCellInst3_LFInst_3_LFInst_2_U10  ( .A1(SubCellInput2[14]), .A2(
        SubCellInst3_LFInst_3_LFInst_2_n20 ), .ZN(
        SubCellInst3_LFInst_3_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst3_LFInst_3_LFInst_2_U9  ( .A1(SubCellInput2[13]), .A2(
        SubCellInst3_LFInst_3_LFInst_2_n19 ), .ZN(
        SubCellInst3_LFInst_3_LFInst_2_n20 ) );
  INV_X1 SubCellInst3_LFInst_3_LFInst_2_U8  ( .A(SubCellInput2[15]), .ZN(
        SubCellInst3_LFInst_3_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst3_LFInst_3_LFInst_2_U7  ( .A1(
        SubCellInst3_LFInst_3_LFInst_2_n18 ), .A2(
        SubCellInst3_LFInst_3_LFInst_2_n17 ), .ZN(
        SubCellInst3_LFInst_3_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst3_LFInst_3_LFInst_2_U6  ( .A(
        SubCellInst3_LFInst_3_LFInst_2_n16 ), .B(SubCellInput2[14]), .Z(
        SubCellInst3_LFInst_3_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst3_LFInst_3_LFInst_2_U5  ( .A1(SubCellInput2[12]), .A2(
        SubCellInput2[13]), .ZN(SubCellInst3_LFInst_3_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst3_LFInst_3_LFInst_2_U4  ( .A1(
        SubCellInst3_LFInst_3_LFInst_2_n15 ), .A2(SubCellInput2[15]), .ZN(
        SubCellInst3_LFInst_3_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst3_LFInst_3_LFInst_2_U3  ( .A(SubCellInput2[12]), .B(
        SubCellInput2[13]), .ZN(SubCellInst3_LFInst_3_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst3_LFInst_3_LFInst_3_U9  ( .A1(
        SubCellInst3_LFInst_3_LFInst_3_n16 ), .A2(
        SubCellInst3_LFInst_3_LFInst_3_n15 ), .ZN(MCInst3_MC1_v3_2 [2]) );
  NAND2_X1 SubCellInst3_LFInst_3_LFInst_3_U8  ( .A1(SubCellInput2[13]), .A2(
        SubCellInst3_LFInst_3_LFInst_3_n14 ), .ZN(
        SubCellInst3_LFInst_3_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst3_LFInst_3_LFInst_3_U7  ( .A(SubCellInput2[15]), .B(
        SubCellInput2[14]), .Z(SubCellInst3_LFInst_3_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst3_LFInst_3_LFInst_3_U6  ( .A1(
        SubCellInst3_LFInst_3_LFInst_3_n13 ), .A2(
        SubCellInst3_LFInst_3_LFInst_3_n12 ), .ZN(
        SubCellInst3_LFInst_3_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst3_LFInst_3_LFInst_3_U5  ( .A1(SubCellInput2[12]), .A2(
        SubCellInput2[14]), .ZN(SubCellInst3_LFInst_3_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst3_LFInst_3_LFInst_3_U4  ( .A(SubCellInput2[12]), .B(
        SubCellInst3_LFInst_3_LFInst_3_n11 ), .ZN(
        SubCellInst3_LFInst_3_LFInst_3_n13 ) );
  OR2_X1 SubCellInst3_LFInst_3_LFInst_3_U3  ( .A1(SubCellInput2[15]), .A2(
        SubCellInput2[13]), .ZN(SubCellInst3_LFInst_3_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst3_LFInst_4_LFInst_0_U6  ( .A1(SubCellInput2[18]), .A2(
        SubCellInst3_LFInst_4_LFInst_0_n4 ), .ZN(
        SubCellInst3_LFInst_4_LFInst_0_n5 ) );
  INV_X1 SubCellInst3_LFInst_4_LFInst_0_U5  ( .A(SubCellInput2[17]), .ZN(
        SubCellInst3_LFInst_4_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst3_LFInst_4_LFInst_0_U4  ( .A(SubCellInput2[16]), .B(
        SubCellInput2[19]), .Z(SubCellInst3_LFInst_4_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst3_LFInst_4_LFInst_0_U3  ( .A(
        SubCellInst3_LFInst_4_LFInst_0_n6 ), .B(
        SubCellInst3_LFInst_4_LFInst_0_n5 ), .ZN(MCInst3_MC1_v2_3 [1]) );
  NAND2_X1 SubCellInst3_LFInst_4_LFInst_1_U12  ( .A1(
        SubCellInst3_LFInst_4_LFInst_1_n18 ), .A2(
        SubCellInst3_LFInst_4_LFInst_1_n17 ), .ZN(MCInst3_MC1_v2_0 [2]) );
  NAND2_X1 SubCellInst3_LFInst_4_LFInst_1_U11  ( .A1(SubCellInput2[17]), .A2(
        SubCellInst3_LFInst_4_LFInst_1_n16 ), .ZN(
        SubCellInst3_LFInst_4_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst3_LFInst_4_LFInst_1_U10  ( .A1(SubCellInput2[19]), .A2(
        SubCellInst3_LFInst_4_LFInst_1_n15 ), .ZN(
        SubCellInst3_LFInst_4_LFInst_1_n16 ) );
  AND2_X1 SubCellInst3_LFInst_4_LFInst_1_U9  ( .A1(SubCellInput2[16]), .A2(
        SubCellInput2[18]), .ZN(SubCellInst3_LFInst_4_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst3_LFInst_4_LFInst_1_U8  ( .A1(SubCellInput2[19]), .A2(
        SubCellInst3_LFInst_4_LFInst_1_n14 ), .ZN(
        SubCellInst3_LFInst_4_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst3_LFInst_4_LFInst_1_U7  ( .A1(
        SubCellInst3_LFInst_4_LFInst_1_n13 ), .A2(
        SubCellInst3_LFInst_4_LFInst_1_n12 ), .ZN(
        SubCellInst3_LFInst_4_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst3_LFInst_4_LFInst_1_U6  ( .A1(SubCellInput2[16]), .A2(
        SubCellInput2[18]), .ZN(SubCellInst3_LFInst_4_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst3_LFInst_4_LFInst_1_U5  ( .A1(
        SubCellInst3_LFInst_4_LFInst_1_n11 ), .A2(
        SubCellInst3_LFInst_4_LFInst_1_n10 ), .ZN(
        SubCellInst3_LFInst_4_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst3_LFInst_4_LFInst_1_U4  ( .A1(SubCellInput2[16]), .A2(
        SubCellInput2[17]), .ZN(SubCellInst3_LFInst_4_LFInst_1_n10 ) );
  INV_X1 SubCellInst3_LFInst_4_LFInst_1_U3  ( .A(SubCellInput2[18]), .ZN(
        SubCellInst3_LFInst_4_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst3_LFInst_4_LFInst_2_U11  ( .A1(
        SubCellInst3_LFInst_4_LFInst_2_n22 ), .A2(
        SubCellInst3_LFInst_4_LFInst_2_n21 ), .ZN(MCInst3_MC1_v2_0 [3]) );
  NAND2_X1 SubCellInst3_LFInst_4_LFInst_2_U10  ( .A1(SubCellInput2[18]), .A2(
        SubCellInst3_LFInst_4_LFInst_2_n20 ), .ZN(
        SubCellInst3_LFInst_4_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst3_LFInst_4_LFInst_2_U9  ( .A1(SubCellInput2[17]), .A2(
        SubCellInst3_LFInst_4_LFInst_2_n19 ), .ZN(
        SubCellInst3_LFInst_4_LFInst_2_n20 ) );
  INV_X1 SubCellInst3_LFInst_4_LFInst_2_U8  ( .A(SubCellInput2[19]), .ZN(
        SubCellInst3_LFInst_4_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst3_LFInst_4_LFInst_2_U7  ( .A1(
        SubCellInst3_LFInst_4_LFInst_2_n18 ), .A2(
        SubCellInst3_LFInst_4_LFInst_2_n17 ), .ZN(
        SubCellInst3_LFInst_4_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst3_LFInst_4_LFInst_2_U6  ( .A(
        SubCellInst3_LFInst_4_LFInst_2_n16 ), .B(SubCellInput2[18]), .Z(
        SubCellInst3_LFInst_4_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst3_LFInst_4_LFInst_2_U5  ( .A1(SubCellInput2[16]), .A2(
        SubCellInput2[17]), .ZN(SubCellInst3_LFInst_4_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst3_LFInst_4_LFInst_2_U4  ( .A1(
        SubCellInst3_LFInst_4_LFInst_2_n15 ), .A2(SubCellInput2[19]), .ZN(
        SubCellInst3_LFInst_4_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst3_LFInst_4_LFInst_2_U3  ( .A(SubCellInput2[16]), .B(
        SubCellInput2[17]), .ZN(SubCellInst3_LFInst_4_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst3_LFInst_4_LFInst_3_U9  ( .A1(
        SubCellInst3_LFInst_4_LFInst_3_n16 ), .A2(
        SubCellInst3_LFInst_4_LFInst_3_n15 ), .ZN(MCInst3_MC1_v2_0 [0]) );
  NAND2_X1 SubCellInst3_LFInst_4_LFInst_3_U8  ( .A1(SubCellInput2[17]), .A2(
        SubCellInst3_LFInst_4_LFInst_3_n14 ), .ZN(
        SubCellInst3_LFInst_4_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst3_LFInst_4_LFInst_3_U7  ( .A(SubCellInput2[19]), .B(
        SubCellInput2[18]), .Z(SubCellInst3_LFInst_4_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst3_LFInst_4_LFInst_3_U6  ( .A1(
        SubCellInst3_LFInst_4_LFInst_3_n13 ), .A2(
        SubCellInst3_LFInst_4_LFInst_3_n12 ), .ZN(
        SubCellInst3_LFInst_4_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst3_LFInst_4_LFInst_3_U5  ( .A1(SubCellInput2[16]), .A2(
        SubCellInput2[18]), .ZN(SubCellInst3_LFInst_4_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst3_LFInst_4_LFInst_3_U4  ( .A(SubCellInput2[16]), .B(
        SubCellInst3_LFInst_4_LFInst_3_n11 ), .ZN(
        SubCellInst3_LFInst_4_LFInst_3_n13 ) );
  OR2_X1 SubCellInst3_LFInst_4_LFInst_3_U3  ( .A1(SubCellInput2[19]), .A2(
        SubCellInput2[17]), .ZN(SubCellInst3_LFInst_4_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst3_LFInst_5_LFInst_0_U6  ( .A1(SubCellInput2[22]), .A2(
        SubCellInst3_LFInst_5_LFInst_0_n4 ), .ZN(
        SubCellInst3_LFInst_5_LFInst_0_n5 ) );
  INV_X1 SubCellInst3_LFInst_5_LFInst_0_U5  ( .A(SubCellInput2[21]), .ZN(
        SubCellInst3_LFInst_5_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst3_LFInst_5_LFInst_0_U4  ( .A(SubCellInput2[20]), .B(
        SubCellInput2[23]), .Z(SubCellInst3_LFInst_5_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst3_LFInst_5_LFInst_0_U3  ( .A(
        SubCellInst3_LFInst_5_LFInst_0_n6 ), .B(
        SubCellInst3_LFInst_5_LFInst_0_n5 ), .ZN(MCInst3_MC0_v2_3 [1]) );
  NAND2_X1 SubCellInst3_LFInst_5_LFInst_1_U12  ( .A1(
        SubCellInst3_LFInst_5_LFInst_1_n18 ), .A2(
        SubCellInst3_LFInst_5_LFInst_1_n17 ), .ZN(MCInst3_MC0_v2_0 [2]) );
  NAND2_X1 SubCellInst3_LFInst_5_LFInst_1_U11  ( .A1(SubCellInput2[21]), .A2(
        SubCellInst3_LFInst_5_LFInst_1_n16 ), .ZN(
        SubCellInst3_LFInst_5_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst3_LFInst_5_LFInst_1_U10  ( .A1(SubCellInput2[23]), .A2(
        SubCellInst3_LFInst_5_LFInst_1_n15 ), .ZN(
        SubCellInst3_LFInst_5_LFInst_1_n16 ) );
  AND2_X1 SubCellInst3_LFInst_5_LFInst_1_U9  ( .A1(SubCellInput2[20]), .A2(
        SubCellInput2[22]), .ZN(SubCellInst3_LFInst_5_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst3_LFInst_5_LFInst_1_U8  ( .A1(SubCellInput2[23]), .A2(
        SubCellInst3_LFInst_5_LFInst_1_n14 ), .ZN(
        SubCellInst3_LFInst_5_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst3_LFInst_5_LFInst_1_U7  ( .A1(
        SubCellInst3_LFInst_5_LFInst_1_n13 ), .A2(
        SubCellInst3_LFInst_5_LFInst_1_n12 ), .ZN(
        SubCellInst3_LFInst_5_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst3_LFInst_5_LFInst_1_U6  ( .A1(SubCellInput2[20]), .A2(
        SubCellInput2[22]), .ZN(SubCellInst3_LFInst_5_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst3_LFInst_5_LFInst_1_U5  ( .A1(
        SubCellInst3_LFInst_5_LFInst_1_n11 ), .A2(
        SubCellInst3_LFInst_5_LFInst_1_n10 ), .ZN(
        SubCellInst3_LFInst_5_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst3_LFInst_5_LFInst_1_U4  ( .A1(SubCellInput2[20]), .A2(
        SubCellInput2[21]), .ZN(SubCellInst3_LFInst_5_LFInst_1_n10 ) );
  INV_X1 SubCellInst3_LFInst_5_LFInst_1_U3  ( .A(SubCellInput2[22]), .ZN(
        SubCellInst3_LFInst_5_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst3_LFInst_5_LFInst_2_U11  ( .A1(
        SubCellInst3_LFInst_5_LFInst_2_n22 ), .A2(
        SubCellInst3_LFInst_5_LFInst_2_n21 ), .ZN(MCInst3_MC0_v2_0 [3]) );
  NAND2_X1 SubCellInst3_LFInst_5_LFInst_2_U10  ( .A1(SubCellInput2[22]), .A2(
        SubCellInst3_LFInst_5_LFInst_2_n20 ), .ZN(
        SubCellInst3_LFInst_5_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst3_LFInst_5_LFInst_2_U9  ( .A1(SubCellInput2[21]), .A2(
        SubCellInst3_LFInst_5_LFInst_2_n19 ), .ZN(
        SubCellInst3_LFInst_5_LFInst_2_n20 ) );
  INV_X1 SubCellInst3_LFInst_5_LFInst_2_U8  ( .A(SubCellInput2[23]), .ZN(
        SubCellInst3_LFInst_5_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst3_LFInst_5_LFInst_2_U7  ( .A1(
        SubCellInst3_LFInst_5_LFInst_2_n18 ), .A2(
        SubCellInst3_LFInst_5_LFInst_2_n17 ), .ZN(
        SubCellInst3_LFInst_5_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst3_LFInst_5_LFInst_2_U6  ( .A(
        SubCellInst3_LFInst_5_LFInst_2_n16 ), .B(SubCellInput2[22]), .Z(
        SubCellInst3_LFInst_5_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst3_LFInst_5_LFInst_2_U5  ( .A1(SubCellInput2[20]), .A2(
        SubCellInput2[21]), .ZN(SubCellInst3_LFInst_5_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst3_LFInst_5_LFInst_2_U4  ( .A1(
        SubCellInst3_LFInst_5_LFInst_2_n15 ), .A2(SubCellInput2[23]), .ZN(
        SubCellInst3_LFInst_5_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst3_LFInst_5_LFInst_2_U3  ( .A(SubCellInput2[20]), .B(
        SubCellInput2[21]), .ZN(SubCellInst3_LFInst_5_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst3_LFInst_5_LFInst_3_U9  ( .A1(
        SubCellInst3_LFInst_5_LFInst_3_n16 ), .A2(
        SubCellInst3_LFInst_5_LFInst_3_n15 ), .ZN(MCInst3_MC0_v2_0 [0]) );
  NAND2_X1 SubCellInst3_LFInst_5_LFInst_3_U8  ( .A1(SubCellInput2[21]), .A2(
        SubCellInst3_LFInst_5_LFInst_3_n14 ), .ZN(
        SubCellInst3_LFInst_5_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst3_LFInst_5_LFInst_3_U7  ( .A(SubCellInput2[23]), .B(
        SubCellInput2[22]), .Z(SubCellInst3_LFInst_5_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst3_LFInst_5_LFInst_3_U6  ( .A1(
        SubCellInst3_LFInst_5_LFInst_3_n13 ), .A2(
        SubCellInst3_LFInst_5_LFInst_3_n12 ), .ZN(
        SubCellInst3_LFInst_5_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst3_LFInst_5_LFInst_3_U5  ( .A1(SubCellInput2[20]), .A2(
        SubCellInput2[22]), .ZN(SubCellInst3_LFInst_5_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst3_LFInst_5_LFInst_3_U4  ( .A(SubCellInput2[20]), .B(
        SubCellInst3_LFInst_5_LFInst_3_n11 ), .ZN(
        SubCellInst3_LFInst_5_LFInst_3_n13 ) );
  OR2_X1 SubCellInst3_LFInst_5_LFInst_3_U3  ( .A1(SubCellInput2[23]), .A2(
        SubCellInput2[21]), .ZN(SubCellInst3_LFInst_5_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst3_LFInst_6_LFInst_0_U6  ( .A1(SubCellInput2[26]), .A2(
        SubCellInst3_LFInst_6_LFInst_0_n4 ), .ZN(
        SubCellInst3_LFInst_6_LFInst_0_n5 ) );
  INV_X1 SubCellInst3_LFInst_6_LFInst_0_U5  ( .A(SubCellInput2[25]), .ZN(
        SubCellInst3_LFInst_6_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst3_LFInst_6_LFInst_0_U4  ( .A(SubCellInput2[24]), .B(
        SubCellInput2[27]), .Z(SubCellInst3_LFInst_6_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst3_LFInst_6_LFInst_0_U3  ( .A(
        SubCellInst3_LFInst_6_LFInst_0_n6 ), .B(
        SubCellInst3_LFInst_6_LFInst_0_n5 ), .ZN(MCInst3_MC3_v2_3 [1]) );
  NAND2_X1 SubCellInst3_LFInst_6_LFInst_1_U12  ( .A1(
        SubCellInst3_LFInst_6_LFInst_1_n18 ), .A2(
        SubCellInst3_LFInst_6_LFInst_1_n17 ), .ZN(MCInst3_MC3_v2_0 [2]) );
  NAND2_X1 SubCellInst3_LFInst_6_LFInst_1_U11  ( .A1(SubCellInput2[25]), .A2(
        SubCellInst3_LFInst_6_LFInst_1_n16 ), .ZN(
        SubCellInst3_LFInst_6_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst3_LFInst_6_LFInst_1_U10  ( .A1(SubCellInput2[27]), .A2(
        SubCellInst3_LFInst_6_LFInst_1_n15 ), .ZN(
        SubCellInst3_LFInst_6_LFInst_1_n16 ) );
  AND2_X1 SubCellInst3_LFInst_6_LFInst_1_U9  ( .A1(SubCellInput2[24]), .A2(
        SubCellInput2[26]), .ZN(SubCellInst3_LFInst_6_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst3_LFInst_6_LFInst_1_U8  ( .A1(SubCellInput2[27]), .A2(
        SubCellInst3_LFInst_6_LFInst_1_n14 ), .ZN(
        SubCellInst3_LFInst_6_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst3_LFInst_6_LFInst_1_U7  ( .A1(
        SubCellInst3_LFInst_6_LFInst_1_n13 ), .A2(
        SubCellInst3_LFInst_6_LFInst_1_n12 ), .ZN(
        SubCellInst3_LFInst_6_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst3_LFInst_6_LFInst_1_U6  ( .A1(SubCellInput2[24]), .A2(
        SubCellInput2[26]), .ZN(SubCellInst3_LFInst_6_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst3_LFInst_6_LFInst_1_U5  ( .A1(
        SubCellInst3_LFInst_6_LFInst_1_n11 ), .A2(
        SubCellInst3_LFInst_6_LFInst_1_n10 ), .ZN(
        SubCellInst3_LFInst_6_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst3_LFInst_6_LFInst_1_U4  ( .A1(SubCellInput2[24]), .A2(
        SubCellInput2[25]), .ZN(SubCellInst3_LFInst_6_LFInst_1_n10 ) );
  INV_X1 SubCellInst3_LFInst_6_LFInst_1_U3  ( .A(SubCellInput2[26]), .ZN(
        SubCellInst3_LFInst_6_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst3_LFInst_6_LFInst_2_U11  ( .A1(
        SubCellInst3_LFInst_6_LFInst_2_n22 ), .A2(
        SubCellInst3_LFInst_6_LFInst_2_n21 ), .ZN(MCInst3_MC3_v2_0 [3]) );
  NAND2_X1 SubCellInst3_LFInst_6_LFInst_2_U10  ( .A1(SubCellInput2[26]), .A2(
        SubCellInst3_LFInst_6_LFInst_2_n20 ), .ZN(
        SubCellInst3_LFInst_6_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst3_LFInst_6_LFInst_2_U9  ( .A1(SubCellInput2[25]), .A2(
        SubCellInst3_LFInst_6_LFInst_2_n19 ), .ZN(
        SubCellInst3_LFInst_6_LFInst_2_n20 ) );
  INV_X1 SubCellInst3_LFInst_6_LFInst_2_U8  ( .A(SubCellInput2[27]), .ZN(
        SubCellInst3_LFInst_6_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst3_LFInst_6_LFInst_2_U7  ( .A1(
        SubCellInst3_LFInst_6_LFInst_2_n18 ), .A2(
        SubCellInst3_LFInst_6_LFInst_2_n17 ), .ZN(
        SubCellInst3_LFInst_6_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst3_LFInst_6_LFInst_2_U6  ( .A(
        SubCellInst3_LFInst_6_LFInst_2_n16 ), .B(SubCellInput2[26]), .Z(
        SubCellInst3_LFInst_6_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst3_LFInst_6_LFInst_2_U5  ( .A1(SubCellInput2[24]), .A2(
        SubCellInput2[25]), .ZN(SubCellInst3_LFInst_6_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst3_LFInst_6_LFInst_2_U4  ( .A1(
        SubCellInst3_LFInst_6_LFInst_2_n15 ), .A2(SubCellInput2[27]), .ZN(
        SubCellInst3_LFInst_6_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst3_LFInst_6_LFInst_2_U3  ( .A(SubCellInput2[24]), .B(
        SubCellInput2[25]), .ZN(SubCellInst3_LFInst_6_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst3_LFInst_6_LFInst_3_U9  ( .A1(
        SubCellInst3_LFInst_6_LFInst_3_n16 ), .A2(
        SubCellInst3_LFInst_6_LFInst_3_n15 ), .ZN(MCInst3_MC3_v2_0 [0]) );
  NAND2_X1 SubCellInst3_LFInst_6_LFInst_3_U8  ( .A1(SubCellInput2[25]), .A2(
        SubCellInst3_LFInst_6_LFInst_3_n14 ), .ZN(
        SubCellInst3_LFInst_6_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst3_LFInst_6_LFInst_3_U7  ( .A(SubCellInput2[27]), .B(
        SubCellInput2[26]), .Z(SubCellInst3_LFInst_6_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst3_LFInst_6_LFInst_3_U6  ( .A1(
        SubCellInst3_LFInst_6_LFInst_3_n13 ), .A2(
        SubCellInst3_LFInst_6_LFInst_3_n12 ), .ZN(
        SubCellInst3_LFInst_6_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst3_LFInst_6_LFInst_3_U5  ( .A1(SubCellInput2[24]), .A2(
        SubCellInput2[26]), .ZN(SubCellInst3_LFInst_6_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst3_LFInst_6_LFInst_3_U4  ( .A(SubCellInput2[24]), .B(
        SubCellInst3_LFInst_6_LFInst_3_n11 ), .ZN(
        SubCellInst3_LFInst_6_LFInst_3_n13 ) );
  OR2_X1 SubCellInst3_LFInst_6_LFInst_3_U3  ( .A1(SubCellInput2[27]), .A2(
        SubCellInput2[25]), .ZN(SubCellInst3_LFInst_6_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst3_LFInst_7_LFInst_0_U6  ( .A1(SubCellInput2[30]), .A2(
        SubCellInst3_LFInst_7_LFInst_0_n4 ), .ZN(
        SubCellInst3_LFInst_7_LFInst_0_n5 ) );
  INV_X1 SubCellInst3_LFInst_7_LFInst_0_U5  ( .A(SubCellInput2[29]), .ZN(
        SubCellInst3_LFInst_7_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst3_LFInst_7_LFInst_0_U4  ( .A(SubCellInput2[28]), .B(
        SubCellInput2[31]), .Z(SubCellInst3_LFInst_7_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst3_LFInst_7_LFInst_0_U3  ( .A(
        SubCellInst3_LFInst_7_LFInst_0_n6 ), .B(
        SubCellInst3_LFInst_7_LFInst_0_n5 ), .ZN(MCInst3_MC2_v2_3 [1]) );
  NAND2_X1 SubCellInst3_LFInst_7_LFInst_1_U12  ( .A1(
        SubCellInst3_LFInst_7_LFInst_1_n18 ), .A2(
        SubCellInst3_LFInst_7_LFInst_1_n17 ), .ZN(MCInst3_MC2_v2_0 [2]) );
  NAND2_X1 SubCellInst3_LFInst_7_LFInst_1_U11  ( .A1(SubCellInput2[29]), .A2(
        SubCellInst3_LFInst_7_LFInst_1_n16 ), .ZN(
        SubCellInst3_LFInst_7_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst3_LFInst_7_LFInst_1_U10  ( .A1(SubCellInput2[31]), .A2(
        SubCellInst3_LFInst_7_LFInst_1_n15 ), .ZN(
        SubCellInst3_LFInst_7_LFInst_1_n16 ) );
  AND2_X1 SubCellInst3_LFInst_7_LFInst_1_U9  ( .A1(SubCellInput2[28]), .A2(
        SubCellInput2[30]), .ZN(SubCellInst3_LFInst_7_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst3_LFInst_7_LFInst_1_U8  ( .A1(SubCellInput2[31]), .A2(
        SubCellInst3_LFInst_7_LFInst_1_n14 ), .ZN(
        SubCellInst3_LFInst_7_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst3_LFInst_7_LFInst_1_U7  ( .A1(
        SubCellInst3_LFInst_7_LFInst_1_n13 ), .A2(
        SubCellInst3_LFInst_7_LFInst_1_n12 ), .ZN(
        SubCellInst3_LFInst_7_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst3_LFInst_7_LFInst_1_U6  ( .A1(SubCellInput2[28]), .A2(
        SubCellInput2[30]), .ZN(SubCellInst3_LFInst_7_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst3_LFInst_7_LFInst_1_U5  ( .A1(
        SubCellInst3_LFInst_7_LFInst_1_n11 ), .A2(
        SubCellInst3_LFInst_7_LFInst_1_n10 ), .ZN(
        SubCellInst3_LFInst_7_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst3_LFInst_7_LFInst_1_U4  ( .A1(SubCellInput2[28]), .A2(
        SubCellInput2[29]), .ZN(SubCellInst3_LFInst_7_LFInst_1_n10 ) );
  INV_X1 SubCellInst3_LFInst_7_LFInst_1_U3  ( .A(SubCellInput2[30]), .ZN(
        SubCellInst3_LFInst_7_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst3_LFInst_7_LFInst_2_U11  ( .A1(
        SubCellInst3_LFInst_7_LFInst_2_n22 ), .A2(
        SubCellInst3_LFInst_7_LFInst_2_n21 ), .ZN(MCInst3_MC2_v2_0 [3]) );
  NAND2_X1 SubCellInst3_LFInst_7_LFInst_2_U10  ( .A1(SubCellInput2[30]), .A2(
        SubCellInst3_LFInst_7_LFInst_2_n20 ), .ZN(
        SubCellInst3_LFInst_7_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst3_LFInst_7_LFInst_2_U9  ( .A1(SubCellInput2[29]), .A2(
        SubCellInst3_LFInst_7_LFInst_2_n19 ), .ZN(
        SubCellInst3_LFInst_7_LFInst_2_n20 ) );
  INV_X1 SubCellInst3_LFInst_7_LFInst_2_U8  ( .A(SubCellInput2[31]), .ZN(
        SubCellInst3_LFInst_7_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst3_LFInst_7_LFInst_2_U7  ( .A1(
        SubCellInst3_LFInst_7_LFInst_2_n18 ), .A2(
        SubCellInst3_LFInst_7_LFInst_2_n17 ), .ZN(
        SubCellInst3_LFInst_7_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst3_LFInst_7_LFInst_2_U6  ( .A(
        SubCellInst3_LFInst_7_LFInst_2_n16 ), .B(SubCellInput2[30]), .Z(
        SubCellInst3_LFInst_7_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst3_LFInst_7_LFInst_2_U5  ( .A1(SubCellInput2[28]), .A2(
        SubCellInput2[29]), .ZN(SubCellInst3_LFInst_7_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst3_LFInst_7_LFInst_2_U4  ( .A1(
        SubCellInst3_LFInst_7_LFInst_2_n15 ), .A2(SubCellInput2[31]), .ZN(
        SubCellInst3_LFInst_7_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst3_LFInst_7_LFInst_2_U3  ( .A(SubCellInput2[28]), .B(
        SubCellInput2[29]), .ZN(SubCellInst3_LFInst_7_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst3_LFInst_7_LFInst_3_U9  ( .A1(
        SubCellInst3_LFInst_7_LFInst_3_n16 ), .A2(
        SubCellInst3_LFInst_7_LFInst_3_n15 ), .ZN(MCInst3_MC2_v2_0 [0]) );
  NAND2_X1 SubCellInst3_LFInst_7_LFInst_3_U8  ( .A1(SubCellInput2[29]), .A2(
        SubCellInst3_LFInst_7_LFInst_3_n14 ), .ZN(
        SubCellInst3_LFInst_7_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst3_LFInst_7_LFInst_3_U7  ( .A(SubCellInput2[31]), .B(
        SubCellInput2[30]), .Z(SubCellInst3_LFInst_7_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst3_LFInst_7_LFInst_3_U6  ( .A1(
        SubCellInst3_LFInst_7_LFInst_3_n13 ), .A2(
        SubCellInst3_LFInst_7_LFInst_3_n12 ), .ZN(
        SubCellInst3_LFInst_7_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst3_LFInst_7_LFInst_3_U5  ( .A1(SubCellInput2[28]), .A2(
        SubCellInput2[30]), .ZN(SubCellInst3_LFInst_7_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst3_LFInst_7_LFInst_3_U4  ( .A(SubCellInput2[28]), .B(
        SubCellInst3_LFInst_7_LFInst_3_n11 ), .ZN(
        SubCellInst3_LFInst_7_LFInst_3_n13 ) );
  OR2_X1 SubCellInst3_LFInst_7_LFInst_3_U3  ( .A1(SubCellInput2[31]), .A2(
        SubCellInput2[29]), .ZN(SubCellInst3_LFInst_7_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst3_LFInst_8_LFInst_0_U6  ( .A1(SubCellInput2[34]), .A2(
        SubCellInst3_LFInst_8_LFInst_0_n4 ), .ZN(
        SubCellInst3_LFInst_8_LFInst_0_n5 ) );
  INV_X1 SubCellInst3_LFInst_8_LFInst_0_U5  ( .A(SubCellInput2[33]), .ZN(
        SubCellInst3_LFInst_8_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst3_LFInst_8_LFInst_0_U4  ( .A(SubCellInput2[32]), .B(
        SubCellInput2[35]), .Z(SubCellInst3_LFInst_8_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst3_LFInst_8_LFInst_0_U3  ( .A(
        SubCellInst3_LFInst_8_LFInst_0_n6 ), .B(
        SubCellInst3_LFInst_8_LFInst_0_n5 ), .ZN(MCInst3_MC2_v1_0 [0]) );
  NAND2_X1 SubCellInst3_LFInst_8_LFInst_1_U12  ( .A1(
        SubCellInst3_LFInst_8_LFInst_1_n18 ), .A2(
        SubCellInst3_LFInst_8_LFInst_1_n17 ), .ZN(MCInst3_MC2_v1_3 [2]) );
  NAND2_X1 SubCellInst3_LFInst_8_LFInst_1_U11  ( .A1(SubCellInput2[33]), .A2(
        SubCellInst3_LFInst_8_LFInst_1_n16 ), .ZN(
        SubCellInst3_LFInst_8_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst3_LFInst_8_LFInst_1_U10  ( .A1(SubCellInput2[35]), .A2(
        SubCellInst3_LFInst_8_LFInst_1_n15 ), .ZN(
        SubCellInst3_LFInst_8_LFInst_1_n16 ) );
  AND2_X1 SubCellInst3_LFInst_8_LFInst_1_U9  ( .A1(SubCellInput2[32]), .A2(
        SubCellInput2[34]), .ZN(SubCellInst3_LFInst_8_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst3_LFInst_8_LFInst_1_U8  ( .A1(SubCellInput2[35]), .A2(
        SubCellInst3_LFInst_8_LFInst_1_n14 ), .ZN(
        SubCellInst3_LFInst_8_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst3_LFInst_8_LFInst_1_U7  ( .A1(
        SubCellInst3_LFInst_8_LFInst_1_n13 ), .A2(
        SubCellInst3_LFInst_8_LFInst_1_n12 ), .ZN(
        SubCellInst3_LFInst_8_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst3_LFInst_8_LFInst_1_U6  ( .A1(SubCellInput2[32]), .A2(
        SubCellInput2[34]), .ZN(SubCellInst3_LFInst_8_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst3_LFInst_8_LFInst_1_U5  ( .A1(
        SubCellInst3_LFInst_8_LFInst_1_n11 ), .A2(
        SubCellInst3_LFInst_8_LFInst_1_n10 ), .ZN(
        SubCellInst3_LFInst_8_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst3_LFInst_8_LFInst_1_U4  ( .A1(SubCellInput2[32]), .A2(
        SubCellInput2[33]), .ZN(SubCellInst3_LFInst_8_LFInst_1_n10 ) );
  INV_X1 SubCellInst3_LFInst_8_LFInst_1_U3  ( .A(SubCellInput2[34]), .ZN(
        SubCellInst3_LFInst_8_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst3_LFInst_8_LFInst_2_U11  ( .A1(
        SubCellInst3_LFInst_8_LFInst_2_n22 ), .A2(
        SubCellInst3_LFInst_8_LFInst_2_n21 ), .ZN(Red_MCInst3_MC2_v1_1[0] )
         );
  NAND2_X1 SubCellInst3_LFInst_8_LFInst_2_U10  ( .A1(SubCellInput2[34]), .A2(
        SubCellInst3_LFInst_8_LFInst_2_n20 ), .ZN(
        SubCellInst3_LFInst_8_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst3_LFInst_8_LFInst_2_U9  ( .A1(SubCellInput2[33]), .A2(
        SubCellInst3_LFInst_8_LFInst_2_n19 ), .ZN(
        SubCellInst3_LFInst_8_LFInst_2_n20 ) );
  INV_X1 SubCellInst3_LFInst_8_LFInst_2_U8  ( .A(SubCellInput2[35]), .ZN(
        SubCellInst3_LFInst_8_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst3_LFInst_8_LFInst_2_U7  ( .A1(
        SubCellInst3_LFInst_8_LFInst_2_n18 ), .A2(
        SubCellInst3_LFInst_8_LFInst_2_n17 ), .ZN(
        SubCellInst3_LFInst_8_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst3_LFInst_8_LFInst_2_U6  ( .A(
        SubCellInst3_LFInst_8_LFInst_2_n16 ), .B(SubCellInput2[34]), .Z(
        SubCellInst3_LFInst_8_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst3_LFInst_8_LFInst_2_U5  ( .A1(SubCellInput2[32]), .A2(
        SubCellInput2[33]), .ZN(SubCellInst3_LFInst_8_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst3_LFInst_8_LFInst_2_U4  ( .A1(
        SubCellInst3_LFInst_8_LFInst_2_n15 ), .A2(SubCellInput2[35]), .ZN(
        SubCellInst3_LFInst_8_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst3_LFInst_8_LFInst_2_U3  ( .A(SubCellInput2[32]), .B(
        SubCellInput2[33]), .ZN(SubCellInst3_LFInst_8_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst3_LFInst_8_LFInst_3_U9  ( .A1(
        SubCellInst3_LFInst_8_LFInst_3_n16 ), .A2(
        SubCellInst3_LFInst_8_LFInst_3_n15 ), .ZN(MCInst3_MC2_v1_0 [3]) );
  NAND2_X1 SubCellInst3_LFInst_8_LFInst_3_U8  ( .A1(SubCellInput2[33]), .A2(
        SubCellInst3_LFInst_8_LFInst_3_n14 ), .ZN(
        SubCellInst3_LFInst_8_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst3_LFInst_8_LFInst_3_U7  ( .A(SubCellInput2[35]), .B(
        SubCellInput2[34]), .Z(SubCellInst3_LFInst_8_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst3_LFInst_8_LFInst_3_U6  ( .A1(
        SubCellInst3_LFInst_8_LFInst_3_n13 ), .A2(
        SubCellInst3_LFInst_8_LFInst_3_n12 ), .ZN(
        SubCellInst3_LFInst_8_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst3_LFInst_8_LFInst_3_U5  ( .A1(SubCellInput2[32]), .A2(
        SubCellInput2[34]), .ZN(SubCellInst3_LFInst_8_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst3_LFInst_8_LFInst_3_U4  ( .A(SubCellInput2[32]), .B(
        SubCellInst3_LFInst_8_LFInst_3_n11 ), .ZN(
        SubCellInst3_LFInst_8_LFInst_3_n13 ) );
  OR2_X1 SubCellInst3_LFInst_8_LFInst_3_U3  ( .A1(SubCellInput2[35]), .A2(
        SubCellInput2[33]), .ZN(SubCellInst3_LFInst_8_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst3_LFInst_9_LFInst_0_U6  ( .A1(SubCellInput2[38]), .A2(
        SubCellInst3_LFInst_9_LFInst_0_n4 ), .ZN(
        SubCellInst3_LFInst_9_LFInst_0_n5 ) );
  INV_X1 SubCellInst3_LFInst_9_LFInst_0_U5  ( .A(SubCellInput2[37]), .ZN(
        SubCellInst3_LFInst_9_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst3_LFInst_9_LFInst_0_U4  ( .A(SubCellInput2[36]), .B(
        SubCellInput2[39]), .Z(SubCellInst3_LFInst_9_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst3_LFInst_9_LFInst_0_U3  ( .A(
        SubCellInst3_LFInst_9_LFInst_0_n6 ), .B(
        SubCellInst3_LFInst_9_LFInst_0_n5 ), .ZN(MCInst3_MC1_v1_0 [0]) );
  NAND2_X1 SubCellInst3_LFInst_9_LFInst_1_U12  ( .A1(
        SubCellInst3_LFInst_9_LFInst_1_n18 ), .A2(
        SubCellInst3_LFInst_9_LFInst_1_n17 ), .ZN(MCInst3_MC1_v1_3 [2]) );
  NAND2_X1 SubCellInst3_LFInst_9_LFInst_1_U11  ( .A1(SubCellInput2[37]), .A2(
        SubCellInst3_LFInst_9_LFInst_1_n16 ), .ZN(
        SubCellInst3_LFInst_9_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst3_LFInst_9_LFInst_1_U10  ( .A1(SubCellInput2[39]), .A2(
        SubCellInst3_LFInst_9_LFInst_1_n15 ), .ZN(
        SubCellInst3_LFInst_9_LFInst_1_n16 ) );
  AND2_X1 SubCellInst3_LFInst_9_LFInst_1_U9  ( .A1(SubCellInput2[36]), .A2(
        SubCellInput2[38]), .ZN(SubCellInst3_LFInst_9_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst3_LFInst_9_LFInst_1_U8  ( .A1(SubCellInput2[39]), .A2(
        SubCellInst3_LFInst_9_LFInst_1_n14 ), .ZN(
        SubCellInst3_LFInst_9_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst3_LFInst_9_LFInst_1_U7  ( .A1(
        SubCellInst3_LFInst_9_LFInst_1_n13 ), .A2(
        SubCellInst3_LFInst_9_LFInst_1_n12 ), .ZN(
        SubCellInst3_LFInst_9_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst3_LFInst_9_LFInst_1_U6  ( .A1(SubCellInput2[36]), .A2(
        SubCellInput2[38]), .ZN(SubCellInst3_LFInst_9_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst3_LFInst_9_LFInst_1_U5  ( .A1(
        SubCellInst3_LFInst_9_LFInst_1_n11 ), .A2(
        SubCellInst3_LFInst_9_LFInst_1_n10 ), .ZN(
        SubCellInst3_LFInst_9_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst3_LFInst_9_LFInst_1_U4  ( .A1(SubCellInput2[36]), .A2(
        SubCellInput2[37]), .ZN(SubCellInst3_LFInst_9_LFInst_1_n10 ) );
  INV_X1 SubCellInst3_LFInst_9_LFInst_1_U3  ( .A(SubCellInput2[38]), .ZN(
        SubCellInst3_LFInst_9_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst3_LFInst_9_LFInst_2_U11  ( .A1(
        SubCellInst3_LFInst_9_LFInst_2_n22 ), .A2(
        SubCellInst3_LFInst_9_LFInst_2_n21 ), .ZN(Red_MCInst3_MC1_v1_1[0] )
         );
  NAND2_X1 SubCellInst3_LFInst_9_LFInst_2_U10  ( .A1(SubCellInput2[38]), .A2(
        SubCellInst3_LFInst_9_LFInst_2_n20 ), .ZN(
        SubCellInst3_LFInst_9_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst3_LFInst_9_LFInst_2_U9  ( .A1(SubCellInput2[37]), .A2(
        SubCellInst3_LFInst_9_LFInst_2_n19 ), .ZN(
        SubCellInst3_LFInst_9_LFInst_2_n20 ) );
  INV_X1 SubCellInst3_LFInst_9_LFInst_2_U8  ( .A(SubCellInput2[39]), .ZN(
        SubCellInst3_LFInst_9_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst3_LFInst_9_LFInst_2_U7  ( .A1(
        SubCellInst3_LFInst_9_LFInst_2_n18 ), .A2(
        SubCellInst3_LFInst_9_LFInst_2_n17 ), .ZN(
        SubCellInst3_LFInst_9_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst3_LFInst_9_LFInst_2_U6  ( .A(
        SubCellInst3_LFInst_9_LFInst_2_n16 ), .B(SubCellInput2[38]), .Z(
        SubCellInst3_LFInst_9_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst3_LFInst_9_LFInst_2_U5  ( .A1(SubCellInput2[36]), .A2(
        SubCellInput2[37]), .ZN(SubCellInst3_LFInst_9_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst3_LFInst_9_LFInst_2_U4  ( .A1(
        SubCellInst3_LFInst_9_LFInst_2_n15 ), .A2(SubCellInput2[39]), .ZN(
        SubCellInst3_LFInst_9_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst3_LFInst_9_LFInst_2_U3  ( .A(SubCellInput2[36]), .B(
        SubCellInput2[37]), .ZN(SubCellInst3_LFInst_9_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst3_LFInst_9_LFInst_3_U9  ( .A1(
        SubCellInst3_LFInst_9_LFInst_3_n16 ), .A2(
        SubCellInst3_LFInst_9_LFInst_3_n15 ), .ZN(MCInst3_MC1_v1_0 [3]) );
  NAND2_X1 SubCellInst3_LFInst_9_LFInst_3_U8  ( .A1(SubCellInput2[37]), .A2(
        SubCellInst3_LFInst_9_LFInst_3_n14 ), .ZN(
        SubCellInst3_LFInst_9_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst3_LFInst_9_LFInst_3_U7  ( .A(SubCellInput2[39]), .B(
        SubCellInput2[38]), .Z(SubCellInst3_LFInst_9_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst3_LFInst_9_LFInst_3_U6  ( .A1(
        SubCellInst3_LFInst_9_LFInst_3_n13 ), .A2(
        SubCellInst3_LFInst_9_LFInst_3_n12 ), .ZN(
        SubCellInst3_LFInst_9_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst3_LFInst_9_LFInst_3_U5  ( .A1(SubCellInput2[36]), .A2(
        SubCellInput2[38]), .ZN(SubCellInst3_LFInst_9_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst3_LFInst_9_LFInst_3_U4  ( .A(SubCellInput2[36]), .B(
        SubCellInst3_LFInst_9_LFInst_3_n11 ), .ZN(
        SubCellInst3_LFInst_9_LFInst_3_n13 ) );
  OR2_X1 SubCellInst3_LFInst_9_LFInst_3_U3  ( .A1(SubCellInput2[39]), .A2(
        SubCellInput2[37]), .ZN(SubCellInst3_LFInst_9_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst3_LFInst_10_LFInst_0_U6  ( .A1(SubCellInput2[42]), .A2(
        SubCellInst3_LFInst_10_LFInst_0_n4 ), .ZN(
        SubCellInst3_LFInst_10_LFInst_0_n5 ) );
  INV_X1 SubCellInst3_LFInst_10_LFInst_0_U5  ( .A(SubCellInput2[41]), .ZN(
        SubCellInst3_LFInst_10_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst3_LFInst_10_LFInst_0_U4  ( .A(SubCellInput2[40]), .B(
        SubCellInput2[43]), .Z(SubCellInst3_LFInst_10_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst3_LFInst_10_LFInst_0_U3  ( .A(
        SubCellInst3_LFInst_10_LFInst_0_n6 ), .B(
        SubCellInst3_LFInst_10_LFInst_0_n5 ), .ZN(MCInst3_MC0_v1_0 [0]) );
  NAND2_X1 SubCellInst3_LFInst_10_LFInst_1_U12  ( .A1(
        SubCellInst3_LFInst_10_LFInst_1_n18 ), .A2(
        SubCellInst3_LFInst_10_LFInst_1_n17 ), .ZN(MCInst3_MC0_v1_3 [2]) );
  NAND2_X1 SubCellInst3_LFInst_10_LFInst_1_U11  ( .A1(SubCellInput2[41]), 
        .A2(SubCellInst3_LFInst_10_LFInst_1_n16 ), .ZN(
        SubCellInst3_LFInst_10_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst3_LFInst_10_LFInst_1_U10  ( .A1(SubCellInput2[43]), .A2(
        SubCellInst3_LFInst_10_LFInst_1_n15 ), .ZN(
        SubCellInst3_LFInst_10_LFInst_1_n16 ) );
  AND2_X1 SubCellInst3_LFInst_10_LFInst_1_U9  ( .A1(SubCellInput2[40]), .A2(
        SubCellInput2[42]), .ZN(SubCellInst3_LFInst_10_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst3_LFInst_10_LFInst_1_U8  ( .A1(SubCellInput2[43]), .A2(
        SubCellInst3_LFInst_10_LFInst_1_n14 ), .ZN(
        SubCellInst3_LFInst_10_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst3_LFInst_10_LFInst_1_U7  ( .A1(
        SubCellInst3_LFInst_10_LFInst_1_n13 ), .A2(
        SubCellInst3_LFInst_10_LFInst_1_n12 ), .ZN(
        SubCellInst3_LFInst_10_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst3_LFInst_10_LFInst_1_U6  ( .A1(SubCellInput2[40]), .A2(
        SubCellInput2[42]), .ZN(SubCellInst3_LFInst_10_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst3_LFInst_10_LFInst_1_U5  ( .A1(
        SubCellInst3_LFInst_10_LFInst_1_n11 ), .A2(
        SubCellInst3_LFInst_10_LFInst_1_n10 ), .ZN(
        SubCellInst3_LFInst_10_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst3_LFInst_10_LFInst_1_U4  ( .A1(SubCellInput2[40]), .A2(
        SubCellInput2[41]), .ZN(SubCellInst3_LFInst_10_LFInst_1_n10 ) );
  INV_X1 SubCellInst3_LFInst_10_LFInst_1_U3  ( .A(SubCellInput2[42]), .ZN(
        SubCellInst3_LFInst_10_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst3_LFInst_10_LFInst_2_U11  ( .A1(
        SubCellInst3_LFInst_10_LFInst_2_n22 ), .A2(
        SubCellInst3_LFInst_10_LFInst_2_n21 ), .ZN(Red_MCInst3_MC0_v1_1[0] )
         );
  NAND2_X1 SubCellInst3_LFInst_10_LFInst_2_U10  ( .A1(SubCellInput2[42]), 
        .A2(SubCellInst3_LFInst_10_LFInst_2_n20 ), .ZN(
        SubCellInst3_LFInst_10_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst3_LFInst_10_LFInst_2_U9  ( .A1(SubCellInput2[41]), .A2(
        SubCellInst3_LFInst_10_LFInst_2_n19 ), .ZN(
        SubCellInst3_LFInst_10_LFInst_2_n20 ) );
  INV_X1 SubCellInst3_LFInst_10_LFInst_2_U8  ( .A(SubCellInput2[43]), .ZN(
        SubCellInst3_LFInst_10_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst3_LFInst_10_LFInst_2_U7  ( .A1(
        SubCellInst3_LFInst_10_LFInst_2_n18 ), .A2(
        SubCellInst3_LFInst_10_LFInst_2_n17 ), .ZN(
        SubCellInst3_LFInst_10_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst3_LFInst_10_LFInst_2_U6  ( .A(
        SubCellInst3_LFInst_10_LFInst_2_n16 ), .B(SubCellInput2[42]), .Z(
        SubCellInst3_LFInst_10_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst3_LFInst_10_LFInst_2_U5  ( .A1(SubCellInput2[40]), .A2(
        SubCellInput2[41]), .ZN(SubCellInst3_LFInst_10_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst3_LFInst_10_LFInst_2_U4  ( .A1(
        SubCellInst3_LFInst_10_LFInst_2_n15 ), .A2(SubCellInput2[43]), .ZN(
        SubCellInst3_LFInst_10_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst3_LFInst_10_LFInst_2_U3  ( .A(SubCellInput2[40]), .B(
        SubCellInput2[41]), .ZN(SubCellInst3_LFInst_10_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst3_LFInst_10_LFInst_3_U9  ( .A1(
        SubCellInst3_LFInst_10_LFInst_3_n16 ), .A2(
        SubCellInst3_LFInst_10_LFInst_3_n15 ), .ZN(MCInst3_MC0_v1_0 [3]) );
  NAND2_X1 SubCellInst3_LFInst_10_LFInst_3_U8  ( .A1(SubCellInput2[41]), .A2(
        SubCellInst3_LFInst_10_LFInst_3_n14 ), .ZN(
        SubCellInst3_LFInst_10_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst3_LFInst_10_LFInst_3_U7  ( .A(SubCellInput2[43]), .B(
        SubCellInput2[42]), .Z(SubCellInst3_LFInst_10_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst3_LFInst_10_LFInst_3_U6  ( .A1(
        SubCellInst3_LFInst_10_LFInst_3_n13 ), .A2(
        SubCellInst3_LFInst_10_LFInst_3_n12 ), .ZN(
        SubCellInst3_LFInst_10_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst3_LFInst_10_LFInst_3_U5  ( .A1(SubCellInput2[40]), .A2(
        SubCellInput2[42]), .ZN(SubCellInst3_LFInst_10_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst3_LFInst_10_LFInst_3_U4  ( .A(SubCellInput2[40]), .B(
        SubCellInst3_LFInst_10_LFInst_3_n11 ), .ZN(
        SubCellInst3_LFInst_10_LFInst_3_n13 ) );
  OR2_X1 SubCellInst3_LFInst_10_LFInst_3_U3  ( .A1(SubCellInput2[43]), .A2(
        SubCellInput2[41]), .ZN(SubCellInst3_LFInst_10_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst3_LFInst_11_LFInst_0_U6  ( .A1(SubCellInput2[46]), .A2(
        SubCellInst3_LFInst_11_LFInst_0_n4 ), .ZN(
        SubCellInst3_LFInst_11_LFInst_0_n5 ) );
  INV_X1 SubCellInst3_LFInst_11_LFInst_0_U5  ( .A(SubCellInput2[45]), .ZN(
        SubCellInst3_LFInst_11_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst3_LFInst_11_LFInst_0_U4  ( .A(SubCellInput2[44]), .B(
        SubCellInput2[47]), .Z(SubCellInst3_LFInst_11_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst3_LFInst_11_LFInst_0_U3  ( .A(
        SubCellInst3_LFInst_11_LFInst_0_n6 ), .B(
        SubCellInst3_LFInst_11_LFInst_0_n5 ), .ZN(MCInst3_MC3_v1_0 [0]) );
  NAND2_X1 SubCellInst3_LFInst_11_LFInst_1_U12  ( .A1(
        SubCellInst3_LFInst_11_LFInst_1_n18 ), .A2(
        SubCellInst3_LFInst_11_LFInst_1_n17 ), .ZN(MCInst3_MC3_v1_3 [2]) );
  NAND2_X1 SubCellInst3_LFInst_11_LFInst_1_U11  ( .A1(SubCellInput2[45]), 
        .A2(SubCellInst3_LFInst_11_LFInst_1_n16 ), .ZN(
        SubCellInst3_LFInst_11_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst3_LFInst_11_LFInst_1_U10  ( .A1(SubCellInput2[47]), .A2(
        SubCellInst3_LFInst_11_LFInst_1_n15 ), .ZN(
        SubCellInst3_LFInst_11_LFInst_1_n16 ) );
  AND2_X1 SubCellInst3_LFInst_11_LFInst_1_U9  ( .A1(SubCellInput2[44]), .A2(
        SubCellInput2[46]), .ZN(SubCellInst3_LFInst_11_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst3_LFInst_11_LFInst_1_U8  ( .A1(SubCellInput2[47]), .A2(
        SubCellInst3_LFInst_11_LFInst_1_n14 ), .ZN(
        SubCellInst3_LFInst_11_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst3_LFInst_11_LFInst_1_U7  ( .A1(
        SubCellInst3_LFInst_11_LFInst_1_n13 ), .A2(
        SubCellInst3_LFInst_11_LFInst_1_n12 ), .ZN(
        SubCellInst3_LFInst_11_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst3_LFInst_11_LFInst_1_U6  ( .A1(SubCellInput2[44]), .A2(
        SubCellInput2[46]), .ZN(SubCellInst3_LFInst_11_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst3_LFInst_11_LFInst_1_U5  ( .A1(
        SubCellInst3_LFInst_11_LFInst_1_n11 ), .A2(
        SubCellInst3_LFInst_11_LFInst_1_n10 ), .ZN(
        SubCellInst3_LFInst_11_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst3_LFInst_11_LFInst_1_U4  ( .A1(SubCellInput2[44]), .A2(
        SubCellInput2[45]), .ZN(SubCellInst3_LFInst_11_LFInst_1_n10 ) );
  INV_X1 SubCellInst3_LFInst_11_LFInst_1_U3  ( .A(SubCellInput2[46]), .ZN(
        SubCellInst3_LFInst_11_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst3_LFInst_11_LFInst_2_U11  ( .A1(
        SubCellInst3_LFInst_11_LFInst_2_n22 ), .A2(
        SubCellInst3_LFInst_11_LFInst_2_n21 ), .ZN(Red_MCInst3_MC3_v1_1[0] )
         );
  NAND2_X1 SubCellInst3_LFInst_11_LFInst_2_U10  ( .A1(SubCellInput2[46]), 
        .A2(SubCellInst3_LFInst_11_LFInst_2_n20 ), .ZN(
        SubCellInst3_LFInst_11_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst3_LFInst_11_LFInst_2_U9  ( .A1(SubCellInput2[45]), .A2(
        SubCellInst3_LFInst_11_LFInst_2_n19 ), .ZN(
        SubCellInst3_LFInst_11_LFInst_2_n20 ) );
  INV_X1 SubCellInst3_LFInst_11_LFInst_2_U8  ( .A(SubCellInput2[47]), .ZN(
        SubCellInst3_LFInst_11_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst3_LFInst_11_LFInst_2_U7  ( .A1(
        SubCellInst3_LFInst_11_LFInst_2_n18 ), .A2(
        SubCellInst3_LFInst_11_LFInst_2_n17 ), .ZN(
        SubCellInst3_LFInst_11_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst3_LFInst_11_LFInst_2_U6  ( .A(
        SubCellInst3_LFInst_11_LFInst_2_n16 ), .B(SubCellInput2[46]), .Z(
        SubCellInst3_LFInst_11_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst3_LFInst_11_LFInst_2_U5  ( .A1(SubCellInput2[44]), .A2(
        SubCellInput2[45]), .ZN(SubCellInst3_LFInst_11_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst3_LFInst_11_LFInst_2_U4  ( .A1(
        SubCellInst3_LFInst_11_LFInst_2_n15 ), .A2(SubCellInput2[47]), .ZN(
        SubCellInst3_LFInst_11_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst3_LFInst_11_LFInst_2_U3  ( .A(SubCellInput2[44]), .B(
        SubCellInput2[45]), .ZN(SubCellInst3_LFInst_11_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst3_LFInst_11_LFInst_3_U9  ( .A1(
        SubCellInst3_LFInst_11_LFInst_3_n16 ), .A2(
        SubCellInst3_LFInst_11_LFInst_3_n15 ), .ZN(MCInst3_MC3_v1_0 [3]) );
  NAND2_X1 SubCellInst3_LFInst_11_LFInst_3_U8  ( .A1(SubCellInput2[45]), .A2(
        SubCellInst3_LFInst_11_LFInst_3_n14 ), .ZN(
        SubCellInst3_LFInst_11_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst3_LFInst_11_LFInst_3_U7  ( .A(SubCellInput2[47]), .B(
        SubCellInput2[46]), .Z(SubCellInst3_LFInst_11_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst3_LFInst_11_LFInst_3_U6  ( .A1(
        SubCellInst3_LFInst_11_LFInst_3_n13 ), .A2(
        SubCellInst3_LFInst_11_LFInst_3_n12 ), .ZN(
        SubCellInst3_LFInst_11_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst3_LFInst_11_LFInst_3_U5  ( .A1(SubCellInput2[44]), .A2(
        SubCellInput2[46]), .ZN(SubCellInst3_LFInst_11_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst3_LFInst_11_LFInst_3_U4  ( .A(SubCellInput2[44]), .B(
        SubCellInst3_LFInst_11_LFInst_3_n11 ), .ZN(
        SubCellInst3_LFInst_11_LFInst_3_n13 ) );
  OR2_X1 SubCellInst3_LFInst_11_LFInst_3_U3  ( .A1(SubCellInput2[47]), .A2(
        SubCellInput2[45]), .ZN(SubCellInst3_LFInst_11_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst3_LFInst_12_LFInst_0_U6  ( .A1(SubCellInput2[50]), .A2(
        SubCellInst3_LFInst_12_LFInst_0_n4 ), .ZN(
        SubCellInst3_LFInst_12_LFInst_0_n5 ) );
  INV_X1 SubCellInst3_LFInst_12_LFInst_0_U5  ( .A(SubCellInput2[49]), .ZN(
        SubCellInst3_LFInst_12_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst3_LFInst_12_LFInst_0_U4  ( .A(SubCellInput2[48]), .B(
        SubCellInput2[51]), .Z(SubCellInst3_LFInst_12_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst3_LFInst_12_LFInst_0_U3  ( .A(
        SubCellInst3_LFInst_12_LFInst_0_n6 ), .B(
        SubCellInst3_LFInst_12_LFInst_0_n5 ), .ZN(Red_MCInst3_MC3_v0_1[0] )
         );
  NAND2_X1 SubCellInst3_LFInst_12_LFInst_1_U12  ( .A1(
        SubCellInst3_LFInst_12_LFInst_1_n18 ), .A2(
        SubCellInst3_LFInst_12_LFInst_1_n17 ), .ZN(MCInst3_MC3_v0_0 [3]) );
  NAND2_X1 SubCellInst3_LFInst_12_LFInst_1_U11  ( .A1(SubCellInput2[49]), 
        .A2(SubCellInst3_LFInst_12_LFInst_1_n16 ), .ZN(
        SubCellInst3_LFInst_12_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst3_LFInst_12_LFInst_1_U10  ( .A1(SubCellInput2[51]), .A2(
        SubCellInst3_LFInst_12_LFInst_1_n15 ), .ZN(
        SubCellInst3_LFInst_12_LFInst_1_n16 ) );
  AND2_X1 SubCellInst3_LFInst_12_LFInst_1_U9  ( .A1(SubCellInput2[48]), .A2(
        SubCellInput2[50]), .ZN(SubCellInst3_LFInst_12_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst3_LFInst_12_LFInst_1_U8  ( .A1(SubCellInput2[51]), .A2(
        SubCellInst3_LFInst_12_LFInst_1_n14 ), .ZN(
        SubCellInst3_LFInst_12_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst3_LFInst_12_LFInst_1_U7  ( .A1(
        SubCellInst3_LFInst_12_LFInst_1_n13 ), .A2(
        SubCellInst3_LFInst_12_LFInst_1_n12 ), .ZN(
        SubCellInst3_LFInst_12_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst3_LFInst_12_LFInst_1_U6  ( .A1(SubCellInput2[48]), .A2(
        SubCellInput2[50]), .ZN(SubCellInst3_LFInst_12_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst3_LFInst_12_LFInst_1_U5  ( .A1(
        SubCellInst3_LFInst_12_LFInst_1_n11 ), .A2(
        SubCellInst3_LFInst_12_LFInst_1_n10 ), .ZN(
        SubCellInst3_LFInst_12_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst3_LFInst_12_LFInst_1_U4  ( .A1(SubCellInput2[48]), .A2(
        SubCellInput2[49]), .ZN(SubCellInst3_LFInst_12_LFInst_1_n10 ) );
  INV_X1 SubCellInst3_LFInst_12_LFInst_1_U3  ( .A(SubCellInput2[50]), .ZN(
        SubCellInst3_LFInst_12_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst3_LFInst_12_LFInst_2_U11  ( .A1(
        SubCellInst3_LFInst_12_LFInst_2_n22 ), .A2(
        SubCellInst3_LFInst_12_LFInst_2_n21 ), .ZN(MCInst3_MC3_v0_3 [3]) );
  NAND2_X1 SubCellInst3_LFInst_12_LFInst_2_U10  ( .A1(SubCellInput2[50]), 
        .A2(SubCellInst3_LFInst_12_LFInst_2_n20 ), .ZN(
        SubCellInst3_LFInst_12_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst3_LFInst_12_LFInst_2_U9  ( .A1(SubCellInput2[49]), .A2(
        SubCellInst3_LFInst_12_LFInst_2_n19 ), .ZN(
        SubCellInst3_LFInst_12_LFInst_2_n20 ) );
  INV_X1 SubCellInst3_LFInst_12_LFInst_2_U8  ( .A(SubCellInput2[51]), .ZN(
        SubCellInst3_LFInst_12_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst3_LFInst_12_LFInst_2_U7  ( .A1(
        SubCellInst3_LFInst_12_LFInst_2_n18 ), .A2(
        SubCellInst3_LFInst_12_LFInst_2_n17 ), .ZN(
        SubCellInst3_LFInst_12_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst3_LFInst_12_LFInst_2_U6  ( .A(
        SubCellInst3_LFInst_12_LFInst_2_n16 ), .B(SubCellInput2[50]), .Z(
        SubCellInst3_LFInst_12_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst3_LFInst_12_LFInst_2_U5  ( .A1(SubCellInput2[48]), .A2(
        SubCellInput2[49]), .ZN(SubCellInst3_LFInst_12_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst3_LFInst_12_LFInst_2_U4  ( .A1(
        SubCellInst3_LFInst_12_LFInst_2_n15 ), .A2(SubCellInput2[51]), .ZN(
        SubCellInst3_LFInst_12_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst3_LFInst_12_LFInst_2_U3  ( .A(SubCellInput2[48]), .B(
        SubCellInput2[49]), .ZN(SubCellInst3_LFInst_12_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst3_LFInst_12_LFInst_3_U9  ( .A1(
        SubCellInst3_LFInst_12_LFInst_3_n16 ), .A2(
        SubCellInst3_LFInst_12_LFInst_3_n15 ), .ZN(MCInst3_MC3_v0_3 [0]) );
  NAND2_X1 SubCellInst3_LFInst_12_LFInst_3_U8  ( .A1(SubCellInput2[49]), .A2(
        SubCellInst3_LFInst_12_LFInst_3_n14 ), .ZN(
        SubCellInst3_LFInst_12_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst3_LFInst_12_LFInst_3_U7  ( .A(SubCellInput2[51]), .B(
        SubCellInput2[50]), .Z(SubCellInst3_LFInst_12_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst3_LFInst_12_LFInst_3_U6  ( .A1(
        SubCellInst3_LFInst_12_LFInst_3_n13 ), .A2(
        SubCellInst3_LFInst_12_LFInst_3_n12 ), .ZN(
        SubCellInst3_LFInst_12_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst3_LFInst_12_LFInst_3_U5  ( .A1(SubCellInput2[48]), .A2(
        SubCellInput2[50]), .ZN(SubCellInst3_LFInst_12_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst3_LFInst_12_LFInst_3_U4  ( .A(SubCellInput2[48]), .B(
        SubCellInst3_LFInst_12_LFInst_3_n11 ), .ZN(
        SubCellInst3_LFInst_12_LFInst_3_n13 ) );
  OR2_X1 SubCellInst3_LFInst_12_LFInst_3_U3  ( .A1(SubCellInput2[51]), .A2(
        SubCellInput2[49]), .ZN(SubCellInst3_LFInst_12_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst3_LFInst_13_LFInst_0_U6  ( .A1(SubCellInput2[54]), .A2(
        SubCellInst3_LFInst_13_LFInst_0_n4 ), .ZN(
        SubCellInst3_LFInst_13_LFInst_0_n5 ) );
  INV_X1 SubCellInst3_LFInst_13_LFInst_0_U5  ( .A(SubCellInput2[53]), .ZN(
        SubCellInst3_LFInst_13_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst3_LFInst_13_LFInst_0_U4  ( .A(SubCellInput2[52]), .B(
        SubCellInput2[55]), .Z(SubCellInst3_LFInst_13_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst3_LFInst_13_LFInst_0_U3  ( .A(
        SubCellInst3_LFInst_13_LFInst_0_n6 ), .B(
        SubCellInst3_LFInst_13_LFInst_0_n5 ), .ZN(Red_MCInst3_MC2_v0_1[0] )
         );
  NAND2_X1 SubCellInst3_LFInst_13_LFInst_1_U12  ( .A1(
        SubCellInst3_LFInst_13_LFInst_1_n18 ), .A2(
        SubCellInst3_LFInst_13_LFInst_1_n17 ), .ZN(MCInst3_MC2_v0_0 [3]) );
  NAND2_X1 SubCellInst3_LFInst_13_LFInst_1_U11  ( .A1(SubCellInput2[53]), 
        .A2(SubCellInst3_LFInst_13_LFInst_1_n16 ), .ZN(
        SubCellInst3_LFInst_13_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst3_LFInst_13_LFInst_1_U10  ( .A1(SubCellInput2[55]), .A2(
        SubCellInst3_LFInst_13_LFInst_1_n15 ), .ZN(
        SubCellInst3_LFInst_13_LFInst_1_n16 ) );
  AND2_X1 SubCellInst3_LFInst_13_LFInst_1_U9  ( .A1(SubCellInput2[52]), .A2(
        SubCellInput2[54]), .ZN(SubCellInst3_LFInst_13_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst3_LFInst_13_LFInst_1_U8  ( .A1(SubCellInput2[55]), .A2(
        SubCellInst3_LFInst_13_LFInst_1_n14 ), .ZN(
        SubCellInst3_LFInst_13_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst3_LFInst_13_LFInst_1_U7  ( .A1(
        SubCellInst3_LFInst_13_LFInst_1_n13 ), .A2(
        SubCellInst3_LFInst_13_LFInst_1_n12 ), .ZN(
        SubCellInst3_LFInst_13_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst3_LFInst_13_LFInst_1_U6  ( .A1(SubCellInput2[52]), .A2(
        SubCellInput2[54]), .ZN(SubCellInst3_LFInst_13_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst3_LFInst_13_LFInst_1_U5  ( .A1(
        SubCellInst3_LFInst_13_LFInst_1_n11 ), .A2(
        SubCellInst3_LFInst_13_LFInst_1_n10 ), .ZN(
        SubCellInst3_LFInst_13_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst3_LFInst_13_LFInst_1_U4  ( .A1(SubCellInput2[52]), .A2(
        SubCellInput2[53]), .ZN(SubCellInst3_LFInst_13_LFInst_1_n10 ) );
  INV_X1 SubCellInst3_LFInst_13_LFInst_1_U3  ( .A(SubCellInput2[54]), .ZN(
        SubCellInst3_LFInst_13_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst3_LFInst_13_LFInst_2_U11  ( .A1(
        SubCellInst3_LFInst_13_LFInst_2_n22 ), .A2(
        SubCellInst3_LFInst_13_LFInst_2_n21 ), .ZN(MCInst3_MC2_v0_3 [3]) );
  NAND2_X1 SubCellInst3_LFInst_13_LFInst_2_U10  ( .A1(SubCellInput2[54]), 
        .A2(SubCellInst3_LFInst_13_LFInst_2_n20 ), .ZN(
        SubCellInst3_LFInst_13_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst3_LFInst_13_LFInst_2_U9  ( .A1(SubCellInput2[53]), .A2(
        SubCellInst3_LFInst_13_LFInst_2_n19 ), .ZN(
        SubCellInst3_LFInst_13_LFInst_2_n20 ) );
  INV_X1 SubCellInst3_LFInst_13_LFInst_2_U8  ( .A(SubCellInput2[55]), .ZN(
        SubCellInst3_LFInst_13_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst3_LFInst_13_LFInst_2_U7  ( .A1(
        SubCellInst3_LFInst_13_LFInst_2_n18 ), .A2(
        SubCellInst3_LFInst_13_LFInst_2_n17 ), .ZN(
        SubCellInst3_LFInst_13_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst3_LFInst_13_LFInst_2_U6  ( .A(
        SubCellInst3_LFInst_13_LFInst_2_n16 ), .B(SubCellInput2[54]), .Z(
        SubCellInst3_LFInst_13_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst3_LFInst_13_LFInst_2_U5  ( .A1(SubCellInput2[52]), .A2(
        SubCellInput2[53]), .ZN(SubCellInst3_LFInst_13_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst3_LFInst_13_LFInst_2_U4  ( .A1(
        SubCellInst3_LFInst_13_LFInst_2_n15 ), .A2(SubCellInput2[55]), .ZN(
        SubCellInst3_LFInst_13_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst3_LFInst_13_LFInst_2_U3  ( .A(SubCellInput2[52]), .B(
        SubCellInput2[53]), .ZN(SubCellInst3_LFInst_13_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst3_LFInst_13_LFInst_3_U9  ( .A1(
        SubCellInst3_LFInst_13_LFInst_3_n16 ), .A2(
        SubCellInst3_LFInst_13_LFInst_3_n15 ), .ZN(MCInst3_MC2_v0_3 [0]) );
  NAND2_X1 SubCellInst3_LFInst_13_LFInst_3_U8  ( .A1(SubCellInput2[53]), .A2(
        SubCellInst3_LFInst_13_LFInst_3_n14 ), .ZN(
        SubCellInst3_LFInst_13_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst3_LFInst_13_LFInst_3_U7  ( .A(SubCellInput2[55]), .B(
        SubCellInput2[54]), .Z(SubCellInst3_LFInst_13_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst3_LFInst_13_LFInst_3_U6  ( .A1(
        SubCellInst3_LFInst_13_LFInst_3_n13 ), .A2(
        SubCellInst3_LFInst_13_LFInst_3_n12 ), .ZN(
        SubCellInst3_LFInst_13_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst3_LFInst_13_LFInst_3_U5  ( .A1(SubCellInput2[52]), .A2(
        SubCellInput2[54]), .ZN(SubCellInst3_LFInst_13_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst3_LFInst_13_LFInst_3_U4  ( .A(SubCellInput2[52]), .B(
        SubCellInst3_LFInst_13_LFInst_3_n11 ), .ZN(
        SubCellInst3_LFInst_13_LFInst_3_n13 ) );
  OR2_X1 SubCellInst3_LFInst_13_LFInst_3_U3  ( .A1(SubCellInput2[55]), .A2(
        SubCellInput2[53]), .ZN(SubCellInst3_LFInst_13_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst3_LFInst_14_LFInst_0_U6  ( .A1(SubCellInput2[58]), .A2(
        SubCellInst3_LFInst_14_LFInst_0_n4 ), .ZN(
        SubCellInst3_LFInst_14_LFInst_0_n5 ) );
  INV_X1 SubCellInst3_LFInst_14_LFInst_0_U5  ( .A(SubCellInput2[57]), .ZN(
        SubCellInst3_LFInst_14_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst3_LFInst_14_LFInst_0_U4  ( .A(SubCellInput2[56]), .B(
        SubCellInput2[59]), .Z(SubCellInst3_LFInst_14_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst3_LFInst_14_LFInst_0_U3  ( .A(
        SubCellInst3_LFInst_14_LFInst_0_n6 ), .B(
        SubCellInst3_LFInst_14_LFInst_0_n5 ), .ZN(Red_MCInst3_MC1_v0_1[0] )
         );
  NAND2_X1 SubCellInst3_LFInst_14_LFInst_1_U12  ( .A1(
        SubCellInst3_LFInst_14_LFInst_1_n18 ), .A2(
        SubCellInst3_LFInst_14_LFInst_1_n17 ), .ZN(MCInst3_MC1_v0_0 [3]) );
  NAND2_X1 SubCellInst3_LFInst_14_LFInst_1_U11  ( .A1(SubCellInput2[57]), 
        .A2(SubCellInst3_LFInst_14_LFInst_1_n16 ), .ZN(
        SubCellInst3_LFInst_14_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst3_LFInst_14_LFInst_1_U10  ( .A1(SubCellInput2[59]), .A2(
        SubCellInst3_LFInst_14_LFInst_1_n15 ), .ZN(
        SubCellInst3_LFInst_14_LFInst_1_n16 ) );
  AND2_X1 SubCellInst3_LFInst_14_LFInst_1_U9  ( .A1(SubCellInput2[56]), .A2(
        SubCellInput2[58]), .ZN(SubCellInst3_LFInst_14_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst3_LFInst_14_LFInst_1_U8  ( .A1(SubCellInput2[59]), .A2(
        SubCellInst3_LFInst_14_LFInst_1_n14 ), .ZN(
        SubCellInst3_LFInst_14_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst3_LFInst_14_LFInst_1_U7  ( .A1(
        SubCellInst3_LFInst_14_LFInst_1_n13 ), .A2(
        SubCellInst3_LFInst_14_LFInst_1_n12 ), .ZN(
        SubCellInst3_LFInst_14_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst3_LFInst_14_LFInst_1_U6  ( .A1(SubCellInput2[56]), .A2(
        SubCellInput2[58]), .ZN(SubCellInst3_LFInst_14_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst3_LFInst_14_LFInst_1_U5  ( .A1(
        SubCellInst3_LFInst_14_LFInst_1_n11 ), .A2(
        SubCellInst3_LFInst_14_LFInst_1_n10 ), .ZN(
        SubCellInst3_LFInst_14_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst3_LFInst_14_LFInst_1_U4  ( .A1(SubCellInput2[56]), .A2(
        SubCellInput2[57]), .ZN(SubCellInst3_LFInst_14_LFInst_1_n10 ) );
  INV_X1 SubCellInst3_LFInst_14_LFInst_1_U3  ( .A(SubCellInput2[58]), .ZN(
        SubCellInst3_LFInst_14_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst3_LFInst_14_LFInst_2_U11  ( .A1(
        SubCellInst3_LFInst_14_LFInst_2_n22 ), .A2(
        SubCellInst3_LFInst_14_LFInst_2_n21 ), .ZN(MCInst3_MC1_v0_3 [3]) );
  NAND2_X1 SubCellInst3_LFInst_14_LFInst_2_U10  ( .A1(SubCellInput2[58]), 
        .A2(SubCellInst3_LFInst_14_LFInst_2_n20 ), .ZN(
        SubCellInst3_LFInst_14_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst3_LFInst_14_LFInst_2_U9  ( .A1(SubCellInput2[57]), .A2(
        SubCellInst3_LFInst_14_LFInst_2_n19 ), .ZN(
        SubCellInst3_LFInst_14_LFInst_2_n20 ) );
  INV_X1 SubCellInst3_LFInst_14_LFInst_2_U8  ( .A(SubCellInput2[59]), .ZN(
        SubCellInst3_LFInst_14_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst3_LFInst_14_LFInst_2_U7  ( .A1(
        SubCellInst3_LFInst_14_LFInst_2_n18 ), .A2(
        SubCellInst3_LFInst_14_LFInst_2_n17 ), .ZN(
        SubCellInst3_LFInst_14_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst3_LFInst_14_LFInst_2_U6  ( .A(
        SubCellInst3_LFInst_14_LFInst_2_n16 ), .B(SubCellInput2[58]), .Z(
        SubCellInst3_LFInst_14_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst3_LFInst_14_LFInst_2_U5  ( .A1(SubCellInput2[56]), .A2(
        SubCellInput2[57]), .ZN(SubCellInst3_LFInst_14_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst3_LFInst_14_LFInst_2_U4  ( .A1(
        SubCellInst3_LFInst_14_LFInst_2_n15 ), .A2(SubCellInput2[59]), .ZN(
        SubCellInst3_LFInst_14_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst3_LFInst_14_LFInst_2_U3  ( .A(SubCellInput2[56]), .B(
        SubCellInput2[57]), .ZN(SubCellInst3_LFInst_14_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst3_LFInst_14_LFInst_3_U9  ( .A1(
        SubCellInst3_LFInst_14_LFInst_3_n16 ), .A2(
        SubCellInst3_LFInst_14_LFInst_3_n15 ), .ZN(MCInst3_MC1_v0_3 [0]) );
  NAND2_X1 SubCellInst3_LFInst_14_LFInst_3_U8  ( .A1(SubCellInput2[57]), .A2(
        SubCellInst3_LFInst_14_LFInst_3_n14 ), .ZN(
        SubCellInst3_LFInst_14_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst3_LFInst_14_LFInst_3_U7  ( .A(SubCellInput2[59]), .B(
        SubCellInput2[58]), .Z(SubCellInst3_LFInst_14_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst3_LFInst_14_LFInst_3_U6  ( .A1(
        SubCellInst3_LFInst_14_LFInst_3_n13 ), .A2(
        SubCellInst3_LFInst_14_LFInst_3_n12 ), .ZN(
        SubCellInst3_LFInst_14_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst3_LFInst_14_LFInst_3_U5  ( .A1(SubCellInput2[56]), .A2(
        SubCellInput2[58]), .ZN(SubCellInst3_LFInst_14_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst3_LFInst_14_LFInst_3_U4  ( .A(SubCellInput2[56]), .B(
        SubCellInst3_LFInst_14_LFInst_3_n11 ), .ZN(
        SubCellInst3_LFInst_14_LFInst_3_n13 ) );
  OR2_X1 SubCellInst3_LFInst_14_LFInst_3_U3  ( .A1(SubCellInput2[59]), .A2(
        SubCellInput2[57]), .ZN(SubCellInst3_LFInst_14_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst3_LFInst_15_LFInst_0_U6  ( .A1(SubCellInput2[62]), .A2(
        SubCellInst3_LFInst_15_LFInst_0_n4 ), .ZN(
        SubCellInst3_LFInst_15_LFInst_0_n5 ) );
  INV_X1 SubCellInst3_LFInst_15_LFInst_0_U5  ( .A(SubCellInput2[61]), .ZN(
        SubCellInst3_LFInst_15_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst3_LFInst_15_LFInst_0_U4  ( .A(SubCellInput2[60]), .B(
        SubCellInput2[63]), .Z(SubCellInst3_LFInst_15_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst3_LFInst_15_LFInst_0_U3  ( .A(
        SubCellInst3_LFInst_15_LFInst_0_n6 ), .B(
        SubCellInst3_LFInst_15_LFInst_0_n5 ), .ZN(Red_MCInst3_MC0_v0_1[0] )
         );
  NAND2_X1 SubCellInst3_LFInst_15_LFInst_1_U12  ( .A1(
        SubCellInst3_LFInst_15_LFInst_1_n18 ), .A2(
        SubCellInst3_LFInst_15_LFInst_1_n17 ), .ZN(MCInst3_MC0_v0_0 [3]) );
  NAND2_X1 SubCellInst3_LFInst_15_LFInst_1_U11  ( .A1(SubCellInput2[61]), 
        .A2(SubCellInst3_LFInst_15_LFInst_1_n16 ), .ZN(
        SubCellInst3_LFInst_15_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst3_LFInst_15_LFInst_1_U10  ( .A1(SubCellInput2[63]), .A2(
        SubCellInst3_LFInst_15_LFInst_1_n15 ), .ZN(
        SubCellInst3_LFInst_15_LFInst_1_n16 ) );
  AND2_X1 SubCellInst3_LFInst_15_LFInst_1_U9  ( .A1(SubCellInput2[60]), .A2(
        SubCellInput2[62]), .ZN(SubCellInst3_LFInst_15_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst3_LFInst_15_LFInst_1_U8  ( .A1(SubCellInput2[63]), .A2(
        SubCellInst3_LFInst_15_LFInst_1_n14 ), .ZN(
        SubCellInst3_LFInst_15_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst3_LFInst_15_LFInst_1_U7  ( .A1(
        SubCellInst3_LFInst_15_LFInst_1_n13 ), .A2(
        SubCellInst3_LFInst_15_LFInst_1_n12 ), .ZN(
        SubCellInst3_LFInst_15_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst3_LFInst_15_LFInst_1_U6  ( .A1(SubCellInput2[60]), .A2(
        SubCellInput2[62]), .ZN(SubCellInst3_LFInst_15_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst3_LFInst_15_LFInst_1_U5  ( .A1(
        SubCellInst3_LFInst_15_LFInst_1_n11 ), .A2(
        SubCellInst3_LFInst_15_LFInst_1_n10 ), .ZN(
        SubCellInst3_LFInst_15_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst3_LFInst_15_LFInst_1_U4  ( .A1(SubCellInput2[60]), .A2(
        SubCellInput2[61]), .ZN(SubCellInst3_LFInst_15_LFInst_1_n10 ) );
  INV_X1 SubCellInst3_LFInst_15_LFInst_1_U3  ( .A(SubCellInput2[62]), .ZN(
        SubCellInst3_LFInst_15_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst3_LFInst_15_LFInst_2_U11  ( .A1(
        SubCellInst3_LFInst_15_LFInst_2_n22 ), .A2(
        SubCellInst3_LFInst_15_LFInst_2_n21 ), .ZN(MCInst3_MC0_v0_3 [3]) );
  NAND2_X1 SubCellInst3_LFInst_15_LFInst_2_U10  ( .A1(SubCellInput2[62]), 
        .A2(SubCellInst3_LFInst_15_LFInst_2_n20 ), .ZN(
        SubCellInst3_LFInst_15_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst3_LFInst_15_LFInst_2_U9  ( .A1(SubCellInput2[61]), .A2(
        SubCellInst3_LFInst_15_LFInst_2_n19 ), .ZN(
        SubCellInst3_LFInst_15_LFInst_2_n20 ) );
  INV_X1 SubCellInst3_LFInst_15_LFInst_2_U8  ( .A(SubCellInput2[63]), .ZN(
        SubCellInst3_LFInst_15_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst3_LFInst_15_LFInst_2_U7  ( .A1(
        SubCellInst3_LFInst_15_LFInst_2_n18 ), .A2(
        SubCellInst3_LFInst_15_LFInst_2_n17 ), .ZN(
        SubCellInst3_LFInst_15_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst3_LFInst_15_LFInst_2_U6  ( .A(
        SubCellInst3_LFInst_15_LFInst_2_n16 ), .B(SubCellInput2[62]), .Z(
        SubCellInst3_LFInst_15_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst3_LFInst_15_LFInst_2_U5  ( .A1(SubCellInput2[60]), .A2(
        SubCellInput2[61]), .ZN(SubCellInst3_LFInst_15_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst3_LFInst_15_LFInst_2_U4  ( .A1(
        SubCellInst3_LFInst_15_LFInst_2_n15 ), .A2(SubCellInput2[63]), .ZN(
        SubCellInst3_LFInst_15_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst3_LFInst_15_LFInst_2_U3  ( .A(SubCellInput2[60]), .B(
        SubCellInput2[61]), .ZN(SubCellInst3_LFInst_15_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst3_LFInst_15_LFInst_3_U9  ( .A1(
        SubCellInst3_LFInst_15_LFInst_3_n16 ), .A2(
        SubCellInst3_LFInst_15_LFInst_3_n15 ), .ZN(MCInst3_MC0_v0_3 [0]) );
  NAND2_X1 SubCellInst3_LFInst_15_LFInst_3_U8  ( .A1(SubCellInput2[61]), .A2(
        SubCellInst3_LFInst_15_LFInst_3_n14 ), .ZN(
        SubCellInst3_LFInst_15_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst3_LFInst_15_LFInst_3_U7  ( .A(SubCellInput2[63]), .B(
        SubCellInput2[62]), .Z(SubCellInst3_LFInst_15_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst3_LFInst_15_LFInst_3_U6  ( .A1(
        SubCellInst3_LFInst_15_LFInst_3_n13 ), .A2(
        SubCellInst3_LFInst_15_LFInst_3_n12 ), .ZN(
        SubCellInst3_LFInst_15_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst3_LFInst_15_LFInst_3_U5  ( .A1(SubCellInput2[60]), .A2(
        SubCellInput2[62]), .ZN(SubCellInst3_LFInst_15_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst3_LFInst_15_LFInst_3_U4  ( .A(SubCellInput2[60]), .B(
        SubCellInst3_LFInst_15_LFInst_3_n11 ), .ZN(
        SubCellInst3_LFInst_15_LFInst_3_n13 ) );
  OR2_X1 SubCellInst3_LFInst_15_LFInst_3_U3  ( .A1(SubCellInput2[63]), .A2(
        SubCellInput2[61]), .ZN(SubCellInst3_LFInst_15_LFInst_3_n11 ) );
  XNOR2_X1 MCInst3_MC0_v0_2Inst_0_U4  ( .A(MCInst3_MC0_v0_2Inst_0_n2 ), .B(
        MCInst3_MC0_v0_0 [3]), .ZN(MCInst3_MC0_v0_2 [0]) );
  XNOR2_X1 MCInst3_MC0_v0_2Inst_0_U3  ( .A(MCInst3_MC0_v0_3 [0]), .B(
        Red_MCInst3_MC0_v0_1[0] ), .ZN(MCInst3_MC0_v0_2Inst_0_n2 ) );
  XOR2_X1 MCInst3_MC0_v1_1Inst_0_U3  ( .A(Red_MCInst3_MC0_v1_1[0] ), .B(
        MCInst3_MC0_v1_0 [3]), .Z(MCInst3_MC0_v1_1 [0]) );
  XNOR2_X1 MCInst3_MC0_v1_2Inst_0_U4  ( .A(MCInst3_MC0_v1_2Inst_0_n2 ), .B(
        Red_MCInst3_MC0_v1_1[0] ), .ZN(MCInst3_MC0_v1_2 [0]) );
  XNOR2_X1 MCInst3_MC0_v1_2Inst_0_U3  ( .A(MCInst3_MC0_v1_0 [3]), .B(
        MCInst3_MC0_v1_3 [2]), .ZN(MCInst3_MC0_v1_2Inst_0_n2 ) );
  XOR2_X1 MCInst3_MC0_v2_1Inst_0_U3  ( .A(MCInst3_MC0_v2_3 [1]), .B(
        MCInst3_MC0_v2_0 [3]), .Z(MCInst3_MC0_v2_1 [0]) );
  XOR2_X1 MCInst3_MC0_v2_2Inst_0_U3  ( .A(MCInst3_MC0_v2_0 [2]), .B(
        MCInst3_MC0_v2_0 [0]), .Z(MCInst3_MC0_v2_2 [0]) );
  XNOR2_X1 MCInst3_MC0_v2_3Inst_0_U5  ( .A(MCInst3_MC0_v2_3Inst_0_n4 ), .B(
        MCInst3_MC0_v2_3Inst_0_n3 ), .ZN(MCInst3_MC0_v2_3 [0]) );
  XNOR2_X1 MCInst3_MC0_v2_3Inst_0_U4  ( .A(MCInst3_MC0_v2_0 [2]), .B(
        MCInst3_MC0_v2_3 [1]), .ZN(MCInst3_MC0_v2_3Inst_0_n3 ) );
  XOR2_X1 MCInst3_MC0_v2_3Inst_0_U3  ( .A(MCInst3_MC0_v2_0 [3]), .B(
        MCInst3_MC0_v2_0 [0]), .Z(MCInst3_MC0_v2_3Inst_0_n4 ) );
  XOR2_X1 MCInst3_MC0_v3_1Inst_0_U3  ( .A(Red_MCInst3_MC0_v3_1[0] ), .B(
        MCInst3_MC0_v3_2 [2]), .Z(MCInst3_MC0_v3_1 [0]) );
  XOR2_X1 MCInst3_MC0_v3_2Inst_0_U3  ( .A(MCInst3_MC0_v3_2 [3]), .B(
        MCInst3_MC0_v3_0 [2]), .Z(MCInst3_MC0_v3_2 [0]) );
  XNOR2_X1 MCInst3_MC0_v3_3Inst_0_U4  ( .A(MCInst3_MC0_v3_3Inst_0_n2 ), .B(
        MCInst3_MC0_v3_0 [2]), .ZN(MCInst3_MC0_v3_3 [0]) );
  XNOR2_X1 MCInst3_MC0_v3_3Inst_0_U3  ( .A(MCInst3_MC0_v3_2 [2]), .B(
        MCInst3_MC0_v3_2 [3]), .ZN(MCInst3_MC0_v3_3Inst_0_n2 ) );
  XOR2_X1 MCInst3_MC0_v0_0Inst_1_U3  ( .A(MCInst3_MC0_v0_3 [3]), .B(
        MCInst3_MC0_v0_3 [0]), .Z(MCInst3_MC0_v0_0 [1]) );
  XOR2_X1 MCInst3_MC0_v0_1Inst_1_U3  ( .A(MCInst3_MC0_v0_0 [3]), .B(
        MCInst3_MC0_v0_3 [3]), .Z(MCInst3_MC0_v0_1 [1]) );
  XNOR2_X1 MCInst3_MC0_v0_2Inst_1_U4  ( .A(MCInst3_MC0_v0_2Inst_1_n2 ), .B(
        MCInst3_MC0_v0_3 [3]), .ZN(MCInst3_MC0_v0_2 [1]) );
  XNOR2_X1 MCInst3_MC0_v0_2Inst_1_U3  ( .A(MCInst3_MC0_v0_3 [0]), .B(
        Red_MCInst3_MC0_v0_1[0] ), .ZN(MCInst3_MC0_v0_2Inst_1_n2 ) );
  XOR2_X1 MCInst3_MC0_v0_3Inst_1_U3  ( .A(Red_MCInst3_MC0_v0_1[0] ), .B(
        MCInst3_MC0_v0_3 [0]), .Z(MCInst3_MC0_v0_3 [1]) );
  XOR2_X1 MCInst3_MC0_v1_1Inst_1_U3  ( .A(MCInst3_MC0_v1_0 [0]), .B(
        Red_MCInst3_MC0_v1_1[0] ), .Z(MCInst3_MC0_v1_1 [1]) );
  XOR2_X1 MCInst3_MC0_v1_2Inst_1_U3  ( .A(MCInst3_MC0_v1_0 [0]), .B(
        MCInst3_MC0_v1_3 [2]), .Z(MCInst3_MC0_v1_2 [1]) );
  XOR2_X1 MCInst3_MC0_v1_3Inst_1_U3  ( .A(MCInst3_MC0_v1_0 [0]), .B(
        MCInst3_MC0_v1_0 [3]), .Z(MCInst3_MC0_v1_3 [1]) );
  XOR2_X1 MCInst3_MC0_v2_0Inst_1_U3  ( .A(MCInst3_MC0_v2_3 [1]), .B(
        MCInst3_MC0_v2_0 [0]), .Z(MCInst3_MC0_v2_0 [1]) );
  XNOR2_X1 MCInst3_MC0_v2_1Inst_1_U4  ( .A(MCInst3_MC0_v2_1Inst_1_n2 ), .B(
        MCInst3_MC0_v2_0 [3]), .ZN(MCInst3_MC0_v2_1 [1]) );
  XNOR2_X1 MCInst3_MC0_v2_1Inst_1_U3  ( .A(MCInst3_MC0_v2_0 [0]), .B(
        MCInst3_MC0_v2_0 [2]), .ZN(MCInst3_MC0_v2_1Inst_1_n2 ) );
  XNOR2_X1 MCInst3_MC0_v2_2Inst_1_U5  ( .A(MCInst3_MC0_v2_2Inst_1_n4 ), .B(
        MCInst3_MC0_v2_2Inst_1_n3 ), .ZN(MCInst3_MC0_v2_2 [1]) );
  XNOR2_X1 MCInst3_MC0_v2_2Inst_1_U4  ( .A(MCInst3_MC0_v2_0 [2]), .B(
        MCInst3_MC0_v2_3 [1]), .ZN(MCInst3_MC0_v2_2Inst_1_n3 ) );
  XOR2_X1 MCInst3_MC0_v2_2Inst_1_U3  ( .A(MCInst3_MC0_v2_0 [3]), .B(
        MCInst3_MC0_v2_0 [0]), .Z(MCInst3_MC0_v2_2Inst_1_n4 ) );
  XOR2_X1 MCInst3_MC0_v3_0Inst_1_U3  ( .A(MCInst3_MC0_v3_2 [3]), .B(
        MCInst3_MC0_v3_2 [2]), .Z(MCInst3_MC0_v3_0 [1]) );
  XOR2_X1 MCInst3_MC0_v3_1Inst_1_U3  ( .A(MCInst3_MC0_v3_2 [3]), .B(
        Red_MCInst3_MC0_v3_1[0] ), .Z(MCInst3_MC0_v3_1 [1]) );
  XNOR2_X1 MCInst3_MC0_v3_3Inst_1_U4  ( .A(MCInst3_MC0_v3_3Inst_1_n2 ), .B(
        Red_MCInst3_MC0_v3_1[0] ), .ZN(MCInst3_MC0_v3_3 [1]) );
  XNOR2_X1 MCInst3_MC0_v3_3Inst_1_U3  ( .A(MCInst3_MC0_v3_2 [2]), .B(
        MCInst3_MC0_v3_2 [3]), .ZN(MCInst3_MC0_v3_3Inst_1_n2 ) );
  XOR2_X1 MCInst3_MC0_v0_0Inst_2_U3  ( .A(Red_MCInst3_MC0_v0_1[0] ), .B(
        MCInst3_MC0_v0_3 [0]), .Z(MCInst3_MC0_v0_0 [2]) );
  XOR2_X1 MCInst3_MC0_v0_1Inst_2_U3  ( .A(MCInst3_MC0_v0_3 [3]), .B(
        MCInst3_MC0_v0_3 [0]), .Z(MCInst3_MC0_v0_1 [2]) );
  XOR2_X1 MCInst3_MC0_v0_2Inst_2_U3  ( .A(MCInst3_MC0_v0_0 [3]), .B(
        MCInst3_MC0_v0_3 [0]), .Z(MCInst3_MC0_v0_2 [2]) );
  XNOR2_X1 MCInst3_MC0_v1_1Inst_2_U4  ( .A(MCInst3_MC0_v1_1Inst_2_n2 ), .B(
        MCInst3_MC0_v1_3 [2]), .ZN(MCInst3_MC0_v1_1 [2]) );
  XNOR2_X1 MCInst3_MC0_v1_1Inst_2_U3  ( .A(MCInst3_MC0_v1_0 [3]), .B(
        MCInst3_MC0_v1_0 [0]), .ZN(MCInst3_MC0_v1_1Inst_2_n2 ) );
  XNOR2_X1 MCInst3_MC0_v1_2Inst_2_U4  ( .A(MCInst3_MC0_v1_2Inst_2_n2 ), .B(
        MCInst3_MC0_v1_3 [2]), .ZN(MCInst3_MC0_v1_2 [2]) );
  XNOR2_X1 MCInst3_MC0_v1_2Inst_2_U3  ( .A(Red_MCInst3_MC0_v1_1[0] ), .B(
        MCInst3_MC0_v1_0 [0]), .ZN(MCInst3_MC0_v1_2Inst_2_n2 ) );
  XNOR2_X1 MCInst3_MC0_v2_1Inst_2_U4  ( .A(MCInst3_MC0_v2_1Inst_2_n2 ), .B(
        MCInst3_MC0_v2_0 [3]), .ZN(MCInst3_MC0_v2_1 [2]) );
  XNOR2_X1 MCInst3_MC0_v2_1Inst_2_U3  ( .A(MCInst3_MC0_v2_0 [0]), .B(
        MCInst3_MC0_v2_3 [1]), .ZN(MCInst3_MC0_v2_1Inst_2_n2 ) );
  XNOR2_X1 MCInst3_MC0_v2_2Inst_2_U4  ( .A(MCInst3_MC0_v2_2Inst_2_n2 ), .B(
        MCInst3_MC0_v2_0 [3]), .ZN(MCInst3_MC0_v2_2 [2]) );
  XNOR2_X1 MCInst3_MC0_v2_2Inst_2_U3  ( .A(MCInst3_MC0_v2_0 [0]), .B(
        MCInst3_MC0_v2_0 [2]), .ZN(MCInst3_MC0_v2_2Inst_2_n2 ) );
  XOR2_X1 MCInst3_MC0_v2_3Inst_2_U3  ( .A(MCInst3_MC0_v2_3 [1]), .B(
        MCInst3_MC0_v2_0 [2]), .Z(MCInst3_MC0_v2_3 [2]) );
  XNOR2_X1 MCInst3_MC0_v3_1Inst_2_U4  ( .A(MCInst3_MC0_v3_1Inst_2_n2 ), .B(
        MCInst3_MC0_v3_0 [2]), .ZN(MCInst3_MC0_v3_1 [2]) );
  XNOR2_X1 MCInst3_MC0_v3_1Inst_2_U3  ( .A(MCInst3_MC0_v3_2 [2]), .B(
        MCInst3_MC0_v3_2 [3]), .ZN(MCInst3_MC0_v3_1Inst_2_n2 ) );
  XOR2_X1 MCInst3_MC0_v3_3Inst_2_U3  ( .A(MCInst3_MC0_v3_0 [2]), .B(
        MCInst3_MC0_v3_2 [2]), .Z(MCInst3_MC0_v3_3 [2]) );
  XOR2_X1 MCInst3_MC0_v0_1Inst_3_U3  ( .A(Red_MCInst3_MC0_v0_1[0] ), .B(
        MCInst3_MC0_v0_3 [0]), .Z(MCInst3_MC0_v0_1 [3]) );
  XOR2_X1 MCInst3_MC0_v0_2Inst_3_U3  ( .A(Red_MCInst3_MC0_v0_1[0] ), .B(
        MCInst3_MC0_v0_3 [3]), .Z(MCInst3_MC0_v0_2 [3]) );
  XOR2_X1 MCInst3_MC0_v1_1Inst_3_U3  ( .A(MCInst3_MC0_v1_3 [2]), .B(
        Red_MCInst3_MC0_v1_1[0] ), .Z(MCInst3_MC0_v1_1 [3]) );
  XNOR2_X1 MCInst3_MC0_v1_2Inst_3_U5  ( .A(MCInst3_MC0_v1_2Inst_3_n4 ), .B(
        MCInst3_MC0_v1_2Inst_3_n3 ), .ZN(MCInst3_MC0_v1_2 [3]) );
  XNOR2_X1 MCInst3_MC0_v1_2Inst_3_U4  ( .A(MCInst3_MC0_v1_3 [2]), .B(
        MCInst3_MC0_v1_0 [0]), .ZN(MCInst3_MC0_v1_2Inst_3_n3 ) );
  XOR2_X1 MCInst3_MC0_v1_2Inst_3_U3  ( .A(Red_MCInst3_MC0_v1_1[0] ), .B(
        MCInst3_MC0_v1_0 [3]), .Z(MCInst3_MC0_v1_2Inst_3_n4 ) );
  XOR2_X1 MCInst3_MC0_v2_1Inst_3_U3  ( .A(MCInst3_MC0_v2_0 [2]), .B(
        MCInst3_MC0_v2_0 [0]), .Z(MCInst3_MC0_v2_1 [3]) );
  XNOR2_X1 MCInst3_MC0_v2_2Inst_3_U4  ( .A(MCInst3_MC0_v2_2Inst_3_n2 ), .B(
        MCInst3_MC0_v2_0 [3]), .ZN(MCInst3_MC0_v2_2 [3]) );
  XNOR2_X1 MCInst3_MC0_v2_2Inst_3_U3  ( .A(MCInst3_MC0_v2_0 [0]), .B(
        MCInst3_MC0_v2_3 [1]), .ZN(MCInst3_MC0_v2_2Inst_3_n2 ) );
  XNOR2_X1 MCInst3_MC0_v2_3Inst_3_U4  ( .A(MCInst3_MC0_v2_3Inst_3_n2 ), .B(
        MCInst3_MC0_v2_0 [2]), .ZN(MCInst3_MC0_v2_3 [3]) );
  XNOR2_X1 MCInst3_MC0_v2_3Inst_3_U3  ( .A(MCInst3_MC0_v2_0 [3]), .B(
        MCInst3_MC0_v2_3 [1]), .ZN(MCInst3_MC0_v2_3Inst_3_n2 ) );
  XOR2_X1 MCInst3_MC0_v3_1Inst_3_U3  ( .A(MCInst3_MC0_v3_0 [2]), .B(
        Red_MCInst3_MC0_v3_1[0] ), .Z(MCInst3_MC0_v3_1 [3]) );
  XOR2_X1 MCInst3_MC0_v3_3Inst_3_U3  ( .A(MCInst3_MC0_v3_2 [3]), .B(
        Red_MCInst3_MC0_v3_1[0] ), .Z(MCInst3_MC0_v3_3 [3]) );
  XNOR2_X1 MCInst3_MC0_r0Inst_XORInst_0_0_U3  ( .A(
        MCInst3_MC0_r0Inst_XORInst_0_0_n5 ), .B(
        MCInst3_MC0_r0Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[60]) );
  XNOR2_X1 MCInst3_MC0_r0Inst_XORInst_0_0_U2  ( .A(MCInst3_MC0_v3_2 [2]), 
        .B(MCInst3_MC0_v2_0 [0]), .ZN(MCInst3_MC0_r0Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst3_MC0_r0Inst_XORInst_0_0_U1  ( .A(MCInst3_MC0_v0_3 [3]), .B(
        MCInst3_MC0_v1_0 [0]), .Z(MCInst3_MC0_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst3_MC0_r0Inst_XORInst_0_1_U3  ( .A(
        MCInst3_MC0_r0Inst_XORInst_0_1_n5 ), .B(
        MCInst3_MC0_r0Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[61]) );
  XNOR2_X1 MCInst3_MC0_r0Inst_XORInst_0_1_U2  ( .A(MCInst3_MC0_v3_0 [1]), 
        .B(MCInst3_MC0_v2_0 [1]), .ZN(MCInst3_MC0_r0Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst3_MC0_r0Inst_XORInst_0_1_U1  ( .A(MCInst3_MC0_v0_0 [1]), .B(
        MCInst3_MC0_v1_3 [2]), .Z(MCInst3_MC0_r0Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst3_MC0_r0Inst_XORInst_0_2_U3  ( .A(
        MCInst3_MC0_r0Inst_XORInst_0_2_n5 ), .B(
        MCInst3_MC0_r0Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[62]) );
  XNOR2_X1 MCInst3_MC0_r0Inst_XORInst_0_2_U2  ( .A(MCInst3_MC0_v3_0 [2]), 
        .B(MCInst3_MC0_v2_0 [2]), .ZN(MCInst3_MC0_r0Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst3_MC0_r0Inst_XORInst_0_2_U1  ( .A(MCInst3_MC0_v0_0 [2]), .B(
        Red_MCInst3_MC0_v1_1[0] ), .Z(MCInst3_MC0_r0Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst3_MC0_r0Inst_XORInst_0_3_U3  ( .A(
        MCInst3_MC0_r0Inst_XORInst_0_3_n5 ), .B(
        MCInst3_MC0_r0Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[63]) );
  XNOR2_X1 MCInst3_MC0_r0Inst_XORInst_0_3_U2  ( .A(Red_MCInst3_MC0_v3_1[0] ), 
        .B(MCInst3_MC0_v2_0 [3]), .ZN(MCInst3_MC0_r0Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst3_MC0_r0Inst_XORInst_0_3_U1  ( .A(MCInst3_MC0_v0_0 [3]), .B(
        MCInst3_MC0_v1_0 [3]), .Z(MCInst3_MC0_r0Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst3_MC0_r1Inst_XORInst_0_0_U3  ( .A(
        MCInst3_MC0_r1Inst_XORInst_0_0_n5 ), .B(
        MCInst3_MC0_r1Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[44]) );
  XNOR2_X1 MCInst3_MC0_r1Inst_XORInst_0_0_U2  ( .A(MCInst3_MC0_v3_1 [0]), 
        .B(MCInst3_MC0_v2_1 [0]), .ZN(MCInst3_MC0_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst3_MC0_r1Inst_XORInst_0_0_U1  ( .A(MCInst3_MC0_v0_0 [3]), .B(
        MCInst3_MC0_v1_1 [0]), .Z(MCInst3_MC0_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst3_MC0_r1Inst_XORInst_0_1_U3  ( .A(
        MCInst3_MC0_r1Inst_XORInst_0_1_n5 ), .B(
        MCInst3_MC0_r1Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[45]) );
  XNOR2_X1 MCInst3_MC0_r1Inst_XORInst_0_1_U2  ( .A(MCInst3_MC0_v3_1 [1]), 
        .B(MCInst3_MC0_v2_1 [1]), .ZN(MCInst3_MC0_r1Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst3_MC0_r1Inst_XORInst_0_1_U1  ( .A(MCInst3_MC0_v0_1 [1]), .B(
        MCInst3_MC0_v1_1 [1]), .Z(MCInst3_MC0_r1Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst3_MC0_r1Inst_XORInst_0_2_U3  ( .A(
        MCInst3_MC0_r1Inst_XORInst_0_2_n5 ), .B(
        MCInst3_MC0_r1Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[46]) );
  XNOR2_X1 MCInst3_MC0_r1Inst_XORInst_0_2_U2  ( .A(MCInst3_MC0_v3_1 [2]), 
        .B(MCInst3_MC0_v2_1 [2]), .ZN(MCInst3_MC0_r1Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst3_MC0_r1Inst_XORInst_0_2_U1  ( .A(MCInst3_MC0_v0_1 [2]), .B(
        MCInst3_MC0_v1_1 [2]), .Z(MCInst3_MC0_r1Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst3_MC0_r1Inst_XORInst_0_3_U3  ( .A(
        MCInst3_MC0_r1Inst_XORInst_0_3_n5 ), .B(
        MCInst3_MC0_r1Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[47]) );
  XNOR2_X1 MCInst3_MC0_r1Inst_XORInst_0_3_U2  ( .A(MCInst3_MC0_v3_1 [3]), 
        .B(MCInst3_MC0_v2_1 [3]), .ZN(MCInst3_MC0_r1Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst3_MC0_r1Inst_XORInst_0_3_U1  ( .A(MCInst3_MC0_v0_1 [3]), .B(
        MCInst3_MC0_v1_1 [3]), .Z(MCInst3_MC0_r1Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst3_MC0_r2Inst_XORInst_0_0_U3  ( .A(
        MCInst3_MC0_r2Inst_XORInst_0_0_n5 ), .B(
        MCInst3_MC0_r2Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[28]) );
  XNOR2_X1 MCInst3_MC0_r2Inst_XORInst_0_0_U2  ( .A(MCInst3_MC0_v3_2 [0]), 
        .B(MCInst3_MC0_v2_2 [0]), .ZN(MCInst3_MC0_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst3_MC0_r2Inst_XORInst_0_0_U1  ( .A(MCInst3_MC0_v0_2 [0]), .B(
        MCInst3_MC0_v1_2 [0]), .Z(MCInst3_MC0_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst3_MC0_r2Inst_XORInst_0_1_U3  ( .A(
        MCInst3_MC0_r2Inst_XORInst_0_1_n5 ), .B(
        MCInst3_MC0_r2Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[29]) );
  XNOR2_X1 MCInst3_MC0_r2Inst_XORInst_0_1_U2  ( .A(Red_MCInst3_MC0_v3_1[0] ), 
        .B(MCInst3_MC0_v2_2 [1]), .ZN(MCInst3_MC0_r2Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst3_MC0_r2Inst_XORInst_0_1_U1  ( .A(MCInst3_MC0_v0_2 [1]), .B(
        MCInst3_MC0_v1_2 [1]), .Z(MCInst3_MC0_r2Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst3_MC0_r2Inst_XORInst_0_2_U3  ( .A(
        MCInst3_MC0_r2Inst_XORInst_0_2_n5 ), .B(
        MCInst3_MC0_r2Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[30]) );
  XNOR2_X1 MCInst3_MC0_r2Inst_XORInst_0_2_U2  ( .A(MCInst3_MC0_v3_2 [2]), 
        .B(MCInst3_MC0_v2_2 [2]), .ZN(MCInst3_MC0_r2Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst3_MC0_r2Inst_XORInst_0_2_U1  ( .A(MCInst3_MC0_v0_2 [2]), .B(
        MCInst3_MC0_v1_2 [2]), .Z(MCInst3_MC0_r2Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst3_MC0_r2Inst_XORInst_0_3_U3  ( .A(
        MCInst3_MC0_r2Inst_XORInst_0_3_n5 ), .B(
        MCInst3_MC0_r2Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[31]) );
  XNOR2_X1 MCInst3_MC0_r2Inst_XORInst_0_3_U2  ( .A(MCInst3_MC0_v3_2 [3]), 
        .B(MCInst3_MC0_v2_2 [3]), .ZN(MCInst3_MC0_r2Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst3_MC0_r2Inst_XORInst_0_3_U1  ( .A(MCInst3_MC0_v0_2 [3]), .B(
        MCInst3_MC0_v1_2 [3]), .Z(MCInst3_MC0_r2Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst3_MC0_r3Inst_XORInst_0_0_U3  ( .A(
        MCInst3_MC0_r3Inst_XORInst_0_0_n5 ), .B(
        MCInst3_MC0_r3Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[12]) );
  XNOR2_X1 MCInst3_MC0_r3Inst_XORInst_0_0_U2  ( .A(MCInst3_MC0_v3_3 [0]), 
        .B(MCInst3_MC0_v2_3 [0]), .ZN(MCInst3_MC0_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst3_MC0_r3Inst_XORInst_0_0_U1  ( .A(MCInst3_MC0_v0_3 [0]), .B(
        MCInst3_MC0_v1_0 [3]), .Z(MCInst3_MC0_r3Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst3_MC0_r3Inst_XORInst_0_1_U3  ( .A(
        MCInst3_MC0_r3Inst_XORInst_0_1_n5 ), .B(
        MCInst3_MC0_r3Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[13]) );
  XNOR2_X1 MCInst3_MC0_r3Inst_XORInst_0_1_U2  ( .A(MCInst3_MC0_v3_3 [1]), 
        .B(MCInst3_MC0_v2_3 [1]), .ZN(MCInst3_MC0_r3Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst3_MC0_r3Inst_XORInst_0_1_U1  ( .A(MCInst3_MC0_v0_3 [1]), .B(
        MCInst3_MC0_v1_3 [1]), .Z(MCInst3_MC0_r3Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst3_MC0_r3Inst_XORInst_0_2_U3  ( .A(
        MCInst3_MC0_r3Inst_XORInst_0_2_n5 ), .B(
        MCInst3_MC0_r3Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[14]) );
  XNOR2_X1 MCInst3_MC0_r3Inst_XORInst_0_2_U2  ( .A(MCInst3_MC0_v3_3 [2]), 
        .B(MCInst3_MC0_v2_3 [2]), .ZN(MCInst3_MC0_r3Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst3_MC0_r3Inst_XORInst_0_2_U1  ( .A(MCInst3_MC0_v0_0 [3]), .B(
        MCInst3_MC0_v1_3 [2]), .Z(MCInst3_MC0_r3Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst3_MC0_r3Inst_XORInst_0_3_U3  ( .A(
        MCInst3_MC0_r3Inst_XORInst_0_3_n5 ), .B(
        MCInst3_MC0_r3Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[15]) );
  XNOR2_X1 MCInst3_MC0_r3Inst_XORInst_0_3_U2  ( .A(MCInst3_MC0_v3_3 [3]), 
        .B(MCInst3_MC0_v2_3 [3]), .ZN(MCInst3_MC0_r3Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst3_MC0_r3Inst_XORInst_0_3_U1  ( .A(MCInst3_MC0_v0_3 [3]), .B(
        Red_MCInst3_MC0_v1_1[0] ), .Z(MCInst3_MC0_r3Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst3_MC1_v0_2Inst_0_U4  ( .A(MCInst3_MC1_v0_2Inst_0_n2 ), .B(
        MCInst3_MC1_v0_0 [3]), .ZN(MCInst3_MC1_v0_2 [0]) );
  XNOR2_X1 MCInst3_MC1_v0_2Inst_0_U3  ( .A(MCInst3_MC1_v0_3 [0]), .B(
        Red_MCInst3_MC1_v0_1[0] ), .ZN(MCInst3_MC1_v0_2Inst_0_n2 ) );
  XOR2_X1 MCInst3_MC1_v1_1Inst_0_U3  ( .A(Red_MCInst3_MC1_v1_1[0] ), .B(
        MCInst3_MC1_v1_0 [3]), .Z(MCInst3_MC1_v1_1 [0]) );
  XNOR2_X1 MCInst3_MC1_v1_2Inst_0_U4  ( .A(MCInst3_MC1_v1_2Inst_0_n2 ), .B(
        Red_MCInst3_MC1_v1_1[0] ), .ZN(MCInst3_MC1_v1_2 [0]) );
  XNOR2_X1 MCInst3_MC1_v1_2Inst_0_U3  ( .A(MCInst3_MC1_v1_0 [3]), .B(
        MCInst3_MC1_v1_3 [2]), .ZN(MCInst3_MC1_v1_2Inst_0_n2 ) );
  XOR2_X1 MCInst3_MC1_v2_1Inst_0_U3  ( .A(MCInst3_MC1_v2_3 [1]), .B(
        MCInst3_MC1_v2_0 [3]), .Z(MCInst3_MC1_v2_1 [0]) );
  XOR2_X1 MCInst3_MC1_v2_2Inst_0_U3  ( .A(MCInst3_MC1_v2_0 [2]), .B(
        MCInst3_MC1_v2_0 [0]), .Z(MCInst3_MC1_v2_2 [0]) );
  XNOR2_X1 MCInst3_MC1_v2_3Inst_0_U5  ( .A(MCInst3_MC1_v2_3Inst_0_n4 ), .B(
        MCInst3_MC1_v2_3Inst_0_n3 ), .ZN(MCInst3_MC1_v2_3 [0]) );
  XNOR2_X1 MCInst3_MC1_v2_3Inst_0_U4  ( .A(MCInst3_MC1_v2_0 [2]), .B(
        MCInst3_MC1_v2_3 [1]), .ZN(MCInst3_MC1_v2_3Inst_0_n3 ) );
  XOR2_X1 MCInst3_MC1_v2_3Inst_0_U3  ( .A(MCInst3_MC1_v2_0 [3]), .B(
        MCInst3_MC1_v2_0 [0]), .Z(MCInst3_MC1_v2_3Inst_0_n4 ) );
  XOR2_X1 MCInst3_MC1_v3_1Inst_0_U3  ( .A(Red_MCInst3_MC1_v3_1[0] ), .B(
        MCInst3_MC1_v3_2 [2]), .Z(MCInst3_MC1_v3_1 [0]) );
  XOR2_X1 MCInst3_MC1_v3_2Inst_0_U3  ( .A(MCInst3_MC1_v3_2 [3]), .B(
        MCInst3_MC1_v3_0 [2]), .Z(MCInst3_MC1_v3_2 [0]) );
  XNOR2_X1 MCInst3_MC1_v3_3Inst_0_U4  ( .A(MCInst3_MC1_v3_3Inst_0_n2 ), .B(
        MCInst3_MC1_v3_0 [2]), .ZN(MCInst3_MC1_v3_3 [0]) );
  XNOR2_X1 MCInst3_MC1_v3_3Inst_0_U3  ( .A(MCInst3_MC1_v3_2 [2]), .B(
        MCInst3_MC1_v3_2 [3]), .ZN(MCInst3_MC1_v3_3Inst_0_n2 ) );
  XOR2_X1 MCInst3_MC1_v0_0Inst_1_U3  ( .A(MCInst3_MC1_v0_3 [3]), .B(
        MCInst3_MC1_v0_3 [0]), .Z(MCInst3_MC1_v0_0 [1]) );
  XOR2_X1 MCInst3_MC1_v0_1Inst_1_U3  ( .A(MCInst3_MC1_v0_0 [3]), .B(
        MCInst3_MC1_v0_3 [3]), .Z(MCInst3_MC1_v0_1 [1]) );
  XNOR2_X1 MCInst3_MC1_v0_2Inst_1_U4  ( .A(MCInst3_MC1_v0_2Inst_1_n2 ), .B(
        MCInst3_MC1_v0_3 [3]), .ZN(MCInst3_MC1_v0_2 [1]) );
  XNOR2_X1 MCInst3_MC1_v0_2Inst_1_U3  ( .A(MCInst3_MC1_v0_3 [0]), .B(
        Red_MCInst3_MC1_v0_1[0] ), .ZN(MCInst3_MC1_v0_2Inst_1_n2 ) );
  XOR2_X1 MCInst3_MC1_v0_3Inst_1_U3  ( .A(Red_MCInst3_MC1_v0_1[0] ), .B(
        MCInst3_MC1_v0_3 [0]), .Z(MCInst3_MC1_v0_3 [1]) );
  XOR2_X1 MCInst3_MC1_v1_1Inst_1_U3  ( .A(MCInst3_MC1_v1_0 [0]), .B(
        Red_MCInst3_MC1_v1_1[0] ), .Z(MCInst3_MC1_v1_1 [1]) );
  XOR2_X1 MCInst3_MC1_v1_2Inst_1_U3  ( .A(MCInst3_MC1_v1_0 [0]), .B(
        MCInst3_MC1_v1_3 [2]), .Z(MCInst3_MC1_v1_2 [1]) );
  XOR2_X1 MCInst3_MC1_v1_3Inst_1_U3  ( .A(MCInst3_MC1_v1_0 [0]), .B(
        MCInst3_MC1_v1_0 [3]), .Z(MCInst3_MC1_v1_3 [1]) );
  XOR2_X1 MCInst3_MC1_v2_0Inst_1_U3  ( .A(MCInst3_MC1_v2_3 [1]), .B(
        MCInst3_MC1_v2_0 [0]), .Z(MCInst3_MC1_v2_0 [1]) );
  XNOR2_X1 MCInst3_MC1_v2_1Inst_1_U4  ( .A(MCInst3_MC1_v2_1Inst_1_n2 ), .B(
        MCInst3_MC1_v2_0 [3]), .ZN(MCInst3_MC1_v2_1 [1]) );
  XNOR2_X1 MCInst3_MC1_v2_1Inst_1_U3  ( .A(MCInst3_MC1_v2_0 [0]), .B(
        MCInst3_MC1_v2_0 [2]), .ZN(MCInst3_MC1_v2_1Inst_1_n2 ) );
  XNOR2_X1 MCInst3_MC1_v2_2Inst_1_U5  ( .A(MCInst3_MC1_v2_2Inst_1_n4 ), .B(
        MCInst3_MC1_v2_2Inst_1_n3 ), .ZN(MCInst3_MC1_v2_2 [1]) );
  XNOR2_X1 MCInst3_MC1_v2_2Inst_1_U4  ( .A(MCInst3_MC1_v2_0 [2]), .B(
        MCInst3_MC1_v2_3 [1]), .ZN(MCInst3_MC1_v2_2Inst_1_n3 ) );
  XOR2_X1 MCInst3_MC1_v2_2Inst_1_U3  ( .A(MCInst3_MC1_v2_0 [3]), .B(
        MCInst3_MC1_v2_0 [0]), .Z(MCInst3_MC1_v2_2Inst_1_n4 ) );
  XOR2_X1 MCInst3_MC1_v3_0Inst_1_U3  ( .A(MCInst3_MC1_v3_2 [3]), .B(
        MCInst3_MC1_v3_2 [2]), .Z(MCInst3_MC1_v3_0 [1]) );
  XOR2_X1 MCInst3_MC1_v3_1Inst_1_U3  ( .A(MCInst3_MC1_v3_2 [3]), .B(
        Red_MCInst3_MC1_v3_1[0] ), .Z(MCInst3_MC1_v3_1 [1]) );
  XNOR2_X1 MCInst3_MC1_v3_3Inst_1_U4  ( .A(MCInst3_MC1_v3_3Inst_1_n2 ), .B(
        Red_MCInst3_MC1_v3_1[0] ), .ZN(MCInst3_MC1_v3_3 [1]) );
  XNOR2_X1 MCInst3_MC1_v3_3Inst_1_U3  ( .A(MCInst3_MC1_v3_2 [2]), .B(
        MCInst3_MC1_v3_2 [3]), .ZN(MCInst3_MC1_v3_3Inst_1_n2 ) );
  XOR2_X1 MCInst3_MC1_v0_0Inst_2_U3  ( .A(Red_MCInst3_MC1_v0_1[0] ), .B(
        MCInst3_MC1_v0_3 [0]), .Z(MCInst3_MC1_v0_0 [2]) );
  XOR2_X1 MCInst3_MC1_v0_1Inst_2_U3  ( .A(MCInst3_MC1_v0_3 [3]), .B(
        MCInst3_MC1_v0_3 [0]), .Z(MCInst3_MC1_v0_1 [2]) );
  XOR2_X1 MCInst3_MC1_v0_2Inst_2_U3  ( .A(MCInst3_MC1_v0_0 [3]), .B(
        MCInst3_MC1_v0_3 [0]), .Z(MCInst3_MC1_v0_2 [2]) );
  XNOR2_X1 MCInst3_MC1_v1_1Inst_2_U4  ( .A(MCInst3_MC1_v1_1Inst_2_n2 ), .B(
        MCInst3_MC1_v1_3 [2]), .ZN(MCInst3_MC1_v1_1 [2]) );
  XNOR2_X1 MCInst3_MC1_v1_1Inst_2_U3  ( .A(MCInst3_MC1_v1_0 [3]), .B(
        MCInst3_MC1_v1_0 [0]), .ZN(MCInst3_MC1_v1_1Inst_2_n2 ) );
  XNOR2_X1 MCInst3_MC1_v1_2Inst_2_U4  ( .A(MCInst3_MC1_v1_2Inst_2_n2 ), .B(
        MCInst3_MC1_v1_3 [2]), .ZN(MCInst3_MC1_v1_2 [2]) );
  XNOR2_X1 MCInst3_MC1_v1_2Inst_2_U3  ( .A(Red_MCInst3_MC1_v1_1[0] ), .B(
        MCInst3_MC1_v1_0 [0]), .ZN(MCInst3_MC1_v1_2Inst_2_n2 ) );
  XNOR2_X1 MCInst3_MC1_v2_1Inst_2_U4  ( .A(MCInst3_MC1_v2_1Inst_2_n2 ), .B(
        MCInst3_MC1_v2_0 [3]), .ZN(MCInst3_MC1_v2_1 [2]) );
  XNOR2_X1 MCInst3_MC1_v2_1Inst_2_U3  ( .A(MCInst3_MC1_v2_0 [0]), .B(
        MCInst3_MC1_v2_3 [1]), .ZN(MCInst3_MC1_v2_1Inst_2_n2 ) );
  XNOR2_X1 MCInst3_MC1_v2_2Inst_2_U4  ( .A(MCInst3_MC1_v2_2Inst_2_n2 ), .B(
        MCInst3_MC1_v2_0 [3]), .ZN(MCInst3_MC1_v2_2 [2]) );
  XNOR2_X1 MCInst3_MC1_v2_2Inst_2_U3  ( .A(MCInst3_MC1_v2_0 [0]), .B(
        MCInst3_MC1_v2_0 [2]), .ZN(MCInst3_MC1_v2_2Inst_2_n2 ) );
  XOR2_X1 MCInst3_MC1_v2_3Inst_2_U3  ( .A(MCInst3_MC1_v2_3 [1]), .B(
        MCInst3_MC1_v2_0 [2]), .Z(MCInst3_MC1_v2_3 [2]) );
  XNOR2_X1 MCInst3_MC1_v3_1Inst_2_U4  ( .A(MCInst3_MC1_v3_1Inst_2_n2 ), .B(
        MCInst3_MC1_v3_0 [2]), .ZN(MCInst3_MC1_v3_1 [2]) );
  XNOR2_X1 MCInst3_MC1_v3_1Inst_2_U3  ( .A(MCInst3_MC1_v3_2 [2]), .B(
        MCInst3_MC1_v3_2 [3]), .ZN(MCInst3_MC1_v3_1Inst_2_n2 ) );
  XOR2_X1 MCInst3_MC1_v3_3Inst_2_U3  ( .A(MCInst3_MC1_v3_0 [2]), .B(
        MCInst3_MC1_v3_2 [2]), .Z(MCInst3_MC1_v3_3 [2]) );
  XOR2_X1 MCInst3_MC1_v0_1Inst_3_U3  ( .A(Red_MCInst3_MC1_v0_1[0] ), .B(
        MCInst3_MC1_v0_3 [0]), .Z(MCInst3_MC1_v0_1 [3]) );
  XOR2_X1 MCInst3_MC1_v0_2Inst_3_U3  ( .A(Red_MCInst3_MC1_v0_1[0] ), .B(
        MCInst3_MC1_v0_3 [3]), .Z(MCInst3_MC1_v0_2 [3]) );
  XOR2_X1 MCInst3_MC1_v1_1Inst_3_U3  ( .A(MCInst3_MC1_v1_3 [2]), .B(
        Red_MCInst3_MC1_v1_1[0] ), .Z(MCInst3_MC1_v1_1 [3]) );
  XNOR2_X1 MCInst3_MC1_v1_2Inst_3_U5  ( .A(MCInst3_MC1_v1_2Inst_3_n4 ), .B(
        MCInst3_MC1_v1_2Inst_3_n3 ), .ZN(MCInst3_MC1_v1_2 [3]) );
  XNOR2_X1 MCInst3_MC1_v1_2Inst_3_U4  ( .A(MCInst3_MC1_v1_3 [2]), .B(
        MCInst3_MC1_v1_0 [0]), .ZN(MCInst3_MC1_v1_2Inst_3_n3 ) );
  XOR2_X1 MCInst3_MC1_v1_2Inst_3_U3  ( .A(Red_MCInst3_MC1_v1_1[0] ), .B(
        MCInst3_MC1_v1_0 [3]), .Z(MCInst3_MC1_v1_2Inst_3_n4 ) );
  XOR2_X1 MCInst3_MC1_v2_1Inst_3_U3  ( .A(MCInst3_MC1_v2_0 [2]), .B(
        MCInst3_MC1_v2_0 [0]), .Z(MCInst3_MC1_v2_1 [3]) );
  XNOR2_X1 MCInst3_MC1_v2_2Inst_3_U4  ( .A(MCInst3_MC1_v2_2Inst_3_n2 ), .B(
        MCInst3_MC1_v2_0 [3]), .ZN(MCInst3_MC1_v2_2 [3]) );
  XNOR2_X1 MCInst3_MC1_v2_2Inst_3_U3  ( .A(MCInst3_MC1_v2_0 [0]), .B(
        MCInst3_MC1_v2_3 [1]), .ZN(MCInst3_MC1_v2_2Inst_3_n2 ) );
  XNOR2_X1 MCInst3_MC1_v2_3Inst_3_U4  ( .A(MCInst3_MC1_v2_3Inst_3_n2 ), .B(
        MCInst3_MC1_v2_0 [2]), .ZN(MCInst3_MC1_v2_3 [3]) );
  XNOR2_X1 MCInst3_MC1_v2_3Inst_3_U3  ( .A(MCInst3_MC1_v2_0 [3]), .B(
        MCInst3_MC1_v2_3 [1]), .ZN(MCInst3_MC1_v2_3Inst_3_n2 ) );
  XOR2_X1 MCInst3_MC1_v3_1Inst_3_U3  ( .A(MCInst3_MC1_v3_0 [2]), .B(
        Red_MCInst3_MC1_v3_1[0] ), .Z(MCInst3_MC1_v3_1 [3]) );
  XOR2_X1 MCInst3_MC1_v3_3Inst_3_U3  ( .A(MCInst3_MC1_v3_2 [3]), .B(
        Red_MCInst3_MC1_v3_1[0] ), .Z(MCInst3_MC1_v3_3 [3]) );
  XNOR2_X1 MCInst3_MC1_r0Inst_XORInst_0_0_U3  ( .A(
        MCInst3_MC1_r0Inst_XORInst_0_0_n5 ), .B(
        MCInst3_MC1_r0Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[56]) );
  XNOR2_X1 MCInst3_MC1_r0Inst_XORInst_0_0_U2  ( .A(MCInst3_MC1_v3_2 [2]), 
        .B(MCInst3_MC1_v2_0 [0]), .ZN(MCInst3_MC1_r0Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst3_MC1_r0Inst_XORInst_0_0_U1  ( .A(MCInst3_MC1_v0_3 [3]), .B(
        MCInst3_MC1_v1_0 [0]), .Z(MCInst3_MC1_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst3_MC1_r0Inst_XORInst_0_1_U3  ( .A(
        MCInst3_MC1_r0Inst_XORInst_0_1_n5 ), .B(
        MCInst3_MC1_r0Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[57]) );
  XNOR2_X1 MCInst3_MC1_r0Inst_XORInst_0_1_U2  ( .A(MCInst3_MC1_v3_0 [1]), 
        .B(MCInst3_MC1_v2_0 [1]), .ZN(MCInst3_MC1_r0Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst3_MC1_r0Inst_XORInst_0_1_U1  ( .A(MCInst3_MC1_v0_0 [1]), .B(
        MCInst3_MC1_v1_3 [2]), .Z(MCInst3_MC1_r0Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst3_MC1_r0Inst_XORInst_0_2_U3  ( .A(
        MCInst3_MC1_r0Inst_XORInst_0_2_n5 ), .B(
        MCInst3_MC1_r0Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[58]) );
  XNOR2_X1 MCInst3_MC1_r0Inst_XORInst_0_2_U2  ( .A(MCInst3_MC1_v3_0 [2]), 
        .B(MCInst3_MC1_v2_0 [2]), .ZN(MCInst3_MC1_r0Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst3_MC1_r0Inst_XORInst_0_2_U1  ( .A(MCInst3_MC1_v0_0 [2]), .B(
        Red_MCInst3_MC1_v1_1[0] ), .Z(MCInst3_MC1_r0Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst3_MC1_r0Inst_XORInst_0_3_U3  ( .A(
        MCInst3_MC1_r0Inst_XORInst_0_3_n5 ), .B(
        MCInst3_MC1_r0Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[59]) );
  XNOR2_X1 MCInst3_MC1_r0Inst_XORInst_0_3_U2  ( .A(Red_MCInst3_MC1_v3_1[0] ), 
        .B(MCInst3_MC1_v2_0 [3]), .ZN(MCInst3_MC1_r0Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst3_MC1_r0Inst_XORInst_0_3_U1  ( .A(MCInst3_MC1_v0_0 [3]), .B(
        MCInst3_MC1_v1_0 [3]), .Z(MCInst3_MC1_r0Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst3_MC1_r1Inst_XORInst_0_0_U3  ( .A(
        MCInst3_MC1_r1Inst_XORInst_0_0_n5 ), .B(
        MCInst3_MC1_r1Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[40]) );
  XNOR2_X1 MCInst3_MC1_r1Inst_XORInst_0_0_U2  ( .A(MCInst3_MC1_v3_1 [0]), 
        .B(MCInst3_MC1_v2_1 [0]), .ZN(MCInst3_MC1_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst3_MC1_r1Inst_XORInst_0_0_U1  ( .A(MCInst3_MC1_v0_0 [3]), .B(
        MCInst3_MC1_v1_1 [0]), .Z(MCInst3_MC1_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst3_MC1_r1Inst_XORInst_0_1_U3  ( .A(
        MCInst3_MC1_r1Inst_XORInst_0_1_n5 ), .B(
        MCInst3_MC1_r1Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[41]) );
  XNOR2_X1 MCInst3_MC1_r1Inst_XORInst_0_1_U2  ( .A(MCInst3_MC1_v3_1 [1]), 
        .B(MCInst3_MC1_v2_1 [1]), .ZN(MCInst3_MC1_r1Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst3_MC1_r1Inst_XORInst_0_1_U1  ( .A(MCInst3_MC1_v0_1 [1]), .B(
        MCInst3_MC1_v1_1 [1]), .Z(MCInst3_MC1_r1Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst3_MC1_r1Inst_XORInst_0_2_U3  ( .A(
        MCInst3_MC1_r1Inst_XORInst_0_2_n5 ), .B(
        MCInst3_MC1_r1Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[42]) );
  XNOR2_X1 MCInst3_MC1_r1Inst_XORInst_0_2_U2  ( .A(MCInst3_MC1_v3_1 [2]), 
        .B(MCInst3_MC1_v2_1 [2]), .ZN(MCInst3_MC1_r1Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst3_MC1_r1Inst_XORInst_0_2_U1  ( .A(MCInst3_MC1_v0_1 [2]), .B(
        MCInst3_MC1_v1_1 [2]), .Z(MCInst3_MC1_r1Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst3_MC1_r1Inst_XORInst_0_3_U3  ( .A(
        MCInst3_MC1_r1Inst_XORInst_0_3_n5 ), .B(
        MCInst3_MC1_r1Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[43]) );
  XNOR2_X1 MCInst3_MC1_r1Inst_XORInst_0_3_U2  ( .A(MCInst3_MC1_v3_1 [3]), 
        .B(MCInst3_MC1_v2_1 [3]), .ZN(MCInst3_MC1_r1Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst3_MC1_r1Inst_XORInst_0_3_U1  ( .A(MCInst3_MC1_v0_1 [3]), .B(
        MCInst3_MC1_v1_1 [3]), .Z(MCInst3_MC1_r1Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst3_MC1_r2Inst_XORInst_0_0_U3  ( .A(
        MCInst3_MC1_r2Inst_XORInst_0_0_n5 ), .B(
        MCInst3_MC1_r2Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[24]) );
  XNOR2_X1 MCInst3_MC1_r2Inst_XORInst_0_0_U2  ( .A(MCInst3_MC1_v3_2 [0]), 
        .B(MCInst3_MC1_v2_2 [0]), .ZN(MCInst3_MC1_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst3_MC1_r2Inst_XORInst_0_0_U1  ( .A(MCInst3_MC1_v0_2 [0]), .B(
        MCInst3_MC1_v1_2 [0]), .Z(MCInst3_MC1_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst3_MC1_r2Inst_XORInst_0_1_U3  ( .A(
        MCInst3_MC1_r2Inst_XORInst_0_1_n5 ), .B(
        MCInst3_MC1_r2Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[25]) );
  XNOR2_X1 MCInst3_MC1_r2Inst_XORInst_0_1_U2  ( .A(Red_MCInst3_MC1_v3_1[0] ), 
        .B(MCInst3_MC1_v2_2 [1]), .ZN(MCInst3_MC1_r2Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst3_MC1_r2Inst_XORInst_0_1_U1  ( .A(MCInst3_MC1_v0_2 [1]), .B(
        MCInst3_MC1_v1_2 [1]), .Z(MCInst3_MC1_r2Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst3_MC1_r2Inst_XORInst_0_2_U3  ( .A(
        MCInst3_MC1_r2Inst_XORInst_0_2_n5 ), .B(
        MCInst3_MC1_r2Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[26]) );
  XNOR2_X1 MCInst3_MC1_r2Inst_XORInst_0_2_U2  ( .A(MCInst3_MC1_v3_2 [2]), 
        .B(MCInst3_MC1_v2_2 [2]), .ZN(MCInst3_MC1_r2Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst3_MC1_r2Inst_XORInst_0_2_U1  ( .A(MCInst3_MC1_v0_2 [2]), .B(
        MCInst3_MC1_v1_2 [2]), .Z(MCInst3_MC1_r2Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst3_MC1_r2Inst_XORInst_0_3_U3  ( .A(
        MCInst3_MC1_r2Inst_XORInst_0_3_n5 ), .B(
        MCInst3_MC1_r2Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[27]) );
  XNOR2_X1 MCInst3_MC1_r2Inst_XORInst_0_3_U2  ( .A(MCInst3_MC1_v3_2 [3]), 
        .B(MCInst3_MC1_v2_2 [3]), .ZN(MCInst3_MC1_r2Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst3_MC1_r2Inst_XORInst_0_3_U1  ( .A(MCInst3_MC1_v0_2 [3]), .B(
        MCInst3_MC1_v1_2 [3]), .Z(MCInst3_MC1_r2Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst3_MC1_r3Inst_XORInst_0_0_U3  ( .A(
        MCInst3_MC1_r3Inst_XORInst_0_0_n5 ), .B(
        MCInst3_MC1_r3Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[8]) );
  XNOR2_X1 MCInst3_MC1_r3Inst_XORInst_0_0_U2  ( .A(MCInst3_MC1_v3_3 [0]), 
        .B(MCInst3_MC1_v2_3 [0]), .ZN(MCInst3_MC1_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst3_MC1_r3Inst_XORInst_0_0_U1  ( .A(MCInst3_MC1_v0_3 [0]), .B(
        MCInst3_MC1_v1_0 [3]), .Z(MCInst3_MC1_r3Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst3_MC1_r3Inst_XORInst_0_1_U3  ( .A(
        MCInst3_MC1_r3Inst_XORInst_0_1_n5 ), .B(
        MCInst3_MC1_r3Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[9]) );
  XNOR2_X1 MCInst3_MC1_r3Inst_XORInst_0_1_U2  ( .A(MCInst3_MC1_v3_3 [1]), 
        .B(MCInst3_MC1_v2_3 [1]), .ZN(MCInst3_MC1_r3Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst3_MC1_r3Inst_XORInst_0_1_U1  ( .A(MCInst3_MC1_v0_3 [1]), .B(
        MCInst3_MC1_v1_3 [1]), .Z(MCInst3_MC1_r3Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst3_MC1_r3Inst_XORInst_0_2_U3  ( .A(
        MCInst3_MC1_r3Inst_XORInst_0_2_n5 ), .B(
        MCInst3_MC1_r3Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[10]) );
  XNOR2_X1 MCInst3_MC1_r3Inst_XORInst_0_2_U2  ( .A(MCInst3_MC1_v3_3 [2]), 
        .B(MCInst3_MC1_v2_3 [2]), .ZN(MCInst3_MC1_r3Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst3_MC1_r3Inst_XORInst_0_2_U1  ( .A(MCInst3_MC1_v0_0 [3]), .B(
        MCInst3_MC1_v1_3 [2]), .Z(MCInst3_MC1_r3Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst3_MC1_r3Inst_XORInst_0_3_U3  ( .A(
        MCInst3_MC1_r3Inst_XORInst_0_3_n5 ), .B(
        MCInst3_MC1_r3Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[11]) );
  XNOR2_X1 MCInst3_MC1_r3Inst_XORInst_0_3_U2  ( .A(MCInst3_MC1_v3_3 [3]), 
        .B(MCInst3_MC1_v2_3 [3]), .ZN(MCInst3_MC1_r3Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst3_MC1_r3Inst_XORInst_0_3_U1  ( .A(MCInst3_MC1_v0_3 [3]), .B(
        Red_MCInst3_MC1_v1_1[0] ), .Z(MCInst3_MC1_r3Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst3_MC2_v0_2Inst_0_U4  ( .A(MCInst3_MC2_v0_2Inst_0_n2 ), .B(
        MCInst3_MC2_v0_0 [3]), .ZN(MCInst3_MC2_v0_2 [0]) );
  XNOR2_X1 MCInst3_MC2_v0_2Inst_0_U3  ( .A(MCInst3_MC2_v0_3 [0]), .B(
        Red_MCInst3_MC2_v0_1[0] ), .ZN(MCInst3_MC2_v0_2Inst_0_n2 ) );
  XOR2_X1 MCInst3_MC2_v1_1Inst_0_U3  ( .A(Red_MCInst3_MC2_v1_1[0] ), .B(
        MCInst3_MC2_v1_0 [3]), .Z(MCInst3_MC2_v1_1 [0]) );
  XNOR2_X1 MCInst3_MC2_v1_2Inst_0_U4  ( .A(MCInst3_MC2_v1_2Inst_0_n2 ), .B(
        Red_MCInst3_MC2_v1_1[0] ), .ZN(MCInst3_MC2_v1_2 [0]) );
  XNOR2_X1 MCInst3_MC2_v1_2Inst_0_U3  ( .A(MCInst3_MC2_v1_0 [3]), .B(
        MCInst3_MC2_v1_3 [2]), .ZN(MCInst3_MC2_v1_2Inst_0_n2 ) );
  XOR2_X1 MCInst3_MC2_v2_1Inst_0_U3  ( .A(MCInst3_MC2_v2_3 [1]), .B(
        MCInst3_MC2_v2_0 [3]), .Z(MCInst3_MC2_v2_1 [0]) );
  XOR2_X1 MCInst3_MC2_v2_2Inst_0_U3  ( .A(MCInst3_MC2_v2_0 [2]), .B(
        MCInst3_MC2_v2_0 [0]), .Z(MCInst3_MC2_v2_2 [0]) );
  XNOR2_X1 MCInst3_MC2_v2_3Inst_0_U5  ( .A(MCInst3_MC2_v2_3Inst_0_n4 ), .B(
        MCInst3_MC2_v2_3Inst_0_n3 ), .ZN(MCInst3_MC2_v2_3 [0]) );
  XNOR2_X1 MCInst3_MC2_v2_3Inst_0_U4  ( .A(MCInst3_MC2_v2_0 [2]), .B(
        MCInst3_MC2_v2_3 [1]), .ZN(MCInst3_MC2_v2_3Inst_0_n3 ) );
  XOR2_X1 MCInst3_MC2_v2_3Inst_0_U3  ( .A(MCInst3_MC2_v2_0 [3]), .B(
        MCInst3_MC2_v2_0 [0]), .Z(MCInst3_MC2_v2_3Inst_0_n4 ) );
  XOR2_X1 MCInst3_MC2_v3_1Inst_0_U3  ( .A(Red_MCInst3_MC2_v3_1[0] ), .B(
        MCInst3_MC2_v3_2 [2]), .Z(MCInst3_MC2_v3_1 [0]) );
  XOR2_X1 MCInst3_MC2_v3_2Inst_0_U3  ( .A(MCInst3_MC2_v3_2 [3]), .B(
        MCInst3_MC2_v3_0 [2]), .Z(MCInst3_MC2_v3_2 [0]) );
  XNOR2_X1 MCInst3_MC2_v3_3Inst_0_U4  ( .A(MCInst3_MC2_v3_3Inst_0_n2 ), .B(
        MCInst3_MC2_v3_0 [2]), .ZN(MCInst3_MC2_v3_3 [0]) );
  XNOR2_X1 MCInst3_MC2_v3_3Inst_0_U3  ( .A(MCInst3_MC2_v3_2 [2]), .B(
        MCInst3_MC2_v3_2 [3]), .ZN(MCInst3_MC2_v3_3Inst_0_n2 ) );
  XOR2_X1 MCInst3_MC2_v0_0Inst_1_U3  ( .A(MCInst3_MC2_v0_3 [3]), .B(
        MCInst3_MC2_v0_3 [0]), .Z(MCInst3_MC2_v0_0 [1]) );
  XOR2_X1 MCInst3_MC2_v0_1Inst_1_U3  ( .A(MCInst3_MC2_v0_0 [3]), .B(
        MCInst3_MC2_v0_3 [3]), .Z(MCInst3_MC2_v0_1 [1]) );
  XNOR2_X1 MCInst3_MC2_v0_2Inst_1_U4  ( .A(MCInst3_MC2_v0_2Inst_1_n2 ), .B(
        MCInst3_MC2_v0_3 [3]), .ZN(MCInst3_MC2_v0_2 [1]) );
  XNOR2_X1 MCInst3_MC2_v0_2Inst_1_U3  ( .A(MCInst3_MC2_v0_3 [0]), .B(
        Red_MCInst3_MC2_v0_1[0] ), .ZN(MCInst3_MC2_v0_2Inst_1_n2 ) );
  XOR2_X1 MCInst3_MC2_v0_3Inst_1_U3  ( .A(Red_MCInst3_MC2_v0_1[0] ), .B(
        MCInst3_MC2_v0_3 [0]), .Z(MCInst3_MC2_v0_3 [1]) );
  XOR2_X1 MCInst3_MC2_v1_1Inst_1_U3  ( .A(MCInst3_MC2_v1_0 [0]), .B(
        Red_MCInst3_MC2_v1_1[0] ), .Z(MCInst3_MC2_v1_1 [1]) );
  XOR2_X1 MCInst3_MC2_v1_2Inst_1_U3  ( .A(MCInst3_MC2_v1_0 [0]), .B(
        MCInst3_MC2_v1_3 [2]), .Z(MCInst3_MC2_v1_2 [1]) );
  XOR2_X1 MCInst3_MC2_v1_3Inst_1_U3  ( .A(MCInst3_MC2_v1_0 [0]), .B(
        MCInst3_MC2_v1_0 [3]), .Z(MCInst3_MC2_v1_3 [1]) );
  XOR2_X1 MCInst3_MC2_v2_0Inst_1_U3  ( .A(MCInst3_MC2_v2_3 [1]), .B(
        MCInst3_MC2_v2_0 [0]), .Z(MCInst3_MC2_v2_0 [1]) );
  XNOR2_X1 MCInst3_MC2_v2_1Inst_1_U4  ( .A(MCInst3_MC2_v2_1Inst_1_n2 ), .B(
        MCInst3_MC2_v2_0 [3]), .ZN(MCInst3_MC2_v2_1 [1]) );
  XNOR2_X1 MCInst3_MC2_v2_1Inst_1_U3  ( .A(MCInst3_MC2_v2_0 [0]), .B(
        MCInst3_MC2_v2_0 [2]), .ZN(MCInst3_MC2_v2_1Inst_1_n2 ) );
  XNOR2_X1 MCInst3_MC2_v2_2Inst_1_U5  ( .A(MCInst3_MC2_v2_2Inst_1_n4 ), .B(
        MCInst3_MC2_v2_2Inst_1_n3 ), .ZN(MCInst3_MC2_v2_2 [1]) );
  XNOR2_X1 MCInst3_MC2_v2_2Inst_1_U4  ( .A(MCInst3_MC2_v2_0 [2]), .B(
        MCInst3_MC2_v2_3 [1]), .ZN(MCInst3_MC2_v2_2Inst_1_n3 ) );
  XOR2_X1 MCInst3_MC2_v2_2Inst_1_U3  ( .A(MCInst3_MC2_v2_0 [3]), .B(
        MCInst3_MC2_v2_0 [0]), .Z(MCInst3_MC2_v2_2Inst_1_n4 ) );
  XOR2_X1 MCInst3_MC2_v3_0Inst_1_U3  ( .A(MCInst3_MC2_v3_2 [3]), .B(
        MCInst3_MC2_v3_2 [2]), .Z(MCInst3_MC2_v3_0 [1]) );
  XOR2_X1 MCInst3_MC2_v3_1Inst_1_U3  ( .A(MCInst3_MC2_v3_2 [3]), .B(
        Red_MCInst3_MC2_v3_1[0] ), .Z(MCInst3_MC2_v3_1 [1]) );
  XNOR2_X1 MCInst3_MC2_v3_3Inst_1_U4  ( .A(MCInst3_MC2_v3_3Inst_1_n2 ), .B(
        Red_MCInst3_MC2_v3_1[0] ), .ZN(MCInst3_MC2_v3_3 [1]) );
  XNOR2_X1 MCInst3_MC2_v3_3Inst_1_U3  ( .A(MCInst3_MC2_v3_2 [2]), .B(
        MCInst3_MC2_v3_2 [3]), .ZN(MCInst3_MC2_v3_3Inst_1_n2 ) );
  XOR2_X1 MCInst3_MC2_v0_0Inst_2_U3  ( .A(Red_MCInst3_MC2_v0_1[0] ), .B(
        MCInst3_MC2_v0_3 [0]), .Z(MCInst3_MC2_v0_0 [2]) );
  XOR2_X1 MCInst3_MC2_v0_1Inst_2_U3  ( .A(MCInst3_MC2_v0_3 [3]), .B(
        MCInst3_MC2_v0_3 [0]), .Z(MCInst3_MC2_v0_1 [2]) );
  XOR2_X1 MCInst3_MC2_v0_2Inst_2_U3  ( .A(MCInst3_MC2_v0_0 [3]), .B(
        MCInst3_MC2_v0_3 [0]), .Z(MCInst3_MC2_v0_2 [2]) );
  XNOR2_X1 MCInst3_MC2_v1_1Inst_2_U4  ( .A(MCInst3_MC2_v1_1Inst_2_n2 ), .B(
        MCInst3_MC2_v1_3 [2]), .ZN(MCInst3_MC2_v1_1 [2]) );
  XNOR2_X1 MCInst3_MC2_v1_1Inst_2_U3  ( .A(MCInst3_MC2_v1_0 [3]), .B(
        MCInst3_MC2_v1_0 [0]), .ZN(MCInst3_MC2_v1_1Inst_2_n2 ) );
  XNOR2_X1 MCInst3_MC2_v1_2Inst_2_U4  ( .A(MCInst3_MC2_v1_2Inst_2_n2 ), .B(
        MCInst3_MC2_v1_3 [2]), .ZN(MCInst3_MC2_v1_2 [2]) );
  XNOR2_X1 MCInst3_MC2_v1_2Inst_2_U3  ( .A(Red_MCInst3_MC2_v1_1[0] ), .B(
        MCInst3_MC2_v1_0 [0]), .ZN(MCInst3_MC2_v1_2Inst_2_n2 ) );
  XNOR2_X1 MCInst3_MC2_v2_1Inst_2_U4  ( .A(MCInst3_MC2_v2_1Inst_2_n2 ), .B(
        MCInst3_MC2_v2_0 [3]), .ZN(MCInst3_MC2_v2_1 [2]) );
  XNOR2_X1 MCInst3_MC2_v2_1Inst_2_U3  ( .A(MCInst3_MC2_v2_0 [0]), .B(
        MCInst3_MC2_v2_3 [1]), .ZN(MCInst3_MC2_v2_1Inst_2_n2 ) );
  XNOR2_X1 MCInst3_MC2_v2_2Inst_2_U4  ( .A(MCInst3_MC2_v2_2Inst_2_n2 ), .B(
        MCInst3_MC2_v2_0 [3]), .ZN(MCInst3_MC2_v2_2 [2]) );
  XNOR2_X1 MCInst3_MC2_v2_2Inst_2_U3  ( .A(MCInst3_MC2_v2_0 [0]), .B(
        MCInst3_MC2_v2_0 [2]), .ZN(MCInst3_MC2_v2_2Inst_2_n2 ) );
  XOR2_X1 MCInst3_MC2_v2_3Inst_2_U3  ( .A(MCInst3_MC2_v2_3 [1]), .B(
        MCInst3_MC2_v2_0 [2]), .Z(MCInst3_MC2_v2_3 [2]) );
  XNOR2_X1 MCInst3_MC2_v3_1Inst_2_U4  ( .A(MCInst3_MC2_v3_1Inst_2_n2 ), .B(
        MCInst3_MC2_v3_0 [2]), .ZN(MCInst3_MC2_v3_1 [2]) );
  XNOR2_X1 MCInst3_MC2_v3_1Inst_2_U3  ( .A(MCInst3_MC2_v3_2 [2]), .B(
        MCInst3_MC2_v3_2 [3]), .ZN(MCInst3_MC2_v3_1Inst_2_n2 ) );
  XOR2_X1 MCInst3_MC2_v3_3Inst_2_U3  ( .A(MCInst3_MC2_v3_0 [2]), .B(
        MCInst3_MC2_v3_2 [2]), .Z(MCInst3_MC2_v3_3 [2]) );
  XOR2_X1 MCInst3_MC2_v0_1Inst_3_U3  ( .A(Red_MCInst3_MC2_v0_1[0] ), .B(
        MCInst3_MC2_v0_3 [0]), .Z(MCInst3_MC2_v0_1 [3]) );
  XOR2_X1 MCInst3_MC2_v0_2Inst_3_U3  ( .A(Red_MCInst3_MC2_v0_1[0] ), .B(
        MCInst3_MC2_v0_3 [3]), .Z(MCInst3_MC2_v0_2 [3]) );
  XOR2_X1 MCInst3_MC2_v1_1Inst_3_U3  ( .A(MCInst3_MC2_v1_3 [2]), .B(
        Red_MCInst3_MC2_v1_1[0] ), .Z(MCInst3_MC2_v1_1 [3]) );
  XNOR2_X1 MCInst3_MC2_v1_2Inst_3_U5  ( .A(MCInst3_MC2_v1_2Inst_3_n4 ), .B(
        MCInst3_MC2_v1_2Inst_3_n3 ), .ZN(MCInst3_MC2_v1_2 [3]) );
  XNOR2_X1 MCInst3_MC2_v1_2Inst_3_U4  ( .A(MCInst3_MC2_v1_3 [2]), .B(
        MCInst3_MC2_v1_0 [0]), .ZN(MCInst3_MC2_v1_2Inst_3_n3 ) );
  XOR2_X1 MCInst3_MC2_v1_2Inst_3_U3  ( .A(Red_MCInst3_MC2_v1_1[0] ), .B(
        MCInst3_MC2_v1_0 [3]), .Z(MCInst3_MC2_v1_2Inst_3_n4 ) );
  XOR2_X1 MCInst3_MC2_v2_1Inst_3_U3  ( .A(MCInst3_MC2_v2_0 [2]), .B(
        MCInst3_MC2_v2_0 [0]), .Z(MCInst3_MC2_v2_1 [3]) );
  XNOR2_X1 MCInst3_MC2_v2_2Inst_3_U4  ( .A(MCInst3_MC2_v2_2Inst_3_n2 ), .B(
        MCInst3_MC2_v2_0 [3]), .ZN(MCInst3_MC2_v2_2 [3]) );
  XNOR2_X1 MCInst3_MC2_v2_2Inst_3_U3  ( .A(MCInst3_MC2_v2_0 [0]), .B(
        MCInst3_MC2_v2_3 [1]), .ZN(MCInst3_MC2_v2_2Inst_3_n2 ) );
  XNOR2_X1 MCInst3_MC2_v2_3Inst_3_U4  ( .A(MCInst3_MC2_v2_3Inst_3_n2 ), .B(
        MCInst3_MC2_v2_0 [2]), .ZN(MCInst3_MC2_v2_3 [3]) );
  XNOR2_X1 MCInst3_MC2_v2_3Inst_3_U3  ( .A(MCInst3_MC2_v2_0 [3]), .B(
        MCInst3_MC2_v2_3 [1]), .ZN(MCInst3_MC2_v2_3Inst_3_n2 ) );
  XOR2_X1 MCInst3_MC2_v3_1Inst_3_U3  ( .A(MCInst3_MC2_v3_0 [2]), .B(
        Red_MCInst3_MC2_v3_1[0] ), .Z(MCInst3_MC2_v3_1 [3]) );
  XOR2_X1 MCInst3_MC2_v3_3Inst_3_U3  ( .A(MCInst3_MC2_v3_2 [3]), .B(
        Red_MCInst3_MC2_v3_1[0] ), .Z(MCInst3_MC2_v3_3 [3]) );
  XNOR2_X1 MCInst3_MC2_r0Inst_XORInst_0_0_U3  ( .A(
        MCInst3_MC2_r0Inst_XORInst_0_0_n5 ), .B(
        MCInst3_MC2_r0Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[52]) );
  XNOR2_X1 MCInst3_MC2_r0Inst_XORInst_0_0_U2  ( .A(MCInst3_MC2_v3_2 [2]), 
        .B(MCInst3_MC2_v2_0 [0]), .ZN(MCInst3_MC2_r0Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst3_MC2_r0Inst_XORInst_0_0_U1  ( .A(MCInst3_MC2_v0_3 [3]), .B(
        MCInst3_MC2_v1_0 [0]), .Z(MCInst3_MC2_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst3_MC2_r0Inst_XORInst_0_1_U3  ( .A(
        MCInst3_MC2_r0Inst_XORInst_0_1_n5 ), .B(
        MCInst3_MC2_r0Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[53]) );
  XNOR2_X1 MCInst3_MC2_r0Inst_XORInst_0_1_U2  ( .A(MCInst3_MC2_v3_0 [1]), 
        .B(MCInst3_MC2_v2_0 [1]), .ZN(MCInst3_MC2_r0Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst3_MC2_r0Inst_XORInst_0_1_U1  ( .A(MCInst3_MC2_v0_0 [1]), .B(
        MCInst3_MC2_v1_3 [2]), .Z(MCInst3_MC2_r0Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst3_MC2_r0Inst_XORInst_0_2_U3  ( .A(
        MCInst3_MC2_r0Inst_XORInst_0_2_n5 ), .B(
        MCInst3_MC2_r0Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[54]) );
  XNOR2_X1 MCInst3_MC2_r0Inst_XORInst_0_2_U2  ( .A(MCInst3_MC2_v3_0 [2]), 
        .B(MCInst3_MC2_v2_0 [2]), .ZN(MCInst3_MC2_r0Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst3_MC2_r0Inst_XORInst_0_2_U1  ( .A(MCInst3_MC2_v0_0 [2]), .B(
        Red_MCInst3_MC2_v1_1[0] ), .Z(MCInst3_MC2_r0Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst3_MC2_r0Inst_XORInst_0_3_U3  ( .A(
        MCInst3_MC2_r0Inst_XORInst_0_3_n5 ), .B(
        MCInst3_MC2_r0Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[55]) );
  XNOR2_X1 MCInst3_MC2_r0Inst_XORInst_0_3_U2  ( .A(Red_MCInst3_MC2_v3_1[0] ), 
        .B(MCInst3_MC2_v2_0 [3]), .ZN(MCInst3_MC2_r0Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst3_MC2_r0Inst_XORInst_0_3_U1  ( .A(MCInst3_MC2_v0_0 [3]), .B(
        MCInst3_MC2_v1_0 [3]), .Z(MCInst3_MC2_r0Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst3_MC2_r1Inst_XORInst_0_0_U3  ( .A(
        MCInst3_MC2_r1Inst_XORInst_0_0_n5 ), .B(
        MCInst3_MC2_r1Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[36]) );
  XNOR2_X1 MCInst3_MC2_r1Inst_XORInst_0_0_U2  ( .A(MCInst3_MC2_v3_1 [0]), 
        .B(MCInst3_MC2_v2_1 [0]), .ZN(MCInst3_MC2_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst3_MC2_r1Inst_XORInst_0_0_U1  ( .A(MCInst3_MC2_v0_0 [3]), .B(
        MCInst3_MC2_v1_1 [0]), .Z(MCInst3_MC2_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst3_MC2_r1Inst_XORInst_0_1_U3  ( .A(
        MCInst3_MC2_r1Inst_XORInst_0_1_n5 ), .B(
        MCInst3_MC2_r1Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[37]) );
  XNOR2_X1 MCInst3_MC2_r1Inst_XORInst_0_1_U2  ( .A(MCInst3_MC2_v3_1 [1]), 
        .B(MCInst3_MC2_v2_1 [1]), .ZN(MCInst3_MC2_r1Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst3_MC2_r1Inst_XORInst_0_1_U1  ( .A(MCInst3_MC2_v0_1 [1]), .B(
        MCInst3_MC2_v1_1 [1]), .Z(MCInst3_MC2_r1Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst3_MC2_r1Inst_XORInst_0_2_U3  ( .A(
        MCInst3_MC2_r1Inst_XORInst_0_2_n5 ), .B(
        MCInst3_MC2_r1Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[38]) );
  XNOR2_X1 MCInst3_MC2_r1Inst_XORInst_0_2_U2  ( .A(MCInst3_MC2_v3_1 [2]), 
        .B(MCInst3_MC2_v2_1 [2]), .ZN(MCInst3_MC2_r1Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst3_MC2_r1Inst_XORInst_0_2_U1  ( .A(MCInst3_MC2_v0_1 [2]), .B(
        MCInst3_MC2_v1_1 [2]), .Z(MCInst3_MC2_r1Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst3_MC2_r1Inst_XORInst_0_3_U3  ( .A(
        MCInst3_MC2_r1Inst_XORInst_0_3_n5 ), .B(
        MCInst3_MC2_r1Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[39]) );
  XNOR2_X1 MCInst3_MC2_r1Inst_XORInst_0_3_U2  ( .A(MCInst3_MC2_v3_1 [3]), 
        .B(MCInst3_MC2_v2_1 [3]), .ZN(MCInst3_MC2_r1Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst3_MC2_r1Inst_XORInst_0_3_U1  ( .A(MCInst3_MC2_v0_1 [3]), .B(
        MCInst3_MC2_v1_1 [3]), .Z(MCInst3_MC2_r1Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst3_MC2_r2Inst_XORInst_0_0_U3  ( .A(
        MCInst3_MC2_r2Inst_XORInst_0_0_n5 ), .B(
        MCInst3_MC2_r2Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[20]) );
  XNOR2_X1 MCInst3_MC2_r2Inst_XORInst_0_0_U2  ( .A(MCInst3_MC2_v3_2 [0]), 
        .B(MCInst3_MC2_v2_2 [0]), .ZN(MCInst3_MC2_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst3_MC2_r2Inst_XORInst_0_0_U1  ( .A(MCInst3_MC2_v0_2 [0]), .B(
        MCInst3_MC2_v1_2 [0]), .Z(MCInst3_MC2_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst3_MC2_r2Inst_XORInst_0_1_U3  ( .A(
        MCInst3_MC2_r2Inst_XORInst_0_1_n5 ), .B(
        MCInst3_MC2_r2Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[21]) );
  XNOR2_X1 MCInst3_MC2_r2Inst_XORInst_0_1_U2  ( .A(Red_MCInst3_MC2_v3_1[0] ), 
        .B(MCInst3_MC2_v2_2 [1]), .ZN(MCInst3_MC2_r2Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst3_MC2_r2Inst_XORInst_0_1_U1  ( .A(MCInst3_MC2_v0_2 [1]), .B(
        MCInst3_MC2_v1_2 [1]), .Z(MCInst3_MC2_r2Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst3_MC2_r2Inst_XORInst_0_2_U3  ( .A(
        MCInst3_MC2_r2Inst_XORInst_0_2_n5 ), .B(
        MCInst3_MC2_r2Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[22]) );
  XNOR2_X1 MCInst3_MC2_r2Inst_XORInst_0_2_U2  ( .A(MCInst3_MC2_v3_2 [2]), 
        .B(MCInst3_MC2_v2_2 [2]), .ZN(MCInst3_MC2_r2Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst3_MC2_r2Inst_XORInst_0_2_U1  ( .A(MCInst3_MC2_v0_2 [2]), .B(
        MCInst3_MC2_v1_2 [2]), .Z(MCInst3_MC2_r2Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst3_MC2_r2Inst_XORInst_0_3_U3  ( .A(
        MCInst3_MC2_r2Inst_XORInst_0_3_n5 ), .B(
        MCInst3_MC2_r2Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[23]) );
  XNOR2_X1 MCInst3_MC2_r2Inst_XORInst_0_3_U2  ( .A(MCInst3_MC2_v3_2 [3]), 
        .B(MCInst3_MC2_v2_2 [3]), .ZN(MCInst3_MC2_r2Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst3_MC2_r2Inst_XORInst_0_3_U1  ( .A(MCInst3_MC2_v0_2 [3]), .B(
        MCInst3_MC2_v1_2 [3]), .Z(MCInst3_MC2_r2Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst3_MC2_r3Inst_XORInst_0_0_U3  ( .A(
        MCInst3_MC2_r3Inst_XORInst_0_0_n5 ), .B(
        MCInst3_MC2_r3Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[4]) );
  XNOR2_X1 MCInst3_MC2_r3Inst_XORInst_0_0_U2  ( .A(MCInst3_MC2_v3_3 [0]), 
        .B(MCInst3_MC2_v2_3 [0]), .ZN(MCInst3_MC2_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst3_MC2_r3Inst_XORInst_0_0_U1  ( .A(MCInst3_MC2_v0_3 [0]), .B(
        MCInst3_MC2_v1_0 [3]), .Z(MCInst3_MC2_r3Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst3_MC2_r3Inst_XORInst_0_1_U3  ( .A(
        MCInst3_MC2_r3Inst_XORInst_0_1_n5 ), .B(
        MCInst3_MC2_r3Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[5]) );
  XNOR2_X1 MCInst3_MC2_r3Inst_XORInst_0_1_U2  ( .A(MCInst3_MC2_v3_3 [1]), 
        .B(MCInst3_MC2_v2_3 [1]), .ZN(MCInst3_MC2_r3Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst3_MC2_r3Inst_XORInst_0_1_U1  ( .A(MCInst3_MC2_v0_3 [1]), .B(
        MCInst3_MC2_v1_3 [1]), .Z(MCInst3_MC2_r3Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst3_MC2_r3Inst_XORInst_0_2_U3  ( .A(
        MCInst3_MC2_r3Inst_XORInst_0_2_n5 ), .B(
        MCInst3_MC2_r3Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[6]) );
  XNOR2_X1 MCInst3_MC2_r3Inst_XORInst_0_2_U2  ( .A(MCInst3_MC2_v3_3 [2]), 
        .B(MCInst3_MC2_v2_3 [2]), .ZN(MCInst3_MC2_r3Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst3_MC2_r3Inst_XORInst_0_2_U1  ( .A(MCInst3_MC2_v0_0 [3]), .B(
        MCInst3_MC2_v1_3 [2]), .Z(MCInst3_MC2_r3Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst3_MC2_r3Inst_XORInst_0_3_U3  ( .A(
        MCInst3_MC2_r3Inst_XORInst_0_3_n5 ), .B(
        MCInst3_MC2_r3Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[7]) );
  XNOR2_X1 MCInst3_MC2_r3Inst_XORInst_0_3_U2  ( .A(MCInst3_MC2_v3_3 [3]), 
        .B(MCInst3_MC2_v2_3 [3]), .ZN(MCInst3_MC2_r3Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst3_MC2_r3Inst_XORInst_0_3_U1  ( .A(MCInst3_MC2_v0_3 [3]), .B(
        Red_MCInst3_MC2_v1_1[0] ), .Z(MCInst3_MC2_r3Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst3_MC3_v0_2Inst_0_U4  ( .A(MCInst3_MC3_v0_2Inst_0_n2 ), .B(
        MCInst3_MC3_v0_0 [3]), .ZN(MCInst3_MC3_v0_2 [0]) );
  XNOR2_X1 MCInst3_MC3_v0_2Inst_0_U3  ( .A(MCInst3_MC3_v0_3 [0]), .B(
        Red_MCInst3_MC3_v0_1[0] ), .ZN(MCInst3_MC3_v0_2Inst_0_n2 ) );
  XOR2_X1 MCInst3_MC3_v1_1Inst_0_U3  ( .A(Red_MCInst3_MC3_v1_1[0] ), .B(
        MCInst3_MC3_v1_0 [3]), .Z(MCInst3_MC3_v1_1 [0]) );
  XNOR2_X1 MCInst3_MC3_v1_2Inst_0_U4  ( .A(MCInst3_MC3_v1_2Inst_0_n2 ), .B(
        Red_MCInst3_MC3_v1_1[0] ), .ZN(MCInst3_MC3_v1_2 [0]) );
  XNOR2_X1 MCInst3_MC3_v1_2Inst_0_U3  ( .A(MCInst3_MC3_v1_0 [3]), .B(
        MCInst3_MC3_v1_3 [2]), .ZN(MCInst3_MC3_v1_2Inst_0_n2 ) );
  XOR2_X1 MCInst3_MC3_v2_1Inst_0_U3  ( .A(MCInst3_MC3_v2_3 [1]), .B(
        MCInst3_MC3_v2_0 [3]), .Z(MCInst3_MC3_v2_1 [0]) );
  XOR2_X1 MCInst3_MC3_v2_2Inst_0_U3  ( .A(MCInst3_MC3_v2_0 [2]), .B(
        MCInst3_MC3_v2_0 [0]), .Z(MCInst3_MC3_v2_2 [0]) );
  XNOR2_X1 MCInst3_MC3_v2_3Inst_0_U5  ( .A(MCInst3_MC3_v2_3Inst_0_n4 ), .B(
        MCInst3_MC3_v2_3Inst_0_n3 ), .ZN(MCInst3_MC3_v2_3 [0]) );
  XNOR2_X1 MCInst3_MC3_v2_3Inst_0_U4  ( .A(MCInst3_MC3_v2_0 [2]), .B(
        MCInst3_MC3_v2_3 [1]), .ZN(MCInst3_MC3_v2_3Inst_0_n3 ) );
  XOR2_X1 MCInst3_MC3_v2_3Inst_0_U3  ( .A(MCInst3_MC3_v2_0 [3]), .B(
        MCInst3_MC3_v2_0 [0]), .Z(MCInst3_MC3_v2_3Inst_0_n4 ) );
  XOR2_X1 MCInst3_MC3_v3_1Inst_0_U3  ( .A(Red_MCInst3_MC3_v3_1[0] ), .B(
        MCInst3_MC3_v3_2 [2]), .Z(MCInst3_MC3_v3_1 [0]) );
  XOR2_X1 MCInst3_MC3_v3_2Inst_0_U3  ( .A(MCInst3_MC3_v3_2 [3]), .B(
        MCInst3_MC3_v3_0 [2]), .Z(MCInst3_MC3_v3_2 [0]) );
  XNOR2_X1 MCInst3_MC3_v3_3Inst_0_U4  ( .A(MCInst3_MC3_v3_3Inst_0_n2 ), .B(
        MCInst3_MC3_v3_0 [2]), .ZN(MCInst3_MC3_v3_3 [0]) );
  XNOR2_X1 MCInst3_MC3_v3_3Inst_0_U3  ( .A(MCInst3_MC3_v3_2 [2]), .B(
        MCInst3_MC3_v3_2 [3]), .ZN(MCInst3_MC3_v3_3Inst_0_n2 ) );
  XOR2_X1 MCInst3_MC3_v0_0Inst_1_U3  ( .A(MCInst3_MC3_v0_3 [3]), .B(
        MCInst3_MC3_v0_3 [0]), .Z(MCInst3_MC3_v0_0 [1]) );
  XOR2_X1 MCInst3_MC3_v0_1Inst_1_U3  ( .A(MCInst3_MC3_v0_0 [3]), .B(
        MCInst3_MC3_v0_3 [3]), .Z(MCInst3_MC3_v0_1 [1]) );
  XNOR2_X1 MCInst3_MC3_v0_2Inst_1_U4  ( .A(MCInst3_MC3_v0_2Inst_1_n2 ), .B(
        MCInst3_MC3_v0_3 [3]), .ZN(MCInst3_MC3_v0_2 [1]) );
  XNOR2_X1 MCInst3_MC3_v0_2Inst_1_U3  ( .A(MCInst3_MC3_v0_3 [0]), .B(
        Red_MCInst3_MC3_v0_1[0] ), .ZN(MCInst3_MC3_v0_2Inst_1_n2 ) );
  XOR2_X1 MCInst3_MC3_v0_3Inst_1_U3  ( .A(Red_MCInst3_MC3_v0_1[0] ), .B(
        MCInst3_MC3_v0_3 [0]), .Z(MCInst3_MC3_v0_3 [1]) );
  XOR2_X1 MCInst3_MC3_v1_1Inst_1_U3  ( .A(MCInst3_MC3_v1_0 [0]), .B(
        Red_MCInst3_MC3_v1_1[0] ), .Z(MCInst3_MC3_v1_1 [1]) );
  XOR2_X1 MCInst3_MC3_v1_2Inst_1_U3  ( .A(MCInst3_MC3_v1_0 [0]), .B(
        MCInst3_MC3_v1_3 [2]), .Z(MCInst3_MC3_v1_2 [1]) );
  XOR2_X1 MCInst3_MC3_v1_3Inst_1_U3  ( .A(MCInst3_MC3_v1_0 [0]), .B(
        MCInst3_MC3_v1_0 [3]), .Z(MCInst3_MC3_v1_3 [1]) );
  XOR2_X1 MCInst3_MC3_v2_0Inst_1_U3  ( .A(MCInst3_MC3_v2_3 [1]), .B(
        MCInst3_MC3_v2_0 [0]), .Z(MCInst3_MC3_v2_0 [1]) );
  XNOR2_X1 MCInst3_MC3_v2_1Inst_1_U4  ( .A(MCInst3_MC3_v2_1Inst_1_n2 ), .B(
        MCInst3_MC3_v2_0 [3]), .ZN(MCInst3_MC3_v2_1 [1]) );
  XNOR2_X1 MCInst3_MC3_v2_1Inst_1_U3  ( .A(MCInst3_MC3_v2_0 [0]), .B(
        MCInst3_MC3_v2_0 [2]), .ZN(MCInst3_MC3_v2_1Inst_1_n2 ) );
  XNOR2_X1 MCInst3_MC3_v2_2Inst_1_U5  ( .A(MCInst3_MC3_v2_2Inst_1_n4 ), .B(
        MCInst3_MC3_v2_2Inst_1_n3 ), .ZN(MCInst3_MC3_v2_2 [1]) );
  XNOR2_X1 MCInst3_MC3_v2_2Inst_1_U4  ( .A(MCInst3_MC3_v2_0 [2]), .B(
        MCInst3_MC3_v2_3 [1]), .ZN(MCInst3_MC3_v2_2Inst_1_n3 ) );
  XOR2_X1 MCInst3_MC3_v2_2Inst_1_U3  ( .A(MCInst3_MC3_v2_0 [3]), .B(
        MCInst3_MC3_v2_0 [0]), .Z(MCInst3_MC3_v2_2Inst_1_n4 ) );
  XOR2_X1 MCInst3_MC3_v3_0Inst_1_U3  ( .A(MCInst3_MC3_v3_2 [3]), .B(
        MCInst3_MC3_v3_2 [2]), .Z(MCInst3_MC3_v3_0 [1]) );
  XOR2_X1 MCInst3_MC3_v3_1Inst_1_U3  ( .A(MCInst3_MC3_v3_2 [3]), .B(
        Red_MCInst3_MC3_v3_1[0] ), .Z(MCInst3_MC3_v3_1 [1]) );
  XNOR2_X1 MCInst3_MC3_v3_3Inst_1_U4  ( .A(MCInst3_MC3_v3_3Inst_1_n2 ), .B(
        Red_MCInst3_MC3_v3_1[0] ), .ZN(MCInst3_MC3_v3_3 [1]) );
  XNOR2_X1 MCInst3_MC3_v3_3Inst_1_U3  ( .A(MCInst3_MC3_v3_2 [2]), .B(
        MCInst3_MC3_v3_2 [3]), .ZN(MCInst3_MC3_v3_3Inst_1_n2 ) );
  XOR2_X1 MCInst3_MC3_v0_0Inst_2_U3  ( .A(Red_MCInst3_MC3_v0_1[0] ), .B(
        MCInst3_MC3_v0_3 [0]), .Z(MCInst3_MC3_v0_0 [2]) );
  XOR2_X1 MCInst3_MC3_v0_1Inst_2_U3  ( .A(MCInst3_MC3_v0_3 [3]), .B(
        MCInst3_MC3_v0_3 [0]), .Z(MCInst3_MC3_v0_1 [2]) );
  XOR2_X1 MCInst3_MC3_v0_2Inst_2_U3  ( .A(MCInst3_MC3_v0_0 [3]), .B(
        MCInst3_MC3_v0_3 [0]), .Z(MCInst3_MC3_v0_2 [2]) );
  XNOR2_X1 MCInst3_MC3_v1_1Inst_2_U4  ( .A(MCInst3_MC3_v1_1Inst_2_n2 ), .B(
        MCInst3_MC3_v1_3 [2]), .ZN(MCInst3_MC3_v1_1 [2]) );
  XNOR2_X1 MCInst3_MC3_v1_1Inst_2_U3  ( .A(MCInst3_MC3_v1_0 [3]), .B(
        MCInst3_MC3_v1_0 [0]), .ZN(MCInst3_MC3_v1_1Inst_2_n2 ) );
  XNOR2_X1 MCInst3_MC3_v1_2Inst_2_U4  ( .A(MCInst3_MC3_v1_2Inst_2_n2 ), .B(
        MCInst3_MC3_v1_3 [2]), .ZN(MCInst3_MC3_v1_2 [2]) );
  XNOR2_X1 MCInst3_MC3_v1_2Inst_2_U3  ( .A(Red_MCInst3_MC3_v1_1[0] ), .B(
        MCInst3_MC3_v1_0 [0]), .ZN(MCInst3_MC3_v1_2Inst_2_n2 ) );
  XNOR2_X1 MCInst3_MC3_v2_1Inst_2_U4  ( .A(MCInst3_MC3_v2_1Inst_2_n2 ), .B(
        MCInst3_MC3_v2_0 [3]), .ZN(MCInst3_MC3_v2_1 [2]) );
  XNOR2_X1 MCInst3_MC3_v2_1Inst_2_U3  ( .A(MCInst3_MC3_v2_0 [0]), .B(
        MCInst3_MC3_v2_3 [1]), .ZN(MCInst3_MC3_v2_1Inst_2_n2 ) );
  XNOR2_X1 MCInst3_MC3_v2_2Inst_2_U4  ( .A(MCInst3_MC3_v2_2Inst_2_n2 ), .B(
        MCInst3_MC3_v2_0 [3]), .ZN(MCInst3_MC3_v2_2 [2]) );
  XNOR2_X1 MCInst3_MC3_v2_2Inst_2_U3  ( .A(MCInst3_MC3_v2_0 [0]), .B(
        MCInst3_MC3_v2_0 [2]), .ZN(MCInst3_MC3_v2_2Inst_2_n2 ) );
  XOR2_X1 MCInst3_MC3_v2_3Inst_2_U3  ( .A(MCInst3_MC3_v2_3 [1]), .B(
        MCInst3_MC3_v2_0 [2]), .Z(MCInst3_MC3_v2_3 [2]) );
  XNOR2_X1 MCInst3_MC3_v3_1Inst_2_U4  ( .A(MCInst3_MC3_v3_1Inst_2_n2 ), .B(
        MCInst3_MC3_v3_0 [2]), .ZN(MCInst3_MC3_v3_1 [2]) );
  XNOR2_X1 MCInst3_MC3_v3_1Inst_2_U3  ( .A(MCInst3_MC3_v3_2 [2]), .B(
        MCInst3_MC3_v3_2 [3]), .ZN(MCInst3_MC3_v3_1Inst_2_n2 ) );
  XOR2_X1 MCInst3_MC3_v3_3Inst_2_U3  ( .A(MCInst3_MC3_v3_0 [2]), .B(
        MCInst3_MC3_v3_2 [2]), .Z(MCInst3_MC3_v3_3 [2]) );
  XOR2_X1 MCInst3_MC3_v0_1Inst_3_U3  ( .A(Red_MCInst3_MC3_v0_1[0] ), .B(
        MCInst3_MC3_v0_3 [0]), .Z(MCInst3_MC3_v0_1 [3]) );
  XOR2_X1 MCInst3_MC3_v0_2Inst_3_U3  ( .A(Red_MCInst3_MC3_v0_1[0] ), .B(
        MCInst3_MC3_v0_3 [3]), .Z(MCInst3_MC3_v0_2 [3]) );
  XOR2_X1 MCInst3_MC3_v1_1Inst_3_U3  ( .A(MCInst3_MC3_v1_3 [2]), .B(
        Red_MCInst3_MC3_v1_1[0] ), .Z(MCInst3_MC3_v1_1 [3]) );
  XNOR2_X1 MCInst3_MC3_v1_2Inst_3_U5  ( .A(MCInst3_MC3_v1_2Inst_3_n4 ), .B(
        MCInst3_MC3_v1_2Inst_3_n3 ), .ZN(MCInst3_MC3_v1_2 [3]) );
  XNOR2_X1 MCInst3_MC3_v1_2Inst_3_U4  ( .A(MCInst3_MC3_v1_3 [2]), .B(
        MCInst3_MC3_v1_0 [0]), .ZN(MCInst3_MC3_v1_2Inst_3_n3 ) );
  XOR2_X1 MCInst3_MC3_v1_2Inst_3_U3  ( .A(Red_MCInst3_MC3_v1_1[0] ), .B(
        MCInst3_MC3_v1_0 [3]), .Z(MCInst3_MC3_v1_2Inst_3_n4 ) );
  XOR2_X1 MCInst3_MC3_v2_1Inst_3_U3  ( .A(MCInst3_MC3_v2_0 [2]), .B(
        MCInst3_MC3_v2_0 [0]), .Z(MCInst3_MC3_v2_1 [3]) );
  XNOR2_X1 MCInst3_MC3_v2_2Inst_3_U4  ( .A(MCInst3_MC3_v2_2Inst_3_n2 ), .B(
        MCInst3_MC3_v2_0 [3]), .ZN(MCInst3_MC3_v2_2 [3]) );
  XNOR2_X1 MCInst3_MC3_v2_2Inst_3_U3  ( .A(MCInst3_MC3_v2_0 [0]), .B(
        MCInst3_MC3_v2_3 [1]), .ZN(MCInst3_MC3_v2_2Inst_3_n2 ) );
  XNOR2_X1 MCInst3_MC3_v2_3Inst_3_U4  ( .A(MCInst3_MC3_v2_3Inst_3_n2 ), .B(
        MCInst3_MC3_v2_0 [2]), .ZN(MCInst3_MC3_v2_3 [3]) );
  XNOR2_X1 MCInst3_MC3_v2_3Inst_3_U3  ( .A(MCInst3_MC3_v2_0 [3]), .B(
        MCInst3_MC3_v2_3 [1]), .ZN(MCInst3_MC3_v2_3Inst_3_n2 ) );
  XOR2_X1 MCInst3_MC3_v3_1Inst_3_U3  ( .A(MCInst3_MC3_v3_0 [2]), .B(
        Red_MCInst3_MC3_v3_1[0] ), .Z(MCInst3_MC3_v3_1 [3]) );
  XOR2_X1 MCInst3_MC3_v3_3Inst_3_U3  ( .A(MCInst3_MC3_v3_2 [3]), .B(
        Red_MCInst3_MC3_v3_1[0] ), .Z(MCInst3_MC3_v3_3 [3]) );
  XNOR2_X1 MCInst3_MC3_r0Inst_XORInst_0_0_U3  ( .A(
        MCInst3_MC3_r0Inst_XORInst_0_0_n5 ), .B(
        MCInst3_MC3_r0Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[48]) );
  XNOR2_X1 MCInst3_MC3_r0Inst_XORInst_0_0_U2  ( .A(MCInst3_MC3_v3_2 [2]), 
        .B(MCInst3_MC3_v2_0 [0]), .ZN(MCInst3_MC3_r0Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst3_MC3_r0Inst_XORInst_0_0_U1  ( .A(MCInst3_MC3_v0_3 [3]), .B(
        MCInst3_MC3_v1_0 [0]), .Z(MCInst3_MC3_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst3_MC3_r0Inst_XORInst_0_1_U3  ( .A(
        MCInst3_MC3_r0Inst_XORInst_0_1_n5 ), .B(
        MCInst3_MC3_r0Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[49]) );
  XNOR2_X1 MCInst3_MC3_r0Inst_XORInst_0_1_U2  ( .A(MCInst3_MC3_v3_0 [1]), 
        .B(MCInst3_MC3_v2_0 [1]), .ZN(MCInst3_MC3_r0Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst3_MC3_r0Inst_XORInst_0_1_U1  ( .A(MCInst3_MC3_v0_0 [1]), .B(
        MCInst3_MC3_v1_3 [2]), .Z(MCInst3_MC3_r0Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst3_MC3_r0Inst_XORInst_0_2_U3  ( .A(
        MCInst3_MC3_r0Inst_XORInst_0_2_n5 ), .B(
        MCInst3_MC3_r0Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[50]) );
  XNOR2_X1 MCInst3_MC3_r0Inst_XORInst_0_2_U2  ( .A(MCInst3_MC3_v3_0 [2]), 
        .B(MCInst3_MC3_v2_0 [2]), .ZN(MCInst3_MC3_r0Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst3_MC3_r0Inst_XORInst_0_2_U1  ( .A(MCInst3_MC3_v0_0 [2]), .B(
        Red_MCInst3_MC3_v1_1[0] ), .Z(MCInst3_MC3_r0Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst3_MC3_r0Inst_XORInst_0_3_U3  ( .A(
        MCInst3_MC3_r0Inst_XORInst_0_3_n5 ), .B(
        MCInst3_MC3_r0Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[51]) );
  XNOR2_X1 MCInst3_MC3_r0Inst_XORInst_0_3_U2  ( .A(Red_MCInst3_MC3_v3_1[0] ), 
        .B(MCInst3_MC3_v2_0 [3]), .ZN(MCInst3_MC3_r0Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst3_MC3_r0Inst_XORInst_0_3_U1  ( .A(MCInst3_MC3_v0_0 [3]), .B(
        MCInst3_MC3_v1_0 [3]), .Z(MCInst3_MC3_r0Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst3_MC3_r1Inst_XORInst_0_0_U3  ( .A(
        MCInst3_MC3_r1Inst_XORInst_0_0_n5 ), .B(
        MCInst3_MC3_r1Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[32]) );
  XNOR2_X1 MCInst3_MC3_r1Inst_XORInst_0_0_U2  ( .A(MCInst3_MC3_v3_1 [0]), 
        .B(MCInst3_MC3_v2_1 [0]), .ZN(MCInst3_MC3_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst3_MC3_r1Inst_XORInst_0_0_U1  ( .A(MCInst3_MC3_v0_0 [3]), .B(
        MCInst3_MC3_v1_1 [0]), .Z(MCInst3_MC3_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst3_MC3_r1Inst_XORInst_0_1_U3  ( .A(
        MCInst3_MC3_r1Inst_XORInst_0_1_n5 ), .B(
        MCInst3_MC3_r1Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[33]) );
  XNOR2_X1 MCInst3_MC3_r1Inst_XORInst_0_1_U2  ( .A(MCInst3_MC3_v3_1 [1]), 
        .B(MCInst3_MC3_v2_1 [1]), .ZN(MCInst3_MC3_r1Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst3_MC3_r1Inst_XORInst_0_1_U1  ( .A(MCInst3_MC3_v0_1 [1]), .B(
        MCInst3_MC3_v1_1 [1]), .Z(MCInst3_MC3_r1Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst3_MC3_r1Inst_XORInst_0_2_U3  ( .A(
        MCInst3_MC3_r1Inst_XORInst_0_2_n5 ), .B(
        MCInst3_MC3_r1Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[34]) );
  XNOR2_X1 MCInst3_MC3_r1Inst_XORInst_0_2_U2  ( .A(MCInst3_MC3_v3_1 [2]), 
        .B(MCInst3_MC3_v2_1 [2]), .ZN(MCInst3_MC3_r1Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst3_MC3_r1Inst_XORInst_0_2_U1  ( .A(MCInst3_MC3_v0_1 [2]), .B(
        MCInst3_MC3_v1_1 [2]), .Z(MCInst3_MC3_r1Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst3_MC3_r1Inst_XORInst_0_3_U3  ( .A(
        MCInst3_MC3_r1Inst_XORInst_0_3_n5 ), .B(
        MCInst3_MC3_r1Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[35]) );
  XNOR2_X1 MCInst3_MC3_r1Inst_XORInst_0_3_U2  ( .A(MCInst3_MC3_v3_1 [3]), 
        .B(MCInst3_MC3_v2_1 [3]), .ZN(MCInst3_MC3_r1Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst3_MC3_r1Inst_XORInst_0_3_U1  ( .A(MCInst3_MC3_v0_1 [3]), .B(
        MCInst3_MC3_v1_1 [3]), .Z(MCInst3_MC3_r1Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst3_MC3_r2Inst_XORInst_0_0_U3  ( .A(
        MCInst3_MC3_r2Inst_XORInst_0_0_n5 ), .B(
        MCInst3_MC3_r2Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[16]) );
  XNOR2_X1 MCInst3_MC3_r2Inst_XORInst_0_0_U2  ( .A(MCInst3_MC3_v3_2 [0]), 
        .B(MCInst3_MC3_v2_2 [0]), .ZN(MCInst3_MC3_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst3_MC3_r2Inst_XORInst_0_0_U1  ( .A(MCInst3_MC3_v0_2 [0]), .B(
        MCInst3_MC3_v1_2 [0]), .Z(MCInst3_MC3_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst3_MC3_r2Inst_XORInst_0_1_U3  ( .A(
        MCInst3_MC3_r2Inst_XORInst_0_1_n5 ), .B(
        MCInst3_MC3_r2Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[17]) );
  XNOR2_X1 MCInst3_MC3_r2Inst_XORInst_0_1_U2  ( .A(Red_MCInst3_MC3_v3_1[0] ), 
        .B(MCInst3_MC3_v2_2 [1]), .ZN(MCInst3_MC3_r2Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst3_MC3_r2Inst_XORInst_0_1_U1  ( .A(MCInst3_MC3_v0_2 [1]), .B(
        MCInst3_MC3_v1_2 [1]), .Z(MCInst3_MC3_r2Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst3_MC3_r2Inst_XORInst_0_2_U3  ( .A(
        MCInst3_MC3_r2Inst_XORInst_0_2_n5 ), .B(
        MCInst3_MC3_r2Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[18]) );
  XNOR2_X1 MCInst3_MC3_r2Inst_XORInst_0_2_U2  ( .A(MCInst3_MC3_v3_2 [2]), 
        .B(MCInst3_MC3_v2_2 [2]), .ZN(MCInst3_MC3_r2Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst3_MC3_r2Inst_XORInst_0_2_U1  ( .A(MCInst3_MC3_v0_2 [2]), .B(
        MCInst3_MC3_v1_2 [2]), .Z(MCInst3_MC3_r2Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst3_MC3_r2Inst_XORInst_0_3_U3  ( .A(
        MCInst3_MC3_r2Inst_XORInst_0_3_n5 ), .B(
        MCInst3_MC3_r2Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[19]) );
  XNOR2_X1 MCInst3_MC3_r2Inst_XORInst_0_3_U2  ( .A(MCInst3_MC3_v3_2 [3]), 
        .B(MCInst3_MC3_v2_2 [3]), .ZN(MCInst3_MC3_r2Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst3_MC3_r2Inst_XORInst_0_3_U1  ( .A(MCInst3_MC3_v0_2 [3]), .B(
        MCInst3_MC3_v1_2 [3]), .Z(MCInst3_MC3_r2Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst3_MC3_r3Inst_XORInst_0_0_U3  ( .A(
        MCInst3_MC3_r3Inst_XORInst_0_0_n5 ), .B(
        MCInst3_MC3_r3Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[0]) );
  XNOR2_X1 MCInst3_MC3_r3Inst_XORInst_0_0_U2  ( .A(MCInst3_MC3_v3_3 [0]), 
        .B(MCInst3_MC3_v2_3 [0]), .ZN(MCInst3_MC3_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst3_MC3_r3Inst_XORInst_0_0_U1  ( .A(MCInst3_MC3_v0_3 [0]), .B(
        MCInst3_MC3_v1_0 [3]), .Z(MCInst3_MC3_r3Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst3_MC3_r3Inst_XORInst_0_1_U3  ( .A(
        MCInst3_MC3_r3Inst_XORInst_0_1_n5 ), .B(
        MCInst3_MC3_r3Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[1]) );
  XNOR2_X1 MCInst3_MC3_r3Inst_XORInst_0_1_U2  ( .A(MCInst3_MC3_v3_3 [1]), 
        .B(MCInst3_MC3_v2_3 [1]), .ZN(MCInst3_MC3_r3Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst3_MC3_r3Inst_XORInst_0_1_U1  ( .A(MCInst3_MC3_v0_3 [1]), .B(
        MCInst3_MC3_v1_3 [1]), .Z(MCInst3_MC3_r3Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst3_MC3_r3Inst_XORInst_0_2_U3  ( .A(
        MCInst3_MC3_r3Inst_XORInst_0_2_n5 ), .B(
        MCInst3_MC3_r3Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[2]) );
  XNOR2_X1 MCInst3_MC3_r3Inst_XORInst_0_2_U2  ( .A(MCInst3_MC3_v3_3 [2]), 
        .B(MCInst3_MC3_v2_3 [2]), .ZN(MCInst3_MC3_r3Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst3_MC3_r3Inst_XORInst_0_2_U1  ( .A(MCInst3_MC3_v0_0 [3]), .B(
        MCInst3_MC3_v1_3 [2]), .Z(MCInst3_MC3_r3Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst3_MC3_r3Inst_XORInst_0_3_U3  ( .A(
        MCInst3_MC3_r3Inst_XORInst_0_3_n5 ), .B(
        MCInst3_MC3_r3Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[3]) );
  XNOR2_X1 MCInst3_MC3_r3Inst_XORInst_0_3_U2  ( .A(MCInst3_MC3_v3_3 [3]), 
        .B(MCInst3_MC3_v2_3 [3]), .ZN(MCInst3_MC3_r3Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst3_MC3_r3Inst_XORInst_0_3_U1  ( .A(MCInst3_MC3_v0_3 [3]), .B(
        Red_MCInst3_MC3_v1_1[0] ), .Z(MCInst3_MC3_r3Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 Red_PlaintextInst_LFInst_0_LFInst_0_U5  ( .A(
        Red_PlaintextInst_LFInst_0_LFInst_0_n4 ), .B(
        Red_PlaintextInst_LFInst_0_LFInst_0_n3 ), .ZN(Red_Plaintext[0]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_0_LFInst_0_U4  ( .A(Plaintext[1]), .B(
        Plaintext[0]), .ZN(Red_PlaintextInst_LFInst_0_LFInst_0_n3 ) );
  XOR2_X1 Red_PlaintextInst_LFInst_0_LFInst_0_U3  ( .A(Plaintext[2]), .B(
        Plaintext[3]), .Z(Red_PlaintextInst_LFInst_0_LFInst_0_n4 ) );
  XNOR2_X1 Red_PlaintextInst_LFInst_1_LFInst_0_U5  ( .A(
        Red_PlaintextInst_LFInst_1_LFInst_0_n4 ), .B(
        Red_PlaintextInst_LFInst_1_LFInst_0_n3 ), .ZN(Red_Plaintext[1]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_1_LFInst_0_U4  ( .A(Plaintext[5]), .B(
        Plaintext[4]), .ZN(Red_PlaintextInst_LFInst_1_LFInst_0_n3 ) );
  XOR2_X1 Red_PlaintextInst_LFInst_1_LFInst_0_U3  ( .A(Plaintext[6]), .B(
        Plaintext[7]), .Z(Red_PlaintextInst_LFInst_1_LFInst_0_n4 ) );
  XNOR2_X1 Red_PlaintextInst_LFInst_2_LFInst_0_U5  ( .A(
        Red_PlaintextInst_LFInst_2_LFInst_0_n4 ), .B(
        Red_PlaintextInst_LFInst_2_LFInst_0_n3 ), .ZN(Red_Plaintext[2]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_2_LFInst_0_U4  ( .A(Plaintext[9]), .B(
        Plaintext[8]), .ZN(Red_PlaintextInst_LFInst_2_LFInst_0_n3 ) );
  XOR2_X1 Red_PlaintextInst_LFInst_2_LFInst_0_U3  ( .A(Plaintext[10]), .B(
        Plaintext[11]), .Z(Red_PlaintextInst_LFInst_2_LFInst_0_n4 ) );
  XNOR2_X1 Red_PlaintextInst_LFInst_3_LFInst_0_U5  ( .A(
        Red_PlaintextInst_LFInst_3_LFInst_0_n4 ), .B(
        Red_PlaintextInst_LFInst_3_LFInst_0_n3 ), .ZN(Red_Plaintext[3]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_3_LFInst_0_U4  ( .A(Plaintext[13]), .B(
        Plaintext[12]), .ZN(Red_PlaintextInst_LFInst_3_LFInst_0_n3 ) );
  XOR2_X1 Red_PlaintextInst_LFInst_3_LFInst_0_U3  ( .A(Plaintext[14]), .B(
        Plaintext[15]), .Z(Red_PlaintextInst_LFInst_3_LFInst_0_n4 ) );
  XNOR2_X1 Red_PlaintextInst_LFInst_4_LFInst_0_U5  ( .A(
        Red_PlaintextInst_LFInst_4_LFInst_0_n4 ), .B(
        Red_PlaintextInst_LFInst_4_LFInst_0_n3 ), .ZN(Red_Plaintext[4]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_4_LFInst_0_U4  ( .A(Plaintext[17]), .B(
        Plaintext[16]), .ZN(Red_PlaintextInst_LFInst_4_LFInst_0_n3 ) );
  XOR2_X1 Red_PlaintextInst_LFInst_4_LFInst_0_U3  ( .A(Plaintext[18]), .B(
        Plaintext[19]), .Z(Red_PlaintextInst_LFInst_4_LFInst_0_n4 ) );
  XNOR2_X1 Red_PlaintextInst_LFInst_5_LFInst_0_U5  ( .A(
        Red_PlaintextInst_LFInst_5_LFInst_0_n4 ), .B(
        Red_PlaintextInst_LFInst_5_LFInst_0_n3 ), .ZN(Red_Plaintext[5]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_5_LFInst_0_U4  ( .A(Plaintext[21]), .B(
        Plaintext[20]), .ZN(Red_PlaintextInst_LFInst_5_LFInst_0_n3 ) );
  XOR2_X1 Red_PlaintextInst_LFInst_5_LFInst_0_U3  ( .A(Plaintext[22]), .B(
        Plaintext[23]), .Z(Red_PlaintextInst_LFInst_5_LFInst_0_n4 ) );
  XNOR2_X1 Red_PlaintextInst_LFInst_6_LFInst_0_U5  ( .A(
        Red_PlaintextInst_LFInst_6_LFInst_0_n4 ), .B(
        Red_PlaintextInst_LFInst_6_LFInst_0_n3 ), .ZN(Red_Plaintext[6]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_6_LFInst_0_U4  ( .A(Plaintext[25]), .B(
        Plaintext[24]), .ZN(Red_PlaintextInst_LFInst_6_LFInst_0_n3 ) );
  XOR2_X1 Red_PlaintextInst_LFInst_6_LFInst_0_U3  ( .A(Plaintext[26]), .B(
        Plaintext[27]), .Z(Red_PlaintextInst_LFInst_6_LFInst_0_n4 ) );
  XNOR2_X1 Red_PlaintextInst_LFInst_7_LFInst_0_U5  ( .A(
        Red_PlaintextInst_LFInst_7_LFInst_0_n4 ), .B(
        Red_PlaintextInst_LFInst_7_LFInst_0_n3 ), .ZN(Red_Plaintext[7]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_7_LFInst_0_U4  ( .A(Plaintext[29]), .B(
        Plaintext[28]), .ZN(Red_PlaintextInst_LFInst_7_LFInst_0_n3 ) );
  XOR2_X1 Red_PlaintextInst_LFInst_7_LFInst_0_U3  ( .A(Plaintext[30]), .B(
        Plaintext[31]), .Z(Red_PlaintextInst_LFInst_7_LFInst_0_n4 ) );
  XNOR2_X1 Red_PlaintextInst_LFInst_8_LFInst_0_U5  ( .A(
        Red_PlaintextInst_LFInst_8_LFInst_0_n4 ), .B(
        Red_PlaintextInst_LFInst_8_LFInst_0_n3 ), .ZN(Red_Plaintext[8]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_8_LFInst_0_U4  ( .A(Plaintext[33]), .B(
        Plaintext[32]), .ZN(Red_PlaintextInst_LFInst_8_LFInst_0_n3 ) );
  XOR2_X1 Red_PlaintextInst_LFInst_8_LFInst_0_U3  ( .A(Plaintext[34]), .B(
        Plaintext[35]), .Z(Red_PlaintextInst_LFInst_8_LFInst_0_n4 ) );
  XNOR2_X1 Red_PlaintextInst_LFInst_9_LFInst_0_U5  ( .A(
        Red_PlaintextInst_LFInst_9_LFInst_0_n4 ), .B(
        Red_PlaintextInst_LFInst_9_LFInst_0_n3 ), .ZN(Red_Plaintext[9]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_9_LFInst_0_U4  ( .A(Plaintext[37]), .B(
        Plaintext[36]), .ZN(Red_PlaintextInst_LFInst_9_LFInst_0_n3 ) );
  XOR2_X1 Red_PlaintextInst_LFInst_9_LFInst_0_U3  ( .A(Plaintext[38]), .B(
        Plaintext[39]), .Z(Red_PlaintextInst_LFInst_9_LFInst_0_n4 ) );
  XNOR2_X1 Red_PlaintextInst_LFInst_10_LFInst_0_U5  ( .A(
        Red_PlaintextInst_LFInst_10_LFInst_0_n4 ), .B(
        Red_PlaintextInst_LFInst_10_LFInst_0_n3 ), .ZN(Red_Plaintext[10]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_10_LFInst_0_U4  ( .A(Plaintext[41]), .B(
        Plaintext[40]), .ZN(Red_PlaintextInst_LFInst_10_LFInst_0_n3 ) );
  XOR2_X1 Red_PlaintextInst_LFInst_10_LFInst_0_U3  ( .A(Plaintext[42]), .B(
        Plaintext[43]), .Z(Red_PlaintextInst_LFInst_10_LFInst_0_n4 ) );
  XNOR2_X1 Red_PlaintextInst_LFInst_11_LFInst_0_U5  ( .A(
        Red_PlaintextInst_LFInst_11_LFInst_0_n4 ), .B(
        Red_PlaintextInst_LFInst_11_LFInst_0_n3 ), .ZN(Red_Plaintext[11]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_11_LFInst_0_U4  ( .A(Plaintext[45]), .B(
        Plaintext[44]), .ZN(Red_PlaintextInst_LFInst_11_LFInst_0_n3 ) );
  XOR2_X1 Red_PlaintextInst_LFInst_11_LFInst_0_U3  ( .A(Plaintext[46]), .B(
        Plaintext[47]), .Z(Red_PlaintextInst_LFInst_11_LFInst_0_n4 ) );
  XNOR2_X1 Red_PlaintextInst_LFInst_12_LFInst_0_U5  ( .A(
        Red_PlaintextInst_LFInst_12_LFInst_0_n4 ), .B(
        Red_PlaintextInst_LFInst_12_LFInst_0_n3 ), .ZN(Red_Plaintext[12]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_12_LFInst_0_U4  ( .A(Plaintext[49]), .B(
        Plaintext[48]), .ZN(Red_PlaintextInst_LFInst_12_LFInst_0_n3 ) );
  XOR2_X1 Red_PlaintextInst_LFInst_12_LFInst_0_U3  ( .A(Plaintext[50]), .B(
        Plaintext[51]), .Z(Red_PlaintextInst_LFInst_12_LFInst_0_n4 ) );
  XNOR2_X1 Red_PlaintextInst_LFInst_13_LFInst_0_U5  ( .A(
        Red_PlaintextInst_LFInst_13_LFInst_0_n4 ), .B(
        Red_PlaintextInst_LFInst_13_LFInst_0_n3 ), .ZN(Red_Plaintext[13]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_13_LFInst_0_U4  ( .A(Plaintext[53]), .B(
        Plaintext[52]), .ZN(Red_PlaintextInst_LFInst_13_LFInst_0_n3 ) );
  XOR2_X1 Red_PlaintextInst_LFInst_13_LFInst_0_U3  ( .A(Plaintext[54]), .B(
        Plaintext[55]), .Z(Red_PlaintextInst_LFInst_13_LFInst_0_n4 ) );
  XNOR2_X1 Red_PlaintextInst_LFInst_14_LFInst_0_U5  ( .A(
        Red_PlaintextInst_LFInst_14_LFInst_0_n4 ), .B(
        Red_PlaintextInst_LFInst_14_LFInst_0_n3 ), .ZN(Red_Plaintext[14]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_14_LFInst_0_U4  ( .A(Plaintext[57]), .B(
        Plaintext[56]), .ZN(Red_PlaintextInst_LFInst_14_LFInst_0_n3 ) );
  XOR2_X1 Red_PlaintextInst_LFInst_14_LFInst_0_U3  ( .A(Plaintext[58]), .B(
        Plaintext[59]), .Z(Red_PlaintextInst_LFInst_14_LFInst_0_n4 ) );
  XNOR2_X1 Red_PlaintextInst_LFInst_15_LFInst_0_U5  ( .A(
        Red_PlaintextInst_LFInst_15_LFInst_0_n4 ), .B(
        Red_PlaintextInst_LFInst_15_LFInst_0_n3 ), .ZN(Red_Plaintext[15]) );
  XNOR2_X1 Red_PlaintextInst_LFInst_15_LFInst_0_U4  ( .A(Plaintext[61]), .B(
        Plaintext[60]), .ZN(Red_PlaintextInst_LFInst_15_LFInst_0_n3 ) );
  XOR2_X1 Red_PlaintextInst_LFInst_15_LFInst_0_U3  ( .A(Plaintext[62]), .B(
        Plaintext[63]), .Z(Red_PlaintextInst_LFInst_15_LFInst_0_n4 ) );
  XOR2_X1 RedAddKeyXOR_XORInst_0_0_U1  ( .A(Red_Plaintext[0]), .B(
        Red_RoundKey[0]), .Z(Red_AddRoundKeyOutput[0]) );
  XOR2_X1 RedAddKeyXOR_XORInst_1_0_U1  ( .A(Red_Plaintext[1]), .B(
        Red_RoundKey[1]), .Z(Red_AddRoundKeyOutput[1]) );
  XOR2_X1 RedAddKeyXOR_XORInst_2_0_U1  ( .A(Red_Plaintext[2]), .B(
        Red_RoundKey[2]), .Z(Red_AddRoundKeyOutput[2]) );
  XOR2_X1 RedAddKeyXOR_XORInst_3_0_U1  ( .A(Red_Plaintext[3]), .B(
        Red_RoundKey[3]), .Z(Red_AddRoundKeyOutput[3]) );
  XOR2_X1 RedAddKeyXOR_XORInst_4_0_U1  ( .A(Red_Plaintext[4]), .B(
        Red_RoundKey[4]), .Z(Red_AddRoundKeyOutput[4]) );
  XOR2_X1 RedAddKeyXOR_XORInst_5_0_U1  ( .A(Red_Plaintext[5]), .B(
        Red_RoundKey[5]), .Z(Red_AddRoundKeyOutput[5]) );
  XOR2_X1 RedAddKeyXOR_XORInst_6_0_U1  ( .A(Red_Plaintext[6]), .B(
        Red_RoundKey[6]), .Z(Red_AddRoundKeyOutput[6]) );
  XOR2_X1 RedAddKeyXOR_XORInst_7_0_U1  ( .A(Red_Plaintext[7]), .B(
        Red_RoundKey[7]), .Z(Red_AddRoundKeyOutput[7]) );
  XOR2_X1 RedAddKeyXOR_XORInst_8_0_U1  ( .A(Red_Plaintext[8]), .B(
        Red_RoundKey[8]), .Z(Red_AddRoundKeyOutput[8]) );
  XOR2_X1 RedAddKeyXOR_XORInst_9_0_U1  ( .A(Red_Plaintext[9]), .B(
        Red_RoundKey[9]), .Z(Red_AddRoundKeyOutput[9]) );
  XOR2_X1 RedAddKeyXOR_XORInst_10_0_U1  ( .A(Red_Plaintext[10]), .B(
        Red_RoundKey[10]), .Z(Red_AddRoundKeyOutput[10]) );
  XOR2_X1 RedAddKeyXOR_XORInst_11_0_U1  ( .A(Red_Plaintext[11]), .B(
        Red_RoundKey[11]), .Z(Red_AddRoundKeyOutput[11]) );
  XOR2_X1 RedAddKeyXOR_XORInst_12_0_U1  ( .A(Red_Plaintext[12]), .B(
        Red_RoundKey[12]), .Z(Red_AddRoundKeyOutput[12]) );
  XOR2_X1 RedAddKeyXOR_XORInst_13_0_U1  ( .A(Red_Plaintext[13]), .B(
        Red_RoundKey[13]), .Z(Red_AddRoundKeyOutput[13]) );
  XOR2_X1 RedAddKeyXOR_XORInst_14_0_U1  ( .A(Red_Plaintext[14]), .B(
        Red_RoundKey[14]), .Z(Red_AddRoundKeyOutput[14]) );
  XOR2_X1 RedAddKeyXOR_XORInst_15_0_U1  ( .A(Red_Plaintext[15]), .B(
        Red_RoundKey[15]), .Z(Red_AddRoundKeyOutput[15]) );
  NAND2_X1 Red_SubCellInst_LFInst_0_LFInst_0_U6  ( .A1(
        Red_SubCellInst_LFInst_0_LFInst_0_n6 ), .A2(
        Red_SubCellInst_LFInst_0_LFInst_0_n5 ), .ZN(Red_ShiftRowsOutput[3])
         );
  NAND2_X1 Red_SubCellInst_LFInst_0_LFInst_0_U5  ( .A1(AddRoundKeyOutput[3]), 
        .A2(AddRoundKeyOutput[2]), .ZN(Red_SubCellInst_LFInst_0_LFInst_0_n5 )
         );
  NAND2_X1 Red_SubCellInst_LFInst_0_LFInst_0_U4  ( .A1(AddRoundKeyOutput[0]), 
        .A2(Red_SubCellInst_LFInst_0_LFInst_0_n4 ), .ZN(
        Red_SubCellInst_LFInst_0_LFInst_0_n6 ) );
  OR2_X1 Red_SubCellInst_LFInst_0_LFInst_0_U3  ( .A1(AddRoundKeyOutput[1]), 
        .A2(AddRoundKeyOutput[3]), .ZN(Red_SubCellInst_LFInst_0_LFInst_0_n4 )
         );
  NAND2_X1 Red_SubCellInst_LFInst_1_LFInst_0_U6  ( .A1(
        Red_SubCellInst_LFInst_1_LFInst_0_n6 ), .A2(
        Red_SubCellInst_LFInst_1_LFInst_0_n5 ), .ZN(Red_ShiftRowsOutput[0])
         );
  NAND2_X1 Red_SubCellInst_LFInst_1_LFInst_0_U5  ( .A1(AddRoundKeyOutput[7]), 
        .A2(AddRoundKeyOutput[6]), .ZN(Red_SubCellInst_LFInst_1_LFInst_0_n5 )
         );
  NAND2_X1 Red_SubCellInst_LFInst_1_LFInst_0_U4  ( .A1(AddRoundKeyOutput[4]), 
        .A2(Red_SubCellInst_LFInst_1_LFInst_0_n4 ), .ZN(
        Red_SubCellInst_LFInst_1_LFInst_0_n6 ) );
  OR2_X1 Red_SubCellInst_LFInst_1_LFInst_0_U3  ( .A1(AddRoundKeyOutput[5]), 
        .A2(AddRoundKeyOutput[7]), .ZN(Red_SubCellInst_LFInst_1_LFInst_0_n4 )
         );
  NAND2_X1 Red_SubCellInst_LFInst_2_LFInst_0_U6  ( .A1(
        Red_SubCellInst_LFInst_2_LFInst_0_n6 ), .A2(
        Red_SubCellInst_LFInst_2_LFInst_0_n5 ), .ZN(Red_ShiftRowsOutput[1])
         );
  NAND2_X1 Red_SubCellInst_LFInst_2_LFInst_0_U5  ( .A1(AddRoundKeyOutput[11]), 
        .A2(AddRoundKeyOutput[10]), .ZN(Red_SubCellInst_LFInst_2_LFInst_0_n5 ) );
  NAND2_X1 Red_SubCellInst_LFInst_2_LFInst_0_U4  ( .A1(AddRoundKeyOutput[8]), 
        .A2(Red_SubCellInst_LFInst_2_LFInst_0_n4 ), .ZN(
        Red_SubCellInst_LFInst_2_LFInst_0_n6 ) );
  OR2_X1 Red_SubCellInst_LFInst_2_LFInst_0_U3  ( .A1(AddRoundKeyOutput[9]), 
        .A2(AddRoundKeyOutput[11]), .ZN(Red_SubCellInst_LFInst_2_LFInst_0_n4 ) );
  NAND2_X1 Red_SubCellInst_LFInst_3_LFInst_0_U6  ( .A1(
        Red_SubCellInst_LFInst_3_LFInst_0_n6 ), .A2(
        Red_SubCellInst_LFInst_3_LFInst_0_n5 ), .ZN(Red_ShiftRowsOutput[2])
         );
  NAND2_X1 Red_SubCellInst_LFInst_3_LFInst_0_U5  ( .A1(AddRoundKeyOutput[15]), 
        .A2(AddRoundKeyOutput[14]), .ZN(Red_SubCellInst_LFInst_3_LFInst_0_n5 ) );
  NAND2_X1 Red_SubCellInst_LFInst_3_LFInst_0_U4  ( .A1(AddRoundKeyOutput[12]), 
        .A2(Red_SubCellInst_LFInst_3_LFInst_0_n4 ), .ZN(
        Red_SubCellInst_LFInst_3_LFInst_0_n6 ) );
  OR2_X1 Red_SubCellInst_LFInst_3_LFInst_0_U3  ( .A1(AddRoundKeyOutput[13]), 
        .A2(AddRoundKeyOutput[15]), .ZN(Red_SubCellInst_LFInst_3_LFInst_0_n4 ) );
  NAND2_X1 Red_SubCellInst_LFInst_4_LFInst_0_U6  ( .A1(
        Red_SubCellInst_LFInst_4_LFInst_0_n6 ), .A2(
        Red_SubCellInst_LFInst_4_LFInst_0_n5 ), .ZN(Red_ShiftRowsOutput[6])
         );
  NAND2_X1 Red_SubCellInst_LFInst_4_LFInst_0_U5  ( .A1(AddRoundKeyOutput[19]), 
        .A2(AddRoundKeyOutput[18]), .ZN(Red_SubCellInst_LFInst_4_LFInst_0_n5 ) );
  NAND2_X1 Red_SubCellInst_LFInst_4_LFInst_0_U4  ( .A1(AddRoundKeyOutput[16]), 
        .A2(Red_SubCellInst_LFInst_4_LFInst_0_n4 ), .ZN(
        Red_SubCellInst_LFInst_4_LFInst_0_n6 ) );
  OR2_X1 Red_SubCellInst_LFInst_4_LFInst_0_U3  ( .A1(AddRoundKeyOutput[17]), 
        .A2(AddRoundKeyOutput[19]), .ZN(Red_SubCellInst_LFInst_4_LFInst_0_n4 ) );
  NAND2_X1 Red_SubCellInst_LFInst_5_LFInst_0_U6  ( .A1(
        Red_SubCellInst_LFInst_5_LFInst_0_n6 ), .A2(
        Red_SubCellInst_LFInst_5_LFInst_0_n5 ), .ZN(Red_ShiftRowsOutput[7])
         );
  NAND2_X1 Red_SubCellInst_LFInst_5_LFInst_0_U5  ( .A1(AddRoundKeyOutput[23]), 
        .A2(AddRoundKeyOutput[22]), .ZN(Red_SubCellInst_LFInst_5_LFInst_0_n5 ) );
  NAND2_X1 Red_SubCellInst_LFInst_5_LFInst_0_U4  ( .A1(AddRoundKeyOutput[20]), 
        .A2(Red_SubCellInst_LFInst_5_LFInst_0_n4 ), .ZN(
        Red_SubCellInst_LFInst_5_LFInst_0_n6 ) );
  OR2_X1 Red_SubCellInst_LFInst_5_LFInst_0_U3  ( .A1(AddRoundKeyOutput[21]), 
        .A2(AddRoundKeyOutput[23]), .ZN(Red_SubCellInst_LFInst_5_LFInst_0_n4 ) );
  NAND2_X1 Red_SubCellInst_LFInst_6_LFInst_0_U6  ( .A1(
        Red_SubCellInst_LFInst_6_LFInst_0_n6 ), .A2(
        Red_SubCellInst_LFInst_6_LFInst_0_n5 ), .ZN(Red_ShiftRowsOutput[4])
         );
  NAND2_X1 Red_SubCellInst_LFInst_6_LFInst_0_U5  ( .A1(AddRoundKeyOutput[27]), 
        .A2(AddRoundKeyOutput[26]), .ZN(Red_SubCellInst_LFInst_6_LFInst_0_n5 ) );
  NAND2_X1 Red_SubCellInst_LFInst_6_LFInst_0_U4  ( .A1(AddRoundKeyOutput[24]), 
        .A2(Red_SubCellInst_LFInst_6_LFInst_0_n4 ), .ZN(
        Red_SubCellInst_LFInst_6_LFInst_0_n6 ) );
  OR2_X1 Red_SubCellInst_LFInst_6_LFInst_0_U3  ( .A1(AddRoundKeyOutput[25]), 
        .A2(AddRoundKeyOutput[27]), .ZN(Red_SubCellInst_LFInst_6_LFInst_0_n4 ) );
  NAND2_X1 Red_SubCellInst_LFInst_7_LFInst_0_U6  ( .A1(
        Red_SubCellInst_LFInst_7_LFInst_0_n6 ), .A2(
        Red_SubCellInst_LFInst_7_LFInst_0_n5 ), .ZN(Red_ShiftRowsOutput[5])
         );
  NAND2_X1 Red_SubCellInst_LFInst_7_LFInst_0_U5  ( .A1(AddRoundKeyOutput[31]), 
        .A2(AddRoundKeyOutput[30]), .ZN(Red_SubCellInst_LFInst_7_LFInst_0_n5 ) );
  NAND2_X1 Red_SubCellInst_LFInst_7_LFInst_0_U4  ( .A1(AddRoundKeyOutput[28]), 
        .A2(Red_SubCellInst_LFInst_7_LFInst_0_n4 ), .ZN(
        Red_SubCellInst_LFInst_7_LFInst_0_n6 ) );
  OR2_X1 Red_SubCellInst_LFInst_7_LFInst_0_U3  ( .A1(AddRoundKeyOutput[29]), 
        .A2(AddRoundKeyOutput[31]), .ZN(Red_SubCellInst_LFInst_7_LFInst_0_n4 ) );
  NAND2_X1 Red_SubCellInst_LFInst_8_LFInst_0_U6  ( .A1(
        Red_SubCellInst_LFInst_8_LFInst_0_n6 ), .A2(
        Red_SubCellInst_LFInst_8_LFInst_0_n5 ), .ZN(Red_ShiftRowsOutput[9])
         );
  NAND2_X1 Red_SubCellInst_LFInst_8_LFInst_0_U5  ( .A1(AddRoundKeyOutput[35]), 
        .A2(AddRoundKeyOutput[34]), .ZN(Red_SubCellInst_LFInst_8_LFInst_0_n5 ) );
  NAND2_X1 Red_SubCellInst_LFInst_8_LFInst_0_U4  ( .A1(AddRoundKeyOutput[32]), 
        .A2(Red_SubCellInst_LFInst_8_LFInst_0_n4 ), .ZN(
        Red_SubCellInst_LFInst_8_LFInst_0_n6 ) );
  OR2_X1 Red_SubCellInst_LFInst_8_LFInst_0_U3  ( .A1(AddRoundKeyOutput[33]), 
        .A2(AddRoundKeyOutput[35]), .ZN(Red_SubCellInst_LFInst_8_LFInst_0_n4 ) );
  NAND2_X1 Red_SubCellInst_LFInst_9_LFInst_0_U6  ( .A1(
        Red_SubCellInst_LFInst_9_LFInst_0_n6 ), .A2(
        Red_SubCellInst_LFInst_9_LFInst_0_n5 ), .ZN(Red_ShiftRowsOutput[10])
         );
  NAND2_X1 Red_SubCellInst_LFInst_9_LFInst_0_U5  ( .A1(AddRoundKeyOutput[39]), 
        .A2(AddRoundKeyOutput[38]), .ZN(Red_SubCellInst_LFInst_9_LFInst_0_n5 ) );
  NAND2_X1 Red_SubCellInst_LFInst_9_LFInst_0_U4  ( .A1(AddRoundKeyOutput[36]), 
        .A2(Red_SubCellInst_LFInst_9_LFInst_0_n4 ), .ZN(
        Red_SubCellInst_LFInst_9_LFInst_0_n6 ) );
  OR2_X1 Red_SubCellInst_LFInst_9_LFInst_0_U3  ( .A1(AddRoundKeyOutput[37]), 
        .A2(AddRoundKeyOutput[39]), .ZN(Red_SubCellInst_LFInst_9_LFInst_0_n4 ) );
  NAND2_X1 Red_SubCellInst_LFInst_10_LFInst_0_U6  ( .A1(
        Red_SubCellInst_LFInst_10_LFInst_0_n6 ), .A2(
        Red_SubCellInst_LFInst_10_LFInst_0_n5 ), .ZN(Red_ShiftRowsOutput[11])
         );
  NAND2_X1 Red_SubCellInst_LFInst_10_LFInst_0_U5  ( .A1(AddRoundKeyOutput[43]), .A2(AddRoundKeyOutput[42]), .ZN(Red_SubCellInst_LFInst_10_LFInst_0_n5 ) );
  NAND2_X1 Red_SubCellInst_LFInst_10_LFInst_0_U4  ( .A1(AddRoundKeyOutput[40]), .A2(Red_SubCellInst_LFInst_10_LFInst_0_n4 ), .ZN(
        Red_SubCellInst_LFInst_10_LFInst_0_n6 ) );
  OR2_X1 Red_SubCellInst_LFInst_10_LFInst_0_U3  ( .A1(AddRoundKeyOutput[41]), 
        .A2(AddRoundKeyOutput[43]), .ZN(
        Red_SubCellInst_LFInst_10_LFInst_0_n4 ) );
  NAND2_X1 Red_SubCellInst_LFInst_11_LFInst_0_U6  ( .A1(
        Red_SubCellInst_LFInst_11_LFInst_0_n6 ), .A2(
        Red_SubCellInst_LFInst_11_LFInst_0_n5 ), .ZN(Red_ShiftRowsOutput[8])
         );
  NAND2_X1 Red_SubCellInst_LFInst_11_LFInst_0_U5  ( .A1(AddRoundKeyOutput[47]), .A2(AddRoundKeyOutput[46]), .ZN(Red_SubCellInst_LFInst_11_LFInst_0_n5 ) );
  NAND2_X1 Red_SubCellInst_LFInst_11_LFInst_0_U4  ( .A1(AddRoundKeyOutput[44]), .A2(Red_SubCellInst_LFInst_11_LFInst_0_n4 ), .ZN(
        Red_SubCellInst_LFInst_11_LFInst_0_n6 ) );
  OR2_X1 Red_SubCellInst_LFInst_11_LFInst_0_U3  ( .A1(AddRoundKeyOutput[45]), 
        .A2(AddRoundKeyOutput[47]), .ZN(
        Red_SubCellInst_LFInst_11_LFInst_0_n4 ) );
  NAND2_X1 Red_SubCellInst_LFInst_12_LFInst_0_U6  ( .A1(
        Red_SubCellInst_LFInst_12_LFInst_0_n6 ), .A2(
        Red_SubCellInst_LFInst_12_LFInst_0_n5 ), .ZN(Red_ShiftRowsOutput[12])
         );
  NAND2_X1 Red_SubCellInst_LFInst_12_LFInst_0_U5  ( .A1(AddRoundKeyOutput[51]), .A2(AddRoundKeyOutput[50]), .ZN(Red_SubCellInst_LFInst_12_LFInst_0_n5 ) );
  NAND2_X1 Red_SubCellInst_LFInst_12_LFInst_0_U4  ( .A1(AddRoundKeyOutput[48]), .A2(Red_SubCellInst_LFInst_12_LFInst_0_n4 ), .ZN(
        Red_SubCellInst_LFInst_12_LFInst_0_n6 ) );
  OR2_X1 Red_SubCellInst_LFInst_12_LFInst_0_U3  ( .A1(AddRoundKeyOutput[49]), 
        .A2(AddRoundKeyOutput[51]), .ZN(
        Red_SubCellInst_LFInst_12_LFInst_0_n4 ) );
  NAND2_X1 Red_SubCellInst_LFInst_13_LFInst_0_U6  ( .A1(
        Red_SubCellInst_LFInst_13_LFInst_0_n6 ), .A2(
        Red_SubCellInst_LFInst_13_LFInst_0_n5 ), .ZN(Red_ShiftRowsOutput[13])
         );
  NAND2_X1 Red_SubCellInst_LFInst_13_LFInst_0_U5  ( .A1(AddRoundKeyOutput[55]), .A2(AddRoundKeyOutput[54]), .ZN(Red_SubCellInst_LFInst_13_LFInst_0_n5 ) );
  NAND2_X1 Red_SubCellInst_LFInst_13_LFInst_0_U4  ( .A1(AddRoundKeyOutput[52]), .A2(Red_SubCellInst_LFInst_13_LFInst_0_n4 ), .ZN(
        Red_SubCellInst_LFInst_13_LFInst_0_n6 ) );
  OR2_X1 Red_SubCellInst_LFInst_13_LFInst_0_U3  ( .A1(AddRoundKeyOutput[53]), 
        .A2(AddRoundKeyOutput[55]), .ZN(
        Red_SubCellInst_LFInst_13_LFInst_0_n4 ) );
  NAND2_X1 Red_SubCellInst_LFInst_14_LFInst_0_U6  ( .A1(
        Red_SubCellInst_LFInst_14_LFInst_0_n6 ), .A2(
        Red_SubCellInst_LFInst_14_LFInst_0_n5 ), .ZN(Red_ShiftRowsOutput[14])
         );
  NAND2_X1 Red_SubCellInst_LFInst_14_LFInst_0_U5  ( .A1(AddRoundKeyOutput[59]), .A2(AddRoundKeyOutput[58]), .ZN(Red_SubCellInst_LFInst_14_LFInst_0_n5 ) );
  NAND2_X1 Red_SubCellInst_LFInst_14_LFInst_0_U4  ( .A1(AddRoundKeyOutput[56]), .A2(Red_SubCellInst_LFInst_14_LFInst_0_n4 ), .ZN(
        Red_SubCellInst_LFInst_14_LFInst_0_n6 ) );
  OR2_X1 Red_SubCellInst_LFInst_14_LFInst_0_U3  ( .A1(AddRoundKeyOutput[57]), 
        .A2(AddRoundKeyOutput[59]), .ZN(
        Red_SubCellInst_LFInst_14_LFInst_0_n4 ) );
  NAND2_X1 Red_SubCellInst_LFInst_15_LFInst_0_U6  ( .A1(
        Red_SubCellInst_LFInst_15_LFInst_0_n6 ), .A2(
        Red_SubCellInst_LFInst_15_LFInst_0_n5 ), .ZN(Red_ShiftRowsOutput[15])
         );
  NAND2_X1 Red_SubCellInst_LFInst_15_LFInst_0_U5  ( .A1(AddRoundKeyOutput[63]), .A2(AddRoundKeyOutput[62]), .ZN(Red_SubCellInst_LFInst_15_LFInst_0_n5 ) );
  NAND2_X1 Red_SubCellInst_LFInst_15_LFInst_0_U4  ( .A1(AddRoundKeyOutput[60]), .A2(Red_SubCellInst_LFInst_15_LFInst_0_n4 ), .ZN(
        Red_SubCellInst_LFInst_15_LFInst_0_n6 ) );
  OR2_X1 Red_SubCellInst_LFInst_15_LFInst_0_U3  ( .A1(AddRoundKeyOutput[61]), 
        .A2(AddRoundKeyOutput[63]), .ZN(
        Red_SubCellInst_LFInst_15_LFInst_0_n4 ) );
  XOR2_X1 Red_MCInst_MC0_v0_0Inst_0_U3  ( .A(Red_MCInst_MC0_v0_1[0] ), .B(
        MCInst_MC0_v0_0 [3]), .Z(Red_MCInst_MC0_v0_0[0] ) );
  XOR2_X1 Red_MCInst_MC0_v0_2Inst_0_U3  ( .A(Red_MCInst_MC0_v0_1[0] ), .B(
        MCInst_MC0_v0_3 [0]), .Z(Red_MCInst_MC0_v0_2[0] ) );
  XNOR2_X1 Red_MCInst_MC0_v0_3Inst_0_U4  ( .A(Red_MCInst_MC0_v0_3Inst_0_n2 ), 
        .B(MCInst_MC0_v0_0 [3]), .ZN(Red_MCInst_MC0_v0_3[0] ) );
  XNOR2_X1 Red_MCInst_MC0_v0_3Inst_0_U3  ( .A(MCInst_MC0_v0_3 [3]), .B(
        Red_MCInst_MC0_v0_1[0] ), .ZN(Red_MCInst_MC0_v0_3Inst_0_n2 ) );
  XNOR2_X1 Red_MCInst_MC0_v1_0Inst_0_U5  ( .A(Red_MCInst_MC0_v1_0Inst_0_n4 ), 
        .B(Red_MCInst_MC0_v1_0Inst_0_n3 ), .ZN(Red_MCInst_MC0_v1_0[0] ) );
  XNOR2_X1 Red_MCInst_MC0_v1_0Inst_0_U4  ( .A(MCInst_MC0_v1_3 [2]), .B(
        MCInst_MC0_v1_0 [0]), .ZN(Red_MCInst_MC0_v1_0Inst_0_n3 ) );
  XOR2_X1 Red_MCInst_MC0_v1_0Inst_0_U3  ( .A(Red_MCInst_MC0_v1_1[0] ), .B(
        MCInst_MC0_v1_0 [3]), .Z(Red_MCInst_MC0_v1_0Inst_0_n4 ) );
  XOR2_X1 Red_MCInst_MC0_v1_2Inst_0_U3  ( .A(MCInst_MC0_v1_0 [0]), .B(
        Red_MCInst_MC0_v1_1[0] ), .Z(Red_MCInst_MC0_v1_2[0] ) );
  XNOR2_X1 Red_MCInst_MC0_v1_3Inst_0_U4  ( .A(Red_MCInst_MC0_v1_3Inst_0_n2 ), 
        .B(MCInst_MC0_v1_3 [2]), .ZN(Red_MCInst_MC0_v1_3[0] ) );
  XNOR2_X1 Red_MCInst_MC0_v1_3Inst_0_U3  ( .A(Red_MCInst_MC0_v1_1[0] ), .B(
        MCInst_MC0_v1_0 [0]), .ZN(Red_MCInst_MC0_v1_3Inst_0_n2 ) );
  XNOR2_X1 Red_MCInst_MC0_v2_0Inst_0_U4  ( .A(Red_MCInst_MC0_v2_0Inst_0_n2 ), 
        .B(MCInst_MC0_v2_0 [2]), .ZN(Red_MCInst_MC0_v2_0[0] ) );
  XNOR2_X1 Red_MCInst_MC0_v2_0Inst_0_U3  ( .A(MCInst_MC0_v2_0 [3]), .B(
        MCInst_MC0_v2_3 [1]), .ZN(Red_MCInst_MC0_v2_0Inst_0_n2 ) );
  XOR2_X1 Red_MCInst_MC0_v2_1Inst_0_U3  ( .A(MCInst_MC0_v2_0 [3]), .B(
        MCInst_MC0_v2_0 [0]), .Z(Red_MCInst_MC0_v2_1[0] ) );
  XOR2_X1 Red_MCInst_MC0_v2_2Inst_0_U3  ( .A(MCInst_MC0_v2_0 [2]), .B(
        MCInst_MC0_v2_0 [3]), .Z(Red_MCInst_MC0_v2_2[0] ) );
  XOR2_X1 Red_MCInst_MC0_v2_3Inst_0_U3  ( .A(MCInst_MC0_v2_0 [2]), .B(
        MCInst_MC0_v2_0 [0]), .Z(Red_MCInst_MC0_v2_3[0] ) );
  XNOR2_X1 Red_MCInst_MC0_v3_0Inst_0_U4  ( .A(Red_MCInst_MC0_v3_0Inst_0_n2 ), 
        .B(MCInst_MC0_v3_0 [2]), .ZN(Red_MCInst_MC0_v3_0[0] ) );
  XNOR2_X1 Red_MCInst_MC0_v3_0Inst_0_U3  ( .A(Red_MCInst_MC0_v3_1[0] ), .B(
        MCInst_MC0_v3_2 [3]), .ZN(Red_MCInst_MC0_v3_0Inst_0_n2 ) );
  XNOR2_X1 Red_MCInst_MC0_v3_2Inst_0_U4  ( .A(Red_MCInst_MC0_v3_2Inst_0_n2 ), 
        .B(Red_MCInst_MC0_v3_1[0] ), .ZN(Red_MCInst_MC0_v3_2[0] ) );
  XNOR2_X1 Red_MCInst_MC0_v3_2Inst_0_U3  ( .A(MCInst_MC0_v3_2 [2]), .B(
        MCInst_MC0_v3_0 [2]), .ZN(Red_MCInst_MC0_v3_2Inst_0_n2 ) );
  XOR2_X1 Red_MCInst_MC0_v3_3Inst_0_U3  ( .A(MCInst_MC0_v3_2 [3]), .B(
        MCInst_MC0_v3_2 [2]), .Z(Red_MCInst_MC0_v3_3[0] ) );
  XNOR2_X1 Red_MCInst_MC0_r0Inst_XORInst_0_0_U3  ( .A(
        Red_MCInst_MC0_r0Inst_XORInst_0_0_n5 ), .B(
        Red_MCInst_MC0_r0Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback[15]) );
  XNOR2_X1 Red_MCInst_MC0_r0Inst_XORInst_0_0_U2  ( .A(
        Red_MCInst_MC0_v3_0[0] ), .B(Red_MCInst_MC0_v2_0[0] ), .ZN(
        Red_MCInst_MC0_r0Inst_XORInst_0_0_n4 ) );
  XOR2_X1 Red_MCInst_MC0_r0Inst_XORInst_0_0_U1  ( .A(Red_MCInst_MC0_v0_0[0] ), .B(Red_MCInst_MC0_v1_0[0] ), .Z(Red_MCInst_MC0_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 Red_MCInst_MC0_r1Inst_XORInst_0_0_U3  ( .A(
        Red_MCInst_MC0_r1Inst_XORInst_0_0_n5 ), .B(
        Red_MCInst_MC0_r1Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback[11]) );
  XNOR2_X1 Red_MCInst_MC0_r1Inst_XORInst_0_0_U2  ( .A(
        Red_MCInst_MC0_v3_1[0] ), .B(Red_MCInst_MC0_v2_1[0] ), .ZN(
        Red_MCInst_MC0_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 Red_MCInst_MC0_r1Inst_XORInst_0_0_U1  ( .A(Red_MCInst_MC0_v0_1[0] ), .B(Red_MCInst_MC0_v1_1[0] ), .Z(Red_MCInst_MC0_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 Red_MCInst_MC0_r2Inst_XORInst_0_0_U3  ( .A(
        Red_MCInst_MC0_r2Inst_XORInst_0_0_n5 ), .B(
        Red_MCInst_MC0_r2Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback[7]) );
  XNOR2_X1 Red_MCInst_MC0_r2Inst_XORInst_0_0_U2  ( .A(
        Red_MCInst_MC0_v3_2[0] ), .B(Red_MCInst_MC0_v2_2[0] ), .ZN(
        Red_MCInst_MC0_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 Red_MCInst_MC0_r2Inst_XORInst_0_0_U1  ( .A(Red_MCInst_MC0_v0_2[0] ), .B(Red_MCInst_MC0_v1_2[0] ), .Z(Red_MCInst_MC0_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 Red_MCInst_MC0_r3Inst_XORInst_0_0_U3  ( .A(
        Red_MCInst_MC0_r3Inst_XORInst_0_0_n5 ), .B(
        Red_MCInst_MC0_r3Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback[3]) );
  XNOR2_X1 Red_MCInst_MC0_r3Inst_XORInst_0_0_U2  ( .A(
        Red_MCInst_MC0_v3_3[0] ), .B(Red_MCInst_MC0_v2_3[0] ), .ZN(
        Red_MCInst_MC0_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 Red_MCInst_MC0_r3Inst_XORInst_0_0_U1  ( .A(Red_MCInst_MC0_v0_3[0] ), .B(Red_MCInst_MC0_v1_3[0] ), .Z(Red_MCInst_MC0_r3Inst_XORInst_0_0_n5 ) );
  XOR2_X1 Red_MCInst_MC1_v0_0Inst_0_U3  ( .A(Red_MCInst_MC1_v0_1[0] ), .B(
        MCInst_MC1_v0_0 [3]), .Z(Red_MCInst_MC1_v0_0[0] ) );
  XOR2_X1 Red_MCInst_MC1_v0_2Inst_0_U3  ( .A(Red_MCInst_MC1_v0_1[0] ), .B(
        MCInst_MC1_v0_3 [0]), .Z(Red_MCInst_MC1_v0_2[0] ) );
  XNOR2_X1 Red_MCInst_MC1_v0_3Inst_0_U4  ( .A(Red_MCInst_MC1_v0_3Inst_0_n2 ), 
        .B(MCInst_MC1_v0_0 [3]), .ZN(Red_MCInst_MC1_v0_3[0] ) );
  XNOR2_X1 Red_MCInst_MC1_v0_3Inst_0_U3  ( .A(MCInst_MC1_v0_3 [3]), .B(
        Red_MCInst_MC1_v0_1[0] ), .ZN(Red_MCInst_MC1_v0_3Inst_0_n2 ) );
  XNOR2_X1 Red_MCInst_MC1_v1_0Inst_0_U5  ( .A(Red_MCInst_MC1_v1_0Inst_0_n4 ), 
        .B(Red_MCInst_MC1_v1_0Inst_0_n3 ), .ZN(Red_MCInst_MC1_v1_0[0] ) );
  XNOR2_X1 Red_MCInst_MC1_v1_0Inst_0_U4  ( .A(MCInst_MC1_v1_3 [2]), .B(
        MCInst_MC1_v1_0 [0]), .ZN(Red_MCInst_MC1_v1_0Inst_0_n3 ) );
  XOR2_X1 Red_MCInst_MC1_v1_0Inst_0_U3  ( .A(Red_MCInst_MC1_v1_1[0] ), .B(
        MCInst_MC1_v1_0 [3]), .Z(Red_MCInst_MC1_v1_0Inst_0_n4 ) );
  XOR2_X1 Red_MCInst_MC1_v1_2Inst_0_U3  ( .A(MCInst_MC1_v1_0 [0]), .B(
        Red_MCInst_MC1_v1_1[0] ), .Z(Red_MCInst_MC1_v1_2[0] ) );
  XNOR2_X1 Red_MCInst_MC1_v1_3Inst_0_U4  ( .A(Red_MCInst_MC1_v1_3Inst_0_n2 ), 
        .B(MCInst_MC1_v1_3 [2]), .ZN(Red_MCInst_MC1_v1_3[0] ) );
  XNOR2_X1 Red_MCInst_MC1_v1_3Inst_0_U3  ( .A(Red_MCInst_MC1_v1_1[0] ), .B(
        MCInst_MC1_v1_0 [0]), .ZN(Red_MCInst_MC1_v1_3Inst_0_n2 ) );
  XNOR2_X1 Red_MCInst_MC1_v2_0Inst_0_U4  ( .A(Red_MCInst_MC1_v2_0Inst_0_n2 ), 
        .B(MCInst_MC1_v2_0 [2]), .ZN(Red_MCInst_MC1_v2_0[0] ) );
  XNOR2_X1 Red_MCInst_MC1_v2_0Inst_0_U3  ( .A(MCInst_MC1_v2_0 [3]), .B(
        MCInst_MC1_v2_3 [1]), .ZN(Red_MCInst_MC1_v2_0Inst_0_n2 ) );
  XOR2_X1 Red_MCInst_MC1_v2_1Inst_0_U3  ( .A(MCInst_MC1_v2_0 [3]), .B(
        MCInst_MC1_v2_0 [0]), .Z(Red_MCInst_MC1_v2_1[0] ) );
  XOR2_X1 Red_MCInst_MC1_v2_2Inst_0_U3  ( .A(MCInst_MC1_v2_0 [2]), .B(
        MCInst_MC1_v2_0 [3]), .Z(Red_MCInst_MC1_v2_2[0] ) );
  XOR2_X1 Red_MCInst_MC1_v2_3Inst_0_U3  ( .A(MCInst_MC1_v2_0 [2]), .B(
        MCInst_MC1_v2_0 [0]), .Z(Red_MCInst_MC1_v2_3[0] ) );
  XNOR2_X1 Red_MCInst_MC1_v3_0Inst_0_U4  ( .A(Red_MCInst_MC1_v3_0Inst_0_n2 ), 
        .B(MCInst_MC1_v3_0 [2]), .ZN(Red_MCInst_MC1_v3_0[0] ) );
  XNOR2_X1 Red_MCInst_MC1_v3_0Inst_0_U3  ( .A(Red_MCInst_MC1_v3_1[0] ), .B(
        MCInst_MC1_v3_2 [3]), .ZN(Red_MCInst_MC1_v3_0Inst_0_n2 ) );
  XNOR2_X1 Red_MCInst_MC1_v3_2Inst_0_U4  ( .A(Red_MCInst_MC1_v3_2Inst_0_n2 ), 
        .B(Red_MCInst_MC1_v3_1[0] ), .ZN(Red_MCInst_MC1_v3_2[0] ) );
  XNOR2_X1 Red_MCInst_MC1_v3_2Inst_0_U3  ( .A(MCInst_MC1_v3_2 [2]), .B(
        MCInst_MC1_v3_0 [2]), .ZN(Red_MCInst_MC1_v3_2Inst_0_n2 ) );
  XOR2_X1 Red_MCInst_MC1_v3_3Inst_0_U3  ( .A(MCInst_MC1_v3_2 [3]), .B(
        MCInst_MC1_v3_2 [2]), .Z(Red_MCInst_MC1_v3_3[0] ) );
  XNOR2_X1 Red_MCInst_MC1_r0Inst_XORInst_0_0_U3  ( .A(
        Red_MCInst_MC1_r0Inst_XORInst_0_0_n5 ), .B(
        Red_MCInst_MC1_r0Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback[14]) );
  XNOR2_X1 Red_MCInst_MC1_r0Inst_XORInst_0_0_U2  ( .A(
        Red_MCInst_MC1_v3_0[0] ), .B(Red_MCInst_MC1_v2_0[0] ), .ZN(
        Red_MCInst_MC1_r0Inst_XORInst_0_0_n4 ) );
  XOR2_X1 Red_MCInst_MC1_r0Inst_XORInst_0_0_U1  ( .A(Red_MCInst_MC1_v0_0[0] ), .B(Red_MCInst_MC1_v1_0[0] ), .Z(Red_MCInst_MC1_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 Red_MCInst_MC1_r1Inst_XORInst_0_0_U3  ( .A(
        Red_MCInst_MC1_r1Inst_XORInst_0_0_n5 ), .B(
        Red_MCInst_MC1_r1Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback[10]) );
  XNOR2_X1 Red_MCInst_MC1_r1Inst_XORInst_0_0_U2  ( .A(
        Red_MCInst_MC1_v3_1[0] ), .B(Red_MCInst_MC1_v2_1[0] ), .ZN(
        Red_MCInst_MC1_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 Red_MCInst_MC1_r1Inst_XORInst_0_0_U1  ( .A(Red_MCInst_MC1_v0_1[0] ), .B(Red_MCInst_MC1_v1_1[0] ), .Z(Red_MCInst_MC1_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 Red_MCInst_MC1_r2Inst_XORInst_0_0_U3  ( .A(
        Red_MCInst_MC1_r2Inst_XORInst_0_0_n5 ), .B(
        Red_MCInst_MC1_r2Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback[6]) );
  XNOR2_X1 Red_MCInst_MC1_r2Inst_XORInst_0_0_U2  ( .A(
        Red_MCInst_MC1_v3_2[0] ), .B(Red_MCInst_MC1_v2_2[0] ), .ZN(
        Red_MCInst_MC1_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 Red_MCInst_MC1_r2Inst_XORInst_0_0_U1  ( .A(Red_MCInst_MC1_v0_2[0] ), .B(Red_MCInst_MC1_v1_2[0] ), .Z(Red_MCInst_MC1_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 Red_MCInst_MC1_r3Inst_XORInst_0_0_U3  ( .A(
        Red_MCInst_MC1_r3Inst_XORInst_0_0_n5 ), .B(
        Red_MCInst_MC1_r3Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback[2]) );
  XNOR2_X1 Red_MCInst_MC1_r3Inst_XORInst_0_0_U2  ( .A(
        Red_MCInst_MC1_v3_3[0] ), .B(Red_MCInst_MC1_v2_3[0] ), .ZN(
        Red_MCInst_MC1_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 Red_MCInst_MC1_r3Inst_XORInst_0_0_U1  ( .A(Red_MCInst_MC1_v0_3[0] ), .B(Red_MCInst_MC1_v1_3[0] ), .Z(Red_MCInst_MC1_r3Inst_XORInst_0_0_n5 ) );
  XOR2_X1 Red_MCInst_MC2_v0_0Inst_0_U3  ( .A(Red_MCInst_MC2_v0_1[0] ), .B(
        MCInst_MC2_v0_0 [3]), .Z(Red_MCInst_MC2_v0_0[0] ) );
  XOR2_X1 Red_MCInst_MC2_v0_2Inst_0_U3  ( .A(Red_MCInst_MC2_v0_1[0] ), .B(
        MCInst_MC2_v0_3 [0]), .Z(Red_MCInst_MC2_v0_2[0] ) );
  XNOR2_X1 Red_MCInst_MC2_v0_3Inst_0_U4  ( .A(Red_MCInst_MC2_v0_3Inst_0_n2 ), 
        .B(MCInst_MC2_v0_0 [3]), .ZN(Red_MCInst_MC2_v0_3[0] ) );
  XNOR2_X1 Red_MCInst_MC2_v0_3Inst_0_U3  ( .A(MCInst_MC2_v0_3 [3]), .B(
        Red_MCInst_MC2_v0_1[0] ), .ZN(Red_MCInst_MC2_v0_3Inst_0_n2 ) );
  XNOR2_X1 Red_MCInst_MC2_v1_0Inst_0_U5  ( .A(Red_MCInst_MC2_v1_0Inst_0_n4 ), 
        .B(Red_MCInst_MC2_v1_0Inst_0_n3 ), .ZN(Red_MCInst_MC2_v1_0[0] ) );
  XNOR2_X1 Red_MCInst_MC2_v1_0Inst_0_U4  ( .A(MCInst_MC2_v1_3 [2]), .B(
        MCInst_MC2_v1_0 [0]), .ZN(Red_MCInst_MC2_v1_0Inst_0_n3 ) );
  XOR2_X1 Red_MCInst_MC2_v1_0Inst_0_U3  ( .A(Red_MCInst_MC2_v1_1[0] ), .B(
        MCInst_MC2_v1_0 [3]), .Z(Red_MCInst_MC2_v1_0Inst_0_n4 ) );
  XOR2_X1 Red_MCInst_MC2_v1_2Inst_0_U3  ( .A(MCInst_MC2_v1_0 [0]), .B(
        Red_MCInst_MC2_v1_1[0] ), .Z(Red_MCInst_MC2_v1_2[0] ) );
  XNOR2_X1 Red_MCInst_MC2_v1_3Inst_0_U4  ( .A(Red_MCInst_MC2_v1_3Inst_0_n2 ), 
        .B(MCInst_MC2_v1_3 [2]), .ZN(Red_MCInst_MC2_v1_3[0] ) );
  XNOR2_X1 Red_MCInst_MC2_v1_3Inst_0_U3  ( .A(Red_MCInst_MC2_v1_1[0] ), .B(
        MCInst_MC2_v1_0 [0]), .ZN(Red_MCInst_MC2_v1_3Inst_0_n2 ) );
  XNOR2_X1 Red_MCInst_MC2_v2_0Inst_0_U4  ( .A(Red_MCInst_MC2_v2_0Inst_0_n2 ), 
        .B(MCInst_MC2_v2_0 [2]), .ZN(Red_MCInst_MC2_v2_0[0] ) );
  XNOR2_X1 Red_MCInst_MC2_v2_0Inst_0_U3  ( .A(MCInst_MC2_v2_0 [3]), .B(
        MCInst_MC2_v2_3 [1]), .ZN(Red_MCInst_MC2_v2_0Inst_0_n2 ) );
  XOR2_X1 Red_MCInst_MC2_v2_1Inst_0_U3  ( .A(MCInst_MC2_v2_0 [3]), .B(
        MCInst_MC2_v2_0 [0]), .Z(Red_MCInst_MC2_v2_1[0] ) );
  XOR2_X1 Red_MCInst_MC2_v2_2Inst_0_U3  ( .A(MCInst_MC2_v2_0 [2]), .B(
        MCInst_MC2_v2_0 [3]), .Z(Red_MCInst_MC2_v2_2[0] ) );
  XOR2_X1 Red_MCInst_MC2_v2_3Inst_0_U3  ( .A(MCInst_MC2_v2_0 [2]), .B(
        MCInst_MC2_v2_0 [0]), .Z(Red_MCInst_MC2_v2_3[0] ) );
  XNOR2_X1 Red_MCInst_MC2_v3_0Inst_0_U4  ( .A(Red_MCInst_MC2_v3_0Inst_0_n2 ), 
        .B(MCInst_MC2_v3_0 [2]), .ZN(Red_MCInst_MC2_v3_0[0] ) );
  XNOR2_X1 Red_MCInst_MC2_v3_0Inst_0_U3  ( .A(Red_MCInst_MC2_v3_1[0] ), .B(
        MCInst_MC2_v3_2 [3]), .ZN(Red_MCInst_MC2_v3_0Inst_0_n2 ) );
  XNOR2_X1 Red_MCInst_MC2_v3_2Inst_0_U4  ( .A(Red_MCInst_MC2_v3_2Inst_0_n2 ), 
        .B(Red_MCInst_MC2_v3_1[0] ), .ZN(Red_MCInst_MC2_v3_2[0] ) );
  XNOR2_X1 Red_MCInst_MC2_v3_2Inst_0_U3  ( .A(MCInst_MC2_v3_2 [2]), .B(
        MCInst_MC2_v3_0 [2]), .ZN(Red_MCInst_MC2_v3_2Inst_0_n2 ) );
  XOR2_X1 Red_MCInst_MC2_v3_3Inst_0_U3  ( .A(MCInst_MC2_v3_2 [3]), .B(
        MCInst_MC2_v3_2 [2]), .Z(Red_MCInst_MC2_v3_3[0] ) );
  XNOR2_X1 Red_MCInst_MC2_r0Inst_XORInst_0_0_U3  ( .A(
        Red_MCInst_MC2_r0Inst_XORInst_0_0_n5 ), .B(
        Red_MCInst_MC2_r0Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback[13]) );
  XNOR2_X1 Red_MCInst_MC2_r0Inst_XORInst_0_0_U2  ( .A(
        Red_MCInst_MC2_v3_0[0] ), .B(Red_MCInst_MC2_v2_0[0] ), .ZN(
        Red_MCInst_MC2_r0Inst_XORInst_0_0_n4 ) );
  XOR2_X1 Red_MCInst_MC2_r0Inst_XORInst_0_0_U1  ( .A(Red_MCInst_MC2_v0_0[0] ), .B(Red_MCInst_MC2_v1_0[0] ), .Z(Red_MCInst_MC2_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 Red_MCInst_MC2_r1Inst_XORInst_0_0_U3  ( .A(
        Red_MCInst_MC2_r1Inst_XORInst_0_0_n5 ), .B(
        Red_MCInst_MC2_r1Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback[9]) );
  XNOR2_X1 Red_MCInst_MC2_r1Inst_XORInst_0_0_U2  ( .A(
        Red_MCInst_MC2_v3_1[0] ), .B(Red_MCInst_MC2_v2_1[0] ), .ZN(
        Red_MCInst_MC2_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 Red_MCInst_MC2_r1Inst_XORInst_0_0_U1  ( .A(Red_MCInst_MC2_v0_1[0] ), .B(Red_MCInst_MC2_v1_1[0] ), .Z(Red_MCInst_MC2_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 Red_MCInst_MC2_r2Inst_XORInst_0_0_U3  ( .A(
        Red_MCInst_MC2_r2Inst_XORInst_0_0_n5 ), .B(
        Red_MCInst_MC2_r2Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback[5]) );
  XNOR2_X1 Red_MCInst_MC2_r2Inst_XORInst_0_0_U2  ( .A(
        Red_MCInst_MC2_v3_2[0] ), .B(Red_MCInst_MC2_v2_2[0] ), .ZN(
        Red_MCInst_MC2_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 Red_MCInst_MC2_r2Inst_XORInst_0_0_U1  ( .A(Red_MCInst_MC2_v0_2[0] ), .B(Red_MCInst_MC2_v1_2[0] ), .Z(Red_MCInst_MC2_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 Red_MCInst_MC2_r3Inst_XORInst_0_0_U3  ( .A(
        Red_MCInst_MC2_r3Inst_XORInst_0_0_n5 ), .B(
        Red_MCInst_MC2_r3Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback[1]) );
  XNOR2_X1 Red_MCInst_MC2_r3Inst_XORInst_0_0_U2  ( .A(
        Red_MCInst_MC2_v3_3[0] ), .B(Red_MCInst_MC2_v2_3[0] ), .ZN(
        Red_MCInst_MC2_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 Red_MCInst_MC2_r3Inst_XORInst_0_0_U1  ( .A(Red_MCInst_MC2_v0_3[0] ), .B(Red_MCInst_MC2_v1_3[0] ), .Z(Red_MCInst_MC2_r3Inst_XORInst_0_0_n5 ) );
  XOR2_X1 Red_MCInst_MC3_v0_0Inst_0_U3  ( .A(Red_MCInst_MC3_v0_1[0] ), .B(
        MCInst_MC3_v0_0 [3]), .Z(Red_MCInst_MC3_v0_0[0] ) );
  XOR2_X1 Red_MCInst_MC3_v0_2Inst_0_U3  ( .A(Red_MCInst_MC3_v0_1[0] ), .B(
        MCInst_MC3_v0_3 [0]), .Z(Red_MCInst_MC3_v0_2[0] ) );
  XNOR2_X1 Red_MCInst_MC3_v0_3Inst_0_U4  ( .A(Red_MCInst_MC3_v0_3Inst_0_n2 ), 
        .B(MCInst_MC3_v0_0 [3]), .ZN(Red_MCInst_MC3_v0_3[0] ) );
  XNOR2_X1 Red_MCInst_MC3_v0_3Inst_0_U3  ( .A(MCInst_MC3_v0_3 [3]), .B(
        Red_MCInst_MC3_v0_1[0] ), .ZN(Red_MCInst_MC3_v0_3Inst_0_n2 ) );
  XNOR2_X1 Red_MCInst_MC3_v1_0Inst_0_U5  ( .A(Red_MCInst_MC3_v1_0Inst_0_n4 ), 
        .B(Red_MCInst_MC3_v1_0Inst_0_n3 ), .ZN(Red_MCInst_MC3_v1_0[0] ) );
  XNOR2_X1 Red_MCInst_MC3_v1_0Inst_0_U4  ( .A(MCInst_MC3_v1_3 [2]), .B(
        MCInst_MC3_v1_0 [0]), .ZN(Red_MCInst_MC3_v1_0Inst_0_n3 ) );
  XOR2_X1 Red_MCInst_MC3_v1_0Inst_0_U3  ( .A(Red_MCInst_MC3_v1_1[0] ), .B(
        MCInst_MC3_v1_0 [3]), .Z(Red_MCInst_MC3_v1_0Inst_0_n4 ) );
  XOR2_X1 Red_MCInst_MC3_v1_2Inst_0_U3  ( .A(MCInst_MC3_v1_0 [0]), .B(
        Red_MCInst_MC3_v1_1[0] ), .Z(Red_MCInst_MC3_v1_2[0] ) );
  XNOR2_X1 Red_MCInst_MC3_v1_3Inst_0_U4  ( .A(Red_MCInst_MC3_v1_3Inst_0_n2 ), 
        .B(MCInst_MC3_v1_3 [2]), .ZN(Red_MCInst_MC3_v1_3[0] ) );
  XNOR2_X1 Red_MCInst_MC3_v1_3Inst_0_U3  ( .A(Red_MCInst_MC3_v1_1[0] ), .B(
        MCInst_MC3_v1_0 [0]), .ZN(Red_MCInst_MC3_v1_3Inst_0_n2 ) );
  XNOR2_X1 Red_MCInst_MC3_v2_0Inst_0_U4  ( .A(Red_MCInst_MC3_v2_0Inst_0_n2 ), 
        .B(MCInst_MC3_v2_0 [2]), .ZN(Red_MCInst_MC3_v2_0[0] ) );
  XNOR2_X1 Red_MCInst_MC3_v2_0Inst_0_U3  ( .A(MCInst_MC3_v2_0 [3]), .B(
        MCInst_MC3_v2_3 [1]), .ZN(Red_MCInst_MC3_v2_0Inst_0_n2 ) );
  XOR2_X1 Red_MCInst_MC3_v2_1Inst_0_U3  ( .A(MCInst_MC3_v2_0 [3]), .B(
        MCInst_MC3_v2_0 [0]), .Z(Red_MCInst_MC3_v2_1[0] ) );
  XOR2_X1 Red_MCInst_MC3_v2_2Inst_0_U3  ( .A(MCInst_MC3_v2_0 [2]), .B(
        MCInst_MC3_v2_0 [3]), .Z(Red_MCInst_MC3_v2_2[0] ) );
  XOR2_X1 Red_MCInst_MC3_v2_3Inst_0_U3  ( .A(MCInst_MC3_v2_0 [2]), .B(
        MCInst_MC3_v2_0 [0]), .Z(Red_MCInst_MC3_v2_3[0] ) );
  XNOR2_X1 Red_MCInst_MC3_v3_0Inst_0_U4  ( .A(Red_MCInst_MC3_v3_0Inst_0_n2 ), 
        .B(MCInst_MC3_v3_0 [2]), .ZN(Red_MCInst_MC3_v3_0[0] ) );
  XNOR2_X1 Red_MCInst_MC3_v3_0Inst_0_U3  ( .A(Red_MCInst_MC3_v3_1[0] ), .B(
        MCInst_MC3_v3_2 [3]), .ZN(Red_MCInst_MC3_v3_0Inst_0_n2 ) );
  XNOR2_X1 Red_MCInst_MC3_v3_2Inst_0_U4  ( .A(Red_MCInst_MC3_v3_2Inst_0_n2 ), 
        .B(Red_MCInst_MC3_v3_1[0] ), .ZN(Red_MCInst_MC3_v3_2[0] ) );
  XNOR2_X1 Red_MCInst_MC3_v3_2Inst_0_U3  ( .A(MCInst_MC3_v3_2 [2]), .B(
        MCInst_MC3_v3_0 [2]), .ZN(Red_MCInst_MC3_v3_2Inst_0_n2 ) );
  XOR2_X1 Red_MCInst_MC3_v3_3Inst_0_U3  ( .A(MCInst_MC3_v3_2 [3]), .B(
        MCInst_MC3_v3_2 [2]), .Z(Red_MCInst_MC3_v3_3[0] ) );
  XNOR2_X1 Red_MCInst_MC3_r0Inst_XORInst_0_0_U3  ( .A(
        Red_MCInst_MC3_r0Inst_XORInst_0_0_n5 ), .B(
        Red_MCInst_MC3_r0Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback[12]) );
  XNOR2_X1 Red_MCInst_MC3_r0Inst_XORInst_0_0_U2  ( .A(
        Red_MCInst_MC3_v3_0[0] ), .B(Red_MCInst_MC3_v2_0[0] ), .ZN(
        Red_MCInst_MC3_r0Inst_XORInst_0_0_n4 ) );
  XOR2_X1 Red_MCInst_MC3_r0Inst_XORInst_0_0_U1  ( .A(Red_MCInst_MC3_v0_0[0] ), .B(Red_MCInst_MC3_v1_0[0] ), .Z(Red_MCInst_MC3_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 Red_MCInst_MC3_r1Inst_XORInst_0_0_U3  ( .A(
        Red_MCInst_MC3_r1Inst_XORInst_0_0_n5 ), .B(
        Red_MCInst_MC3_r1Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback[8]) );
  XNOR2_X1 Red_MCInst_MC3_r1Inst_XORInst_0_0_U2  ( .A(
        Red_MCInst_MC3_v3_1[0] ), .B(Red_MCInst_MC3_v2_1[0] ), .ZN(
        Red_MCInst_MC3_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 Red_MCInst_MC3_r1Inst_XORInst_0_0_U1  ( .A(Red_MCInst_MC3_v0_1[0] ), .B(Red_MCInst_MC3_v1_1[0] ), .Z(Red_MCInst_MC3_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 Red_MCInst_MC3_r2Inst_XORInst_0_0_U3  ( .A(
        Red_MCInst_MC3_r2Inst_XORInst_0_0_n5 ), .B(
        Red_MCInst_MC3_r2Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback[4]) );
  XNOR2_X1 Red_MCInst_MC3_r2Inst_XORInst_0_0_U2  ( .A(
        Red_MCInst_MC3_v3_2[0] ), .B(Red_MCInst_MC3_v2_2[0] ), .ZN(
        Red_MCInst_MC3_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 Red_MCInst_MC3_r2Inst_XORInst_0_0_U1  ( .A(Red_MCInst_MC3_v0_2[0] ), .B(Red_MCInst_MC3_v1_2[0] ), .Z(Red_MCInst_MC3_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 Red_MCInst_MC3_r3Inst_XORInst_0_0_U3  ( .A(
        Red_MCInst_MC3_r3Inst_XORInst_0_0_n5 ), .B(
        Red_MCInst_MC3_r3Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback[0]) );
  XNOR2_X1 Red_MCInst_MC3_r3Inst_XORInst_0_0_U2  ( .A(
        Red_MCInst_MC3_v3_3[0] ), .B(Red_MCInst_MC3_v2_3[0] ), .ZN(
        Red_MCInst_MC3_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 Red_MCInst_MC3_r3Inst_XORInst_0_0_U1  ( .A(Red_MCInst_MC3_v0_3[0] ), .B(Red_MCInst_MC3_v1_3[0] ), .Z(Red_MCInst_MC3_r3Inst_XORInst_0_0_n5 ) );
  DFF_X1 RedStateReg_s_current_state_reg[0]  ( .D(Red_Feedback[0]), .CK(clk), 
        .Q(Red_SubCellInput[0]) );
  DFF_X1 RedStateReg_s_current_state_reg[1]  ( .D(Red_Feedback[1]), .CK(clk), 
        .Q(Red_SubCellInput[1]) );
  DFF_X1 RedStateReg_s_current_state_reg[2]  ( .D(Red_Feedback[2]), .CK(clk), 
        .Q(Red_SubCellInput[2]) );
  DFF_X1 RedStateReg_s_current_state_reg[3]  ( .D(Red_Feedback[3]), .CK(clk), 
        .Q(Red_SubCellInput[3]) );
  DFF_X1 RedStateReg_s_current_state_reg[4]  ( .D(Red_Feedback[4]), .CK(clk), 
        .Q(Red_SubCellInput[4]) );
  DFF_X1 RedStateReg_s_current_state_reg[5]  ( .D(Red_Feedback[5]), .CK(clk), 
        .Q(Red_SubCellInput[5]) );
  DFF_X1 RedStateReg_s_current_state_reg[6]  ( .D(Red_Feedback[6]), .CK(clk), 
        .Q(Red_SubCellInput[6]) );
  DFF_X1 RedStateReg_s_current_state_reg[7]  ( .D(Red_Feedback[7]), .CK(clk), 
        .Q(Red_SubCellInput[7]) );
  DFF_X1 RedStateReg_s_current_state_reg[8]  ( .D(Red_Feedback[8]), .CK(clk), 
        .Q(Red_SubCellInput[8]) );
  DFF_X1 RedStateReg_s_current_state_reg[9]  ( .D(Red_Feedback[9]), .CK(clk), 
        .Q(Red_SubCellInput[9]) );
  DFF_X1 RedStateReg_s_current_state_reg[10]  ( .D(Red_Feedback[10]), .CK(clk), .Q(Red_SubCellInput[10]) );
  DFF_X1 RedStateReg_s_current_state_reg[11]  ( .D(Red_Feedback[11]), .CK(clk), .Q(Red_SubCellInput[11]) );
  DFF_X1 RedStateReg_s_current_state_reg[12]  ( .D(Red_Feedback[12]), .CK(clk), .Q(Red_SubCellInput[12]) );
  DFF_X1 RedStateReg_s_current_state_reg[13]  ( .D(Red_Feedback[13]), .CK(clk), .Q(Red_SubCellInput[13]) );
  DFF_X1 RedStateReg_s_current_state_reg[14]  ( .D(Red_Feedback[14]), .CK(clk), .Q(Red_SubCellInput[14]) );
  DFF_X1 RedStateReg_s_current_state_reg[15]  ( .D(Red_Feedback[15]), .CK(clk), .Q(Red_SubCellInput[15]) );
  NAND2_X1 Red_SubCellInst2_LFInst_0_LFInst_0_U6  ( .A1(
        Red_SubCellInst2_LFInst_0_LFInst_0_n6 ), .A2(
        Red_SubCellInst2_LFInst_0_LFInst_0_n5 ), .ZN(Red_ShiftRowsOutput2[3])
         );
  NAND2_X1 Red_SubCellInst2_LFInst_0_LFInst_0_U5  ( .A1(SubCellInput[3]), 
        .A2(SubCellInput[2]), .ZN(Red_SubCellInst2_LFInst_0_LFInst_0_n5 ) );
  NAND2_X1 Red_SubCellInst2_LFInst_0_LFInst_0_U4  ( .A1(SubCellInput[0]), 
        .A2(Red_SubCellInst2_LFInst_0_LFInst_0_n4 ), .ZN(
        Red_SubCellInst2_LFInst_0_LFInst_0_n6 ) );
  OR2_X1 Red_SubCellInst2_LFInst_0_LFInst_0_U3  ( .A1(SubCellInput[1]), .A2(
        SubCellInput[3]), .ZN(Red_SubCellInst2_LFInst_0_LFInst_0_n4 ) );
  NAND2_X1 Red_SubCellInst2_LFInst_1_LFInst_0_U6  ( .A1(
        Red_SubCellInst2_LFInst_1_LFInst_0_n6 ), .A2(
        Red_SubCellInst2_LFInst_1_LFInst_0_n5 ), .ZN(Red_ShiftRowsOutput2[0])
         );
  NAND2_X1 Red_SubCellInst2_LFInst_1_LFInst_0_U5  ( .A1(SubCellInput[7]), 
        .A2(SubCellInput[6]), .ZN(Red_SubCellInst2_LFInst_1_LFInst_0_n5 ) );
  NAND2_X1 Red_SubCellInst2_LFInst_1_LFInst_0_U4  ( .A1(SubCellInput[4]), 
        .A2(Red_SubCellInst2_LFInst_1_LFInst_0_n4 ), .ZN(
        Red_SubCellInst2_LFInst_1_LFInst_0_n6 ) );
  OR2_X1 Red_SubCellInst2_LFInst_1_LFInst_0_U3  ( .A1(SubCellInput[5]), .A2(
        SubCellInput[7]), .ZN(Red_SubCellInst2_LFInst_1_LFInst_0_n4 ) );
  NAND2_X1 Red_SubCellInst2_LFInst_2_LFInst_0_U6  ( .A1(
        Red_SubCellInst2_LFInst_2_LFInst_0_n6 ), .A2(
        Red_SubCellInst2_LFInst_2_LFInst_0_n5 ), .ZN(Red_ShiftRowsOutput2[1])
         );
  NAND2_X1 Red_SubCellInst2_LFInst_2_LFInst_0_U5  ( .A1(SubCellInput[11]), 
        .A2(SubCellInput[10]), .ZN(Red_SubCellInst2_LFInst_2_LFInst_0_n5 ) );
  NAND2_X1 Red_SubCellInst2_LFInst_2_LFInst_0_U4  ( .A1(SubCellInput[8]), 
        .A2(Red_SubCellInst2_LFInst_2_LFInst_0_n4 ), .ZN(
        Red_SubCellInst2_LFInst_2_LFInst_0_n6 ) );
  OR2_X1 Red_SubCellInst2_LFInst_2_LFInst_0_U3  ( .A1(SubCellInput[9]), .A2(
        SubCellInput[11]), .ZN(Red_SubCellInst2_LFInst_2_LFInst_0_n4 ) );
  NAND2_X1 Red_SubCellInst2_LFInst_3_LFInst_0_U6  ( .A1(
        Red_SubCellInst2_LFInst_3_LFInst_0_n6 ), .A2(
        Red_SubCellInst2_LFInst_3_LFInst_0_n5 ), .ZN(Red_ShiftRowsOutput2[2])
         );
  NAND2_X1 Red_SubCellInst2_LFInst_3_LFInst_0_U5  ( .A1(SubCellInput[15]), 
        .A2(SubCellInput[14]), .ZN(Red_SubCellInst2_LFInst_3_LFInst_0_n5 ) );
  NAND2_X1 Red_SubCellInst2_LFInst_3_LFInst_0_U4  ( .A1(SubCellInput[12]), 
        .A2(Red_SubCellInst2_LFInst_3_LFInst_0_n4 ), .ZN(
        Red_SubCellInst2_LFInst_3_LFInst_0_n6 ) );
  OR2_X1 Red_SubCellInst2_LFInst_3_LFInst_0_U3  ( .A1(SubCellInput[13]), .A2(
        SubCellInput[15]), .ZN(Red_SubCellInst2_LFInst_3_LFInst_0_n4 ) );
  NAND2_X1 Red_SubCellInst2_LFInst_4_LFInst_0_U6  ( .A1(
        Red_SubCellInst2_LFInst_4_LFInst_0_n6 ), .A2(
        Red_SubCellInst2_LFInst_4_LFInst_0_n5 ), .ZN(Red_ShiftRowsOutput2[6])
         );
  NAND2_X1 Red_SubCellInst2_LFInst_4_LFInst_0_U5  ( .A1(SubCellInput[19]), 
        .A2(SubCellInput[18]), .ZN(Red_SubCellInst2_LFInst_4_LFInst_0_n5 ) );
  NAND2_X1 Red_SubCellInst2_LFInst_4_LFInst_0_U4  ( .A1(SubCellInput[16]), 
        .A2(Red_SubCellInst2_LFInst_4_LFInst_0_n4 ), .ZN(
        Red_SubCellInst2_LFInst_4_LFInst_0_n6 ) );
  OR2_X1 Red_SubCellInst2_LFInst_4_LFInst_0_U3  ( .A1(SubCellInput[17]), .A2(
        SubCellInput[19]), .ZN(Red_SubCellInst2_LFInst_4_LFInst_0_n4 ) );
  NAND2_X1 Red_SubCellInst2_LFInst_5_LFInst_0_U6  ( .A1(
        Red_SubCellInst2_LFInst_5_LFInst_0_n6 ), .A2(
        Red_SubCellInst2_LFInst_5_LFInst_0_n5 ), .ZN(Red_ShiftRowsOutput2[7])
         );
  NAND2_X1 Red_SubCellInst2_LFInst_5_LFInst_0_U5  ( .A1(SubCellInput[23]), 
        .A2(SubCellInput[22]), .ZN(Red_SubCellInst2_LFInst_5_LFInst_0_n5 ) );
  NAND2_X1 Red_SubCellInst2_LFInst_5_LFInst_0_U4  ( .A1(SubCellInput[20]), 
        .A2(Red_SubCellInst2_LFInst_5_LFInst_0_n4 ), .ZN(
        Red_SubCellInst2_LFInst_5_LFInst_0_n6 ) );
  OR2_X1 Red_SubCellInst2_LFInst_5_LFInst_0_U3  ( .A1(SubCellInput[21]), .A2(
        SubCellInput[23]), .ZN(Red_SubCellInst2_LFInst_5_LFInst_0_n4 ) );
  NAND2_X1 Red_SubCellInst2_LFInst_6_LFInst_0_U6  ( .A1(
        Red_SubCellInst2_LFInst_6_LFInst_0_n6 ), .A2(
        Red_SubCellInst2_LFInst_6_LFInst_0_n5 ), .ZN(Red_ShiftRowsOutput2[4])
         );
  NAND2_X1 Red_SubCellInst2_LFInst_6_LFInst_0_U5  ( .A1(SubCellInput[27]), 
        .A2(SubCellInput[26]), .ZN(Red_SubCellInst2_LFInst_6_LFInst_0_n5 ) );
  NAND2_X1 Red_SubCellInst2_LFInst_6_LFInst_0_U4  ( .A1(SubCellInput[24]), 
        .A2(Red_SubCellInst2_LFInst_6_LFInst_0_n4 ), .ZN(
        Red_SubCellInst2_LFInst_6_LFInst_0_n6 ) );
  OR2_X1 Red_SubCellInst2_LFInst_6_LFInst_0_U3  ( .A1(SubCellInput[25]), .A2(
        SubCellInput[27]), .ZN(Red_SubCellInst2_LFInst_6_LFInst_0_n4 ) );
  NAND2_X1 Red_SubCellInst2_LFInst_7_LFInst_0_U6  ( .A1(
        Red_SubCellInst2_LFInst_7_LFInst_0_n6 ), .A2(
        Red_SubCellInst2_LFInst_7_LFInst_0_n5 ), .ZN(Red_ShiftRowsOutput2[5])
         );
  NAND2_X1 Red_SubCellInst2_LFInst_7_LFInst_0_U5  ( .A1(SubCellInput[31]), 
        .A2(SubCellInput[30]), .ZN(Red_SubCellInst2_LFInst_7_LFInst_0_n5 ) );
  NAND2_X1 Red_SubCellInst2_LFInst_7_LFInst_0_U4  ( .A1(SubCellInput[28]), 
        .A2(Red_SubCellInst2_LFInst_7_LFInst_0_n4 ), .ZN(
        Red_SubCellInst2_LFInst_7_LFInst_0_n6 ) );
  OR2_X1 Red_SubCellInst2_LFInst_7_LFInst_0_U3  ( .A1(SubCellInput[29]), .A2(
        SubCellInput[31]), .ZN(Red_SubCellInst2_LFInst_7_LFInst_0_n4 ) );
  NAND2_X1 Red_SubCellInst2_LFInst_8_LFInst_0_U6  ( .A1(
        Red_SubCellInst2_LFInst_8_LFInst_0_n6 ), .A2(
        Red_SubCellInst2_LFInst_8_LFInst_0_n5 ), .ZN(Red_ShiftRowsOutput2[9])
         );
  NAND2_X1 Red_SubCellInst2_LFInst_8_LFInst_0_U5  ( .A1(SubCellInput[35]), 
        .A2(SubCellInput[34]), .ZN(Red_SubCellInst2_LFInst_8_LFInst_0_n5 ) );
  NAND2_X1 Red_SubCellInst2_LFInst_8_LFInst_0_U4  ( .A1(SubCellInput[32]), 
        .A2(Red_SubCellInst2_LFInst_8_LFInst_0_n4 ), .ZN(
        Red_SubCellInst2_LFInst_8_LFInst_0_n6 ) );
  OR2_X1 Red_SubCellInst2_LFInst_8_LFInst_0_U3  ( .A1(SubCellInput[33]), .A2(
        SubCellInput[35]), .ZN(Red_SubCellInst2_LFInst_8_LFInst_0_n4 ) );
  NAND2_X1 Red_SubCellInst2_LFInst_9_LFInst_0_U6  ( .A1(
        Red_SubCellInst2_LFInst_9_LFInst_0_n6 ), .A2(
        Red_SubCellInst2_LFInst_9_LFInst_0_n5 ), .ZN(Red_ShiftRowsOutput2[10]) );
  NAND2_X1 Red_SubCellInst2_LFInst_9_LFInst_0_U5  ( .A1(SubCellInput[39]), 
        .A2(SubCellInput[38]), .ZN(Red_SubCellInst2_LFInst_9_LFInst_0_n5 ) );
  NAND2_X1 Red_SubCellInst2_LFInst_9_LFInst_0_U4  ( .A1(SubCellInput[36]), 
        .A2(Red_SubCellInst2_LFInst_9_LFInst_0_n4 ), .ZN(
        Red_SubCellInst2_LFInst_9_LFInst_0_n6 ) );
  OR2_X1 Red_SubCellInst2_LFInst_9_LFInst_0_U3  ( .A1(SubCellInput[37]), .A2(
        SubCellInput[39]), .ZN(Red_SubCellInst2_LFInst_9_LFInst_0_n4 ) );
  NAND2_X1 Red_SubCellInst2_LFInst_10_LFInst_0_U6  ( .A1(
        Red_SubCellInst2_LFInst_10_LFInst_0_n6 ), .A2(
        Red_SubCellInst2_LFInst_10_LFInst_0_n5 ), .ZN(
        Red_ShiftRowsOutput2[11]) );
  NAND2_X1 Red_SubCellInst2_LFInst_10_LFInst_0_U5  ( .A1(SubCellInput[43]), 
        .A2(SubCellInput[42]), .ZN(Red_SubCellInst2_LFInst_10_LFInst_0_n5 )
         );
  NAND2_X1 Red_SubCellInst2_LFInst_10_LFInst_0_U4  ( .A1(SubCellInput[40]), 
        .A2(Red_SubCellInst2_LFInst_10_LFInst_0_n4 ), .ZN(
        Red_SubCellInst2_LFInst_10_LFInst_0_n6 ) );
  OR2_X1 Red_SubCellInst2_LFInst_10_LFInst_0_U3  ( .A1(SubCellInput[41]), 
        .A2(SubCellInput[43]), .ZN(Red_SubCellInst2_LFInst_10_LFInst_0_n4 )
         );
  NAND2_X1 Red_SubCellInst2_LFInst_11_LFInst_0_U6  ( .A1(
        Red_SubCellInst2_LFInst_11_LFInst_0_n6 ), .A2(
        Red_SubCellInst2_LFInst_11_LFInst_0_n5 ), .ZN(Red_ShiftRowsOutput2[8]) );
  NAND2_X1 Red_SubCellInst2_LFInst_11_LFInst_0_U5  ( .A1(SubCellInput[47]), 
        .A2(SubCellInput[46]), .ZN(Red_SubCellInst2_LFInst_11_LFInst_0_n5 )
         );
  NAND2_X1 Red_SubCellInst2_LFInst_11_LFInst_0_U4  ( .A1(SubCellInput[44]), 
        .A2(Red_SubCellInst2_LFInst_11_LFInst_0_n4 ), .ZN(
        Red_SubCellInst2_LFInst_11_LFInst_0_n6 ) );
  OR2_X1 Red_SubCellInst2_LFInst_11_LFInst_0_U3  ( .A1(SubCellInput[45]), 
        .A2(SubCellInput[47]), .ZN(Red_SubCellInst2_LFInst_11_LFInst_0_n4 )
         );
  NAND2_X1 Red_SubCellInst2_LFInst_12_LFInst_0_U6  ( .A1(
        Red_SubCellInst2_LFInst_12_LFInst_0_n6 ), .A2(
        Red_SubCellInst2_LFInst_12_LFInst_0_n5 ), .ZN(
        Red_ShiftRowsOutput2[12]) );
  NAND2_X1 Red_SubCellInst2_LFInst_12_LFInst_0_U5  ( .A1(SubCellInput[51]), 
        .A2(SubCellInput[50]), .ZN(Red_SubCellInst2_LFInst_12_LFInst_0_n5 )
         );
  NAND2_X1 Red_SubCellInst2_LFInst_12_LFInst_0_U4  ( .A1(SubCellInput[48]), 
        .A2(Red_SubCellInst2_LFInst_12_LFInst_0_n4 ), .ZN(
        Red_SubCellInst2_LFInst_12_LFInst_0_n6 ) );
  OR2_X1 Red_SubCellInst2_LFInst_12_LFInst_0_U3  ( .A1(SubCellInput[49]), 
        .A2(SubCellInput[51]), .ZN(Red_SubCellInst2_LFInst_12_LFInst_0_n4 )
         );
  NAND2_X1 Red_SubCellInst2_LFInst_13_LFInst_0_U6  ( .A1(
        Red_SubCellInst2_LFInst_13_LFInst_0_n6 ), .A2(
        Red_SubCellInst2_LFInst_13_LFInst_0_n5 ), .ZN(
        Red_ShiftRowsOutput2[13]) );
  NAND2_X1 Red_SubCellInst2_LFInst_13_LFInst_0_U5  ( .A1(SubCellInput[55]), 
        .A2(SubCellInput[54]), .ZN(Red_SubCellInst2_LFInst_13_LFInst_0_n5 )
         );
  NAND2_X1 Red_SubCellInst2_LFInst_13_LFInst_0_U4  ( .A1(SubCellInput[52]), 
        .A2(Red_SubCellInst2_LFInst_13_LFInst_0_n4 ), .ZN(
        Red_SubCellInst2_LFInst_13_LFInst_0_n6 ) );
  OR2_X1 Red_SubCellInst2_LFInst_13_LFInst_0_U3  ( .A1(SubCellInput[53]), 
        .A2(SubCellInput[55]), .ZN(Red_SubCellInst2_LFInst_13_LFInst_0_n4 )
         );
  NAND2_X1 Red_SubCellInst2_LFInst_14_LFInst_0_U6  ( .A1(
        Red_SubCellInst2_LFInst_14_LFInst_0_n6 ), .A2(
        Red_SubCellInst2_LFInst_14_LFInst_0_n5 ), .ZN(
        Red_ShiftRowsOutput2[14]) );
  NAND2_X1 Red_SubCellInst2_LFInst_14_LFInst_0_U5  ( .A1(SubCellInput[59]), 
        .A2(SubCellInput[58]), .ZN(Red_SubCellInst2_LFInst_14_LFInst_0_n5 )
         );
  NAND2_X1 Red_SubCellInst2_LFInst_14_LFInst_0_U4  ( .A1(SubCellInput[56]), 
        .A2(Red_SubCellInst2_LFInst_14_LFInst_0_n4 ), .ZN(
        Red_SubCellInst2_LFInst_14_LFInst_0_n6 ) );
  OR2_X1 Red_SubCellInst2_LFInst_14_LFInst_0_U3  ( .A1(SubCellInput[57]), 
        .A2(SubCellInput[59]), .ZN(Red_SubCellInst2_LFInst_14_LFInst_0_n4 )
         );
  NAND2_X1 Red_SubCellInst2_LFInst_15_LFInst_0_U6  ( .A1(
        Red_SubCellInst2_LFInst_15_LFInst_0_n6 ), .A2(
        Red_SubCellInst2_LFInst_15_LFInst_0_n5 ), .ZN(
        Red_ShiftRowsOutput2[15]) );
  NAND2_X1 Red_SubCellInst2_LFInst_15_LFInst_0_U5  ( .A1(SubCellInput[63]), 
        .A2(SubCellInput[62]), .ZN(Red_SubCellInst2_LFInst_15_LFInst_0_n5 )
         );
  NAND2_X1 Red_SubCellInst2_LFInst_15_LFInst_0_U4  ( .A1(SubCellInput[60]), 
        .A2(Red_SubCellInst2_LFInst_15_LFInst_0_n4 ), .ZN(
        Red_SubCellInst2_LFInst_15_LFInst_0_n6 ) );
  OR2_X1 Red_SubCellInst2_LFInst_15_LFInst_0_U3  ( .A1(SubCellInput[61]), 
        .A2(SubCellInput[63]), .ZN(Red_SubCellInst2_LFInst_15_LFInst_0_n4 )
         );
  XOR2_X1 Red_MCInst2_MC0_v0_0Inst_0_U3  ( .A(Red_MCInst2_MC0_v0_1[0] ), .B(
        MCInst2_MC0_v0_0 [3]), .Z(Red_MCInst2_MC0_v0_0[0] ) );
  XOR2_X1 Red_MCInst2_MC0_v0_2Inst_0_U3  ( .A(Red_MCInst2_MC0_v0_1[0] ), .B(
        MCInst2_MC0_v0_3 [0]), .Z(Red_MCInst2_MC0_v0_2[0] ) );
  XNOR2_X1 Red_MCInst2_MC0_v0_3Inst_0_U4  ( .A(
        Red_MCInst2_MC0_v0_3Inst_0_n2 ), .B(MCInst2_MC0_v0_0 [3]), .ZN(
        Red_MCInst2_MC0_v0_3[0] ) );
  XNOR2_X1 Red_MCInst2_MC0_v0_3Inst_0_U3  ( .A(MCInst2_MC0_v0_3 [3]), .B(
        Red_MCInst2_MC0_v0_1[0] ), .ZN(Red_MCInst2_MC0_v0_3Inst_0_n2 ) );
  XNOR2_X1 Red_MCInst2_MC0_v1_0Inst_0_U5  ( .A(
        Red_MCInst2_MC0_v1_0Inst_0_n4 ), .B(Red_MCInst2_MC0_v1_0Inst_0_n3 ), 
        .ZN(Red_MCInst2_MC0_v1_0[0] ) );
  XNOR2_X1 Red_MCInst2_MC0_v1_0Inst_0_U4  ( .A(MCInst2_MC0_v1_3 [2]), .B(
        MCInst2_MC0_v1_0 [0]), .ZN(Red_MCInst2_MC0_v1_0Inst_0_n3 ) );
  XOR2_X1 Red_MCInst2_MC0_v1_0Inst_0_U3  ( .A(Red_MCInst2_MC0_v1_1[0] ), .B(
        MCInst2_MC0_v1_0 [3]), .Z(Red_MCInst2_MC0_v1_0Inst_0_n4 ) );
  XOR2_X1 Red_MCInst2_MC0_v1_2Inst_0_U3  ( .A(MCInst2_MC0_v1_0 [0]), .B(
        Red_MCInst2_MC0_v1_1[0] ), .Z(Red_MCInst2_MC0_v1_2[0] ) );
  XNOR2_X1 Red_MCInst2_MC0_v1_3Inst_0_U4  ( .A(
        Red_MCInst2_MC0_v1_3Inst_0_n2 ), .B(MCInst2_MC0_v1_3 [2]), .ZN(
        Red_MCInst2_MC0_v1_3[0] ) );
  XNOR2_X1 Red_MCInst2_MC0_v1_3Inst_0_U3  ( .A(Red_MCInst2_MC0_v1_1[0] ), 
        .B(MCInst2_MC0_v1_0 [0]), .ZN(Red_MCInst2_MC0_v1_3Inst_0_n2 ) );
  XNOR2_X1 Red_MCInst2_MC0_v2_0Inst_0_U4  ( .A(
        Red_MCInst2_MC0_v2_0Inst_0_n2 ), .B(MCInst2_MC0_v2_0 [2]), .ZN(
        Red_MCInst2_MC0_v2_0[0] ) );
  XNOR2_X1 Red_MCInst2_MC0_v2_0Inst_0_U3  ( .A(MCInst2_MC0_v2_0 [3]), .B(
        MCInst2_MC0_v2_3 [1]), .ZN(Red_MCInst2_MC0_v2_0Inst_0_n2 ) );
  XOR2_X1 Red_MCInst2_MC0_v2_1Inst_0_U3  ( .A(MCInst2_MC0_v2_0 [3]), .B(
        MCInst2_MC0_v2_0 [0]), .Z(Red_MCInst2_MC0_v2_1[0] ) );
  XOR2_X1 Red_MCInst2_MC0_v2_2Inst_0_U3  ( .A(MCInst2_MC0_v2_0 [2]), .B(
        MCInst2_MC0_v2_0 [3]), .Z(Red_MCInst2_MC0_v2_2[0] ) );
  XOR2_X1 Red_MCInst2_MC0_v2_3Inst_0_U3  ( .A(MCInst2_MC0_v2_0 [2]), .B(
        MCInst2_MC0_v2_0 [0]), .Z(Red_MCInst2_MC0_v2_3[0] ) );
  XNOR2_X1 Red_MCInst2_MC0_v3_0Inst_0_U4  ( .A(
        Red_MCInst2_MC0_v3_0Inst_0_n2 ), .B(MCInst2_MC0_v3_0 [2]), .ZN(
        Red_MCInst2_MC0_v3_0[0] ) );
  XNOR2_X1 Red_MCInst2_MC0_v3_0Inst_0_U3  ( .A(Red_MCInst2_MC0_v3_1[0] ), 
        .B(MCInst2_MC0_v3_2 [3]), .ZN(Red_MCInst2_MC0_v3_0Inst_0_n2 ) );
  XNOR2_X1 Red_MCInst2_MC0_v3_2Inst_0_U4  ( .A(
        Red_MCInst2_MC0_v3_2Inst_0_n2 ), .B(Red_MCInst2_MC0_v3_1[0] ), .ZN(
        Red_MCInst2_MC0_v3_2[0] ) );
  XNOR2_X1 Red_MCInst2_MC0_v3_2Inst_0_U3  ( .A(MCInst2_MC0_v3_2 [2]), .B(
        MCInst2_MC0_v3_0 [2]), .ZN(Red_MCInst2_MC0_v3_2Inst_0_n2 ) );
  XOR2_X1 Red_MCInst2_MC0_v3_3Inst_0_U3  ( .A(MCInst2_MC0_v3_2 [3]), .B(
        MCInst2_MC0_v3_2 [2]), .Z(Red_MCInst2_MC0_v3_3[0] ) );
  XNOR2_X1 Red_MCInst2_MC0_r0Inst_XORInst_0_0_U3  ( .A(
        Red_MCInst2_MC0_r0Inst_XORInst_0_0_n5 ), .B(
        Red_MCInst2_MC0_r0Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback2[15]) );
  XNOR2_X1 Red_MCInst2_MC0_r0Inst_XORInst_0_0_U2  ( .A(
        Red_MCInst2_MC0_v3_0[0] ), .B(Red_MCInst2_MC0_v2_0[0] ), .ZN(
        Red_MCInst2_MC0_r0Inst_XORInst_0_0_n4 ) );
  XOR2_X1 Red_MCInst2_MC0_r0Inst_XORInst_0_0_U1  ( .A(
        Red_MCInst2_MC0_v0_0[0] ), .B(Red_MCInst2_MC0_v1_0[0] ), .Z(
        Red_MCInst2_MC0_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 Red_MCInst2_MC0_r1Inst_XORInst_0_0_U3  ( .A(
        Red_MCInst2_MC0_r1Inst_XORInst_0_0_n5 ), .B(
        Red_MCInst2_MC0_r1Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback2[11]) );
  XNOR2_X1 Red_MCInst2_MC0_r1Inst_XORInst_0_0_U2  ( .A(
        Red_MCInst2_MC0_v3_1[0] ), .B(Red_MCInst2_MC0_v2_1[0] ), .ZN(
        Red_MCInst2_MC0_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 Red_MCInst2_MC0_r1Inst_XORInst_0_0_U1  ( .A(
        Red_MCInst2_MC0_v0_1[0] ), .B(Red_MCInst2_MC0_v1_1[0] ), .Z(
        Red_MCInst2_MC0_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 Red_MCInst2_MC0_r2Inst_XORInst_0_0_U3  ( .A(
        Red_MCInst2_MC0_r2Inst_XORInst_0_0_n5 ), .B(
        Red_MCInst2_MC0_r2Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback2[7]) );
  XNOR2_X1 Red_MCInst2_MC0_r2Inst_XORInst_0_0_U2  ( .A(
        Red_MCInst2_MC0_v3_2[0] ), .B(Red_MCInst2_MC0_v2_2[0] ), .ZN(
        Red_MCInst2_MC0_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 Red_MCInst2_MC0_r2Inst_XORInst_0_0_U1  ( .A(
        Red_MCInst2_MC0_v0_2[0] ), .B(Red_MCInst2_MC0_v1_2[0] ), .Z(
        Red_MCInst2_MC0_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 Red_MCInst2_MC0_r3Inst_XORInst_0_0_U3  ( .A(
        Red_MCInst2_MC0_r3Inst_XORInst_0_0_n5 ), .B(
        Red_MCInst2_MC0_r3Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback2[3]) );
  XNOR2_X1 Red_MCInst2_MC0_r3Inst_XORInst_0_0_U2  ( .A(
        Red_MCInst2_MC0_v3_3[0] ), .B(Red_MCInst2_MC0_v2_3[0] ), .ZN(
        Red_MCInst2_MC0_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 Red_MCInst2_MC0_r3Inst_XORInst_0_0_U1  ( .A(
        Red_MCInst2_MC0_v0_3[0] ), .B(Red_MCInst2_MC0_v1_3[0] ), .Z(
        Red_MCInst2_MC0_r3Inst_XORInst_0_0_n5 ) );
  XOR2_X1 Red_MCInst2_MC1_v0_0Inst_0_U3  ( .A(Red_MCInst2_MC1_v0_1[0] ), .B(
        MCInst2_MC1_v0_0 [3]), .Z(Red_MCInst2_MC1_v0_0[0] ) );
  XOR2_X1 Red_MCInst2_MC1_v0_2Inst_0_U3  ( .A(Red_MCInst2_MC1_v0_1[0] ), .B(
        MCInst2_MC1_v0_3 [0]), .Z(Red_MCInst2_MC1_v0_2[0] ) );
  XNOR2_X1 Red_MCInst2_MC1_v0_3Inst_0_U4  ( .A(
        Red_MCInst2_MC1_v0_3Inst_0_n2 ), .B(MCInst2_MC1_v0_0 [3]), .ZN(
        Red_MCInst2_MC1_v0_3[0] ) );
  XNOR2_X1 Red_MCInst2_MC1_v0_3Inst_0_U3  ( .A(MCInst2_MC1_v0_3 [3]), .B(
        Red_MCInst2_MC1_v0_1[0] ), .ZN(Red_MCInst2_MC1_v0_3Inst_0_n2 ) );
  XNOR2_X1 Red_MCInst2_MC1_v1_0Inst_0_U5  ( .A(
        Red_MCInst2_MC1_v1_0Inst_0_n4 ), .B(Red_MCInst2_MC1_v1_0Inst_0_n3 ), 
        .ZN(Red_MCInst2_MC1_v1_0[0] ) );
  XNOR2_X1 Red_MCInst2_MC1_v1_0Inst_0_U4  ( .A(MCInst2_MC1_v1_3 [2]), .B(
        MCInst2_MC1_v1_0 [0]), .ZN(Red_MCInst2_MC1_v1_0Inst_0_n3 ) );
  XOR2_X1 Red_MCInst2_MC1_v1_0Inst_0_U3  ( .A(Red_MCInst2_MC1_v1_1[0] ), .B(
        MCInst2_MC1_v1_0 [3]), .Z(Red_MCInst2_MC1_v1_0Inst_0_n4 ) );
  XOR2_X1 Red_MCInst2_MC1_v1_2Inst_0_U3  ( .A(MCInst2_MC1_v1_0 [0]), .B(
        Red_MCInst2_MC1_v1_1[0] ), .Z(Red_MCInst2_MC1_v1_2[0] ) );
  XNOR2_X1 Red_MCInst2_MC1_v1_3Inst_0_U4  ( .A(
        Red_MCInst2_MC1_v1_3Inst_0_n2 ), .B(MCInst2_MC1_v1_3 [2]), .ZN(
        Red_MCInst2_MC1_v1_3[0] ) );
  XNOR2_X1 Red_MCInst2_MC1_v1_3Inst_0_U3  ( .A(Red_MCInst2_MC1_v1_1[0] ), 
        .B(MCInst2_MC1_v1_0 [0]), .ZN(Red_MCInst2_MC1_v1_3Inst_0_n2 ) );
  XNOR2_X1 Red_MCInst2_MC1_v2_0Inst_0_U4  ( .A(
        Red_MCInst2_MC1_v2_0Inst_0_n2 ), .B(MCInst2_MC1_v2_0 [2]), .ZN(
        Red_MCInst2_MC1_v2_0[0] ) );
  XNOR2_X1 Red_MCInst2_MC1_v2_0Inst_0_U3  ( .A(MCInst2_MC1_v2_0 [3]), .B(
        MCInst2_MC1_v2_3 [1]), .ZN(Red_MCInst2_MC1_v2_0Inst_0_n2 ) );
  XOR2_X1 Red_MCInst2_MC1_v2_1Inst_0_U3  ( .A(MCInst2_MC1_v2_0 [3]), .B(
        MCInst2_MC1_v2_0 [0]), .Z(Red_MCInst2_MC1_v2_1[0] ) );
  XOR2_X1 Red_MCInst2_MC1_v2_2Inst_0_U3  ( .A(MCInst2_MC1_v2_0 [2]), .B(
        MCInst2_MC1_v2_0 [3]), .Z(Red_MCInst2_MC1_v2_2[0] ) );
  XOR2_X1 Red_MCInst2_MC1_v2_3Inst_0_U3  ( .A(MCInst2_MC1_v2_0 [2]), .B(
        MCInst2_MC1_v2_0 [0]), .Z(Red_MCInst2_MC1_v2_3[0] ) );
  XNOR2_X1 Red_MCInst2_MC1_v3_0Inst_0_U4  ( .A(
        Red_MCInst2_MC1_v3_0Inst_0_n2 ), .B(MCInst2_MC1_v3_0 [2]), .ZN(
        Red_MCInst2_MC1_v3_0[0] ) );
  XNOR2_X1 Red_MCInst2_MC1_v3_0Inst_0_U3  ( .A(Red_MCInst2_MC1_v3_1[0] ), 
        .B(MCInst2_MC1_v3_2 [3]), .ZN(Red_MCInst2_MC1_v3_0Inst_0_n2 ) );
  XNOR2_X1 Red_MCInst2_MC1_v3_2Inst_0_U4  ( .A(
        Red_MCInst2_MC1_v3_2Inst_0_n2 ), .B(Red_MCInst2_MC1_v3_1[0] ), .ZN(
        Red_MCInst2_MC1_v3_2[0] ) );
  XNOR2_X1 Red_MCInst2_MC1_v3_2Inst_0_U3  ( .A(MCInst2_MC1_v3_2 [2]), .B(
        MCInst2_MC1_v3_0 [2]), .ZN(Red_MCInst2_MC1_v3_2Inst_0_n2 ) );
  XOR2_X1 Red_MCInst2_MC1_v3_3Inst_0_U3  ( .A(MCInst2_MC1_v3_2 [3]), .B(
        MCInst2_MC1_v3_2 [2]), .Z(Red_MCInst2_MC1_v3_3[0] ) );
  XNOR2_X1 Red_MCInst2_MC1_r0Inst_XORInst_0_0_U3  ( .A(
        Red_MCInst2_MC1_r0Inst_XORInst_0_0_n5 ), .B(
        Red_MCInst2_MC1_r0Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback2[14]) );
  XNOR2_X1 Red_MCInst2_MC1_r0Inst_XORInst_0_0_U2  ( .A(
        Red_MCInst2_MC1_v3_0[0] ), .B(Red_MCInst2_MC1_v2_0[0] ), .ZN(
        Red_MCInst2_MC1_r0Inst_XORInst_0_0_n4 ) );
  XOR2_X1 Red_MCInst2_MC1_r0Inst_XORInst_0_0_U1  ( .A(
        Red_MCInst2_MC1_v0_0[0] ), .B(Red_MCInst2_MC1_v1_0[0] ), .Z(
        Red_MCInst2_MC1_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 Red_MCInst2_MC1_r1Inst_XORInst_0_0_U3  ( .A(
        Red_MCInst2_MC1_r1Inst_XORInst_0_0_n5 ), .B(
        Red_MCInst2_MC1_r1Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback2[10]) );
  XNOR2_X1 Red_MCInst2_MC1_r1Inst_XORInst_0_0_U2  ( .A(
        Red_MCInst2_MC1_v3_1[0] ), .B(Red_MCInst2_MC1_v2_1[0] ), .ZN(
        Red_MCInst2_MC1_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 Red_MCInst2_MC1_r1Inst_XORInst_0_0_U1  ( .A(
        Red_MCInst2_MC1_v0_1[0] ), .B(Red_MCInst2_MC1_v1_1[0] ), .Z(
        Red_MCInst2_MC1_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 Red_MCInst2_MC1_r2Inst_XORInst_0_0_U3  ( .A(
        Red_MCInst2_MC1_r2Inst_XORInst_0_0_n5 ), .B(
        Red_MCInst2_MC1_r2Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback2[6]) );
  XNOR2_X1 Red_MCInst2_MC1_r2Inst_XORInst_0_0_U2  ( .A(
        Red_MCInst2_MC1_v3_2[0] ), .B(Red_MCInst2_MC1_v2_2[0] ), .ZN(
        Red_MCInst2_MC1_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 Red_MCInst2_MC1_r2Inst_XORInst_0_0_U1  ( .A(
        Red_MCInst2_MC1_v0_2[0] ), .B(Red_MCInst2_MC1_v1_2[0] ), .Z(
        Red_MCInst2_MC1_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 Red_MCInst2_MC1_r3Inst_XORInst_0_0_U3  ( .A(
        Red_MCInst2_MC1_r3Inst_XORInst_0_0_n5 ), .B(
        Red_MCInst2_MC1_r3Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback2[2]) );
  XNOR2_X1 Red_MCInst2_MC1_r3Inst_XORInst_0_0_U2  ( .A(
        Red_MCInst2_MC1_v3_3[0] ), .B(Red_MCInst2_MC1_v2_3[0] ), .ZN(
        Red_MCInst2_MC1_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 Red_MCInst2_MC1_r3Inst_XORInst_0_0_U1  ( .A(
        Red_MCInst2_MC1_v0_3[0] ), .B(Red_MCInst2_MC1_v1_3[0] ), .Z(
        Red_MCInst2_MC1_r3Inst_XORInst_0_0_n5 ) );
  XOR2_X1 Red_MCInst2_MC2_v0_0Inst_0_U3  ( .A(Red_MCInst2_MC2_v0_1[0] ), .B(
        MCInst2_MC2_v0_0 [3]), .Z(Red_MCInst2_MC2_v0_0[0] ) );
  XOR2_X1 Red_MCInst2_MC2_v0_2Inst_0_U3  ( .A(Red_MCInst2_MC2_v0_1[0] ), .B(
        MCInst2_MC2_v0_3 [0]), .Z(Red_MCInst2_MC2_v0_2[0] ) );
  XNOR2_X1 Red_MCInst2_MC2_v0_3Inst_0_U4  ( .A(
        Red_MCInst2_MC2_v0_3Inst_0_n2 ), .B(MCInst2_MC2_v0_0 [3]), .ZN(
        Red_MCInst2_MC2_v0_3[0] ) );
  XNOR2_X1 Red_MCInst2_MC2_v0_3Inst_0_U3  ( .A(MCInst2_MC2_v0_3 [3]), .B(
        Red_MCInst2_MC2_v0_1[0] ), .ZN(Red_MCInst2_MC2_v0_3Inst_0_n2 ) );
  XNOR2_X1 Red_MCInst2_MC2_v1_0Inst_0_U5  ( .A(
        Red_MCInst2_MC2_v1_0Inst_0_n4 ), .B(Red_MCInst2_MC2_v1_0Inst_0_n3 ), 
        .ZN(Red_MCInst2_MC2_v1_0[0] ) );
  XNOR2_X1 Red_MCInst2_MC2_v1_0Inst_0_U4  ( .A(MCInst2_MC2_v1_3 [2]), .B(
        MCInst2_MC2_v1_0 [0]), .ZN(Red_MCInst2_MC2_v1_0Inst_0_n3 ) );
  XOR2_X1 Red_MCInst2_MC2_v1_0Inst_0_U3  ( .A(Red_MCInst2_MC2_v1_1[0] ), .B(
        MCInst2_MC2_v1_0 [3]), .Z(Red_MCInst2_MC2_v1_0Inst_0_n4 ) );
  XOR2_X1 Red_MCInst2_MC2_v1_2Inst_0_U3  ( .A(MCInst2_MC2_v1_0 [0]), .B(
        Red_MCInst2_MC2_v1_1[0] ), .Z(Red_MCInst2_MC2_v1_2[0] ) );
  XNOR2_X1 Red_MCInst2_MC2_v1_3Inst_0_U4  ( .A(
        Red_MCInst2_MC2_v1_3Inst_0_n2 ), .B(MCInst2_MC2_v1_3 [2]), .ZN(
        Red_MCInst2_MC2_v1_3[0] ) );
  XNOR2_X1 Red_MCInst2_MC2_v1_3Inst_0_U3  ( .A(Red_MCInst2_MC2_v1_1[0] ), 
        .B(MCInst2_MC2_v1_0 [0]), .ZN(Red_MCInst2_MC2_v1_3Inst_0_n2 ) );
  XNOR2_X1 Red_MCInst2_MC2_v2_0Inst_0_U4  ( .A(
        Red_MCInst2_MC2_v2_0Inst_0_n2 ), .B(MCInst2_MC2_v2_0 [2]), .ZN(
        Red_MCInst2_MC2_v2_0[0] ) );
  XNOR2_X1 Red_MCInst2_MC2_v2_0Inst_0_U3  ( .A(MCInst2_MC2_v2_0 [3]), .B(
        MCInst2_MC2_v2_3 [1]), .ZN(Red_MCInst2_MC2_v2_0Inst_0_n2 ) );
  XOR2_X1 Red_MCInst2_MC2_v2_1Inst_0_U3  ( .A(MCInst2_MC2_v2_0 [3]), .B(
        MCInst2_MC2_v2_0 [0]), .Z(Red_MCInst2_MC2_v2_1[0] ) );
  XOR2_X1 Red_MCInst2_MC2_v2_2Inst_0_U3  ( .A(MCInst2_MC2_v2_0 [2]), .B(
        MCInst2_MC2_v2_0 [3]), .Z(Red_MCInst2_MC2_v2_2[0] ) );
  XOR2_X1 Red_MCInst2_MC2_v2_3Inst_0_U3  ( .A(MCInst2_MC2_v2_0 [2]), .B(
        MCInst2_MC2_v2_0 [0]), .Z(Red_MCInst2_MC2_v2_3[0] ) );
  XNOR2_X1 Red_MCInst2_MC2_v3_0Inst_0_U4  ( .A(
        Red_MCInst2_MC2_v3_0Inst_0_n2 ), .B(MCInst2_MC2_v3_0 [2]), .ZN(
        Red_MCInst2_MC2_v3_0[0] ) );
  XNOR2_X1 Red_MCInst2_MC2_v3_0Inst_0_U3  ( .A(Red_MCInst2_MC2_v3_1[0] ), 
        .B(MCInst2_MC2_v3_2 [3]), .ZN(Red_MCInst2_MC2_v3_0Inst_0_n2 ) );
  XNOR2_X1 Red_MCInst2_MC2_v3_2Inst_0_U4  ( .A(
        Red_MCInst2_MC2_v3_2Inst_0_n2 ), .B(Red_MCInst2_MC2_v3_1[0] ), .ZN(
        Red_MCInst2_MC2_v3_2[0] ) );
  XNOR2_X1 Red_MCInst2_MC2_v3_2Inst_0_U3  ( .A(MCInst2_MC2_v3_2 [2]), .B(
        MCInst2_MC2_v3_0 [2]), .ZN(Red_MCInst2_MC2_v3_2Inst_0_n2 ) );
  XOR2_X1 Red_MCInst2_MC2_v3_3Inst_0_U3  ( .A(MCInst2_MC2_v3_2 [3]), .B(
        MCInst2_MC2_v3_2 [2]), .Z(Red_MCInst2_MC2_v3_3[0] ) );
  XNOR2_X1 Red_MCInst2_MC2_r0Inst_XORInst_0_0_U3  ( .A(
        Red_MCInst2_MC2_r0Inst_XORInst_0_0_n5 ), .B(
        Red_MCInst2_MC2_r0Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback2[13]) );
  XNOR2_X1 Red_MCInst2_MC2_r0Inst_XORInst_0_0_U2  ( .A(
        Red_MCInst2_MC2_v3_0[0] ), .B(Red_MCInst2_MC2_v2_0[0] ), .ZN(
        Red_MCInst2_MC2_r0Inst_XORInst_0_0_n4 ) );
  XOR2_X1 Red_MCInst2_MC2_r0Inst_XORInst_0_0_U1  ( .A(
        Red_MCInst2_MC2_v0_0[0] ), .B(Red_MCInst2_MC2_v1_0[0] ), .Z(
        Red_MCInst2_MC2_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 Red_MCInst2_MC2_r1Inst_XORInst_0_0_U3  ( .A(
        Red_MCInst2_MC2_r1Inst_XORInst_0_0_n5 ), .B(
        Red_MCInst2_MC2_r1Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback2[9]) );
  XNOR2_X1 Red_MCInst2_MC2_r1Inst_XORInst_0_0_U2  ( .A(
        Red_MCInst2_MC2_v3_1[0] ), .B(Red_MCInst2_MC2_v2_1[0] ), .ZN(
        Red_MCInst2_MC2_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 Red_MCInst2_MC2_r1Inst_XORInst_0_0_U1  ( .A(
        Red_MCInst2_MC2_v0_1[0] ), .B(Red_MCInst2_MC2_v1_1[0] ), .Z(
        Red_MCInst2_MC2_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 Red_MCInst2_MC2_r2Inst_XORInst_0_0_U3  ( .A(
        Red_MCInst2_MC2_r2Inst_XORInst_0_0_n5 ), .B(
        Red_MCInst2_MC2_r2Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback2[5]) );
  XNOR2_X1 Red_MCInst2_MC2_r2Inst_XORInst_0_0_U2  ( .A(
        Red_MCInst2_MC2_v3_2[0] ), .B(Red_MCInst2_MC2_v2_2[0] ), .ZN(
        Red_MCInst2_MC2_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 Red_MCInst2_MC2_r2Inst_XORInst_0_0_U1  ( .A(
        Red_MCInst2_MC2_v0_2[0] ), .B(Red_MCInst2_MC2_v1_2[0] ), .Z(
        Red_MCInst2_MC2_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 Red_MCInst2_MC2_r3Inst_XORInst_0_0_U3  ( .A(
        Red_MCInst2_MC2_r3Inst_XORInst_0_0_n5 ), .B(
        Red_MCInst2_MC2_r3Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback2[1]) );
  XNOR2_X1 Red_MCInst2_MC2_r3Inst_XORInst_0_0_U2  ( .A(
        Red_MCInst2_MC2_v3_3[0] ), .B(Red_MCInst2_MC2_v2_3[0] ), .ZN(
        Red_MCInst2_MC2_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 Red_MCInst2_MC2_r3Inst_XORInst_0_0_U1  ( .A(
        Red_MCInst2_MC2_v0_3[0] ), .B(Red_MCInst2_MC2_v1_3[0] ), .Z(
        Red_MCInst2_MC2_r3Inst_XORInst_0_0_n5 ) );
  XOR2_X1 Red_MCInst2_MC3_v0_0Inst_0_U3  ( .A(Red_MCInst2_MC3_v0_1[0] ), .B(
        MCInst2_MC3_v0_0 [3]), .Z(Red_MCInst2_MC3_v0_0[0] ) );
  XOR2_X1 Red_MCInst2_MC3_v0_2Inst_0_U3  ( .A(Red_MCInst2_MC3_v0_1[0] ), .B(
        MCInst2_MC3_v0_3 [0]), .Z(Red_MCInst2_MC3_v0_2[0] ) );
  XNOR2_X1 Red_MCInst2_MC3_v0_3Inst_0_U4  ( .A(
        Red_MCInst2_MC3_v0_3Inst_0_n2 ), .B(MCInst2_MC3_v0_0 [3]), .ZN(
        Red_MCInst2_MC3_v0_3[0] ) );
  XNOR2_X1 Red_MCInst2_MC3_v0_3Inst_0_U3  ( .A(MCInst2_MC3_v0_3 [3]), .B(
        Red_MCInst2_MC3_v0_1[0] ), .ZN(Red_MCInst2_MC3_v0_3Inst_0_n2 ) );
  XNOR2_X1 Red_MCInst2_MC3_v1_0Inst_0_U5  ( .A(
        Red_MCInst2_MC3_v1_0Inst_0_n4 ), .B(Red_MCInst2_MC3_v1_0Inst_0_n3 ), 
        .ZN(Red_MCInst2_MC3_v1_0[0] ) );
  XNOR2_X1 Red_MCInst2_MC3_v1_0Inst_0_U4  ( .A(MCInst2_MC3_v1_3 [2]), .B(
        MCInst2_MC3_v1_0 [0]), .ZN(Red_MCInst2_MC3_v1_0Inst_0_n3 ) );
  XOR2_X1 Red_MCInst2_MC3_v1_0Inst_0_U3  ( .A(Red_MCInst2_MC3_v1_1[0] ), .B(
        MCInst2_MC3_v1_0 [3]), .Z(Red_MCInst2_MC3_v1_0Inst_0_n4 ) );
  XOR2_X1 Red_MCInst2_MC3_v1_2Inst_0_U3  ( .A(MCInst2_MC3_v1_0 [0]), .B(
        Red_MCInst2_MC3_v1_1[0] ), .Z(Red_MCInst2_MC3_v1_2[0] ) );
  XNOR2_X1 Red_MCInst2_MC3_v1_3Inst_0_U4  ( .A(
        Red_MCInst2_MC3_v1_3Inst_0_n2 ), .B(MCInst2_MC3_v1_3 [2]), .ZN(
        Red_MCInst2_MC3_v1_3[0] ) );
  XNOR2_X1 Red_MCInst2_MC3_v1_3Inst_0_U3  ( .A(Red_MCInst2_MC3_v1_1[0] ), 
        .B(MCInst2_MC3_v1_0 [0]), .ZN(Red_MCInst2_MC3_v1_3Inst_0_n2 ) );
  XNOR2_X1 Red_MCInst2_MC3_v2_0Inst_0_U4  ( .A(
        Red_MCInst2_MC3_v2_0Inst_0_n2 ), .B(MCInst2_MC3_v2_0 [2]), .ZN(
        Red_MCInst2_MC3_v2_0[0] ) );
  XNOR2_X1 Red_MCInst2_MC3_v2_0Inst_0_U3  ( .A(MCInst2_MC3_v2_0 [3]), .B(
        MCInst2_MC3_v2_3 [1]), .ZN(Red_MCInst2_MC3_v2_0Inst_0_n2 ) );
  XOR2_X1 Red_MCInst2_MC3_v2_1Inst_0_U3  ( .A(MCInst2_MC3_v2_0 [3]), .B(
        MCInst2_MC3_v2_0 [0]), .Z(Red_MCInst2_MC3_v2_1[0] ) );
  XOR2_X1 Red_MCInst2_MC3_v2_2Inst_0_U3  ( .A(MCInst2_MC3_v2_0 [2]), .B(
        MCInst2_MC3_v2_0 [3]), .Z(Red_MCInst2_MC3_v2_2[0] ) );
  XOR2_X1 Red_MCInst2_MC3_v2_3Inst_0_U3  ( .A(MCInst2_MC3_v2_0 [2]), .B(
        MCInst2_MC3_v2_0 [0]), .Z(Red_MCInst2_MC3_v2_3[0] ) );
  XNOR2_X1 Red_MCInst2_MC3_v3_0Inst_0_U4  ( .A(
        Red_MCInst2_MC3_v3_0Inst_0_n2 ), .B(MCInst2_MC3_v3_0 [2]), .ZN(
        Red_MCInst2_MC3_v3_0[0] ) );
  XNOR2_X1 Red_MCInst2_MC3_v3_0Inst_0_U3  ( .A(Red_MCInst2_MC3_v3_1[0] ), 
        .B(MCInst2_MC3_v3_2 [3]), .ZN(Red_MCInst2_MC3_v3_0Inst_0_n2 ) );
  XNOR2_X1 Red_MCInst2_MC3_v3_2Inst_0_U4  ( .A(
        Red_MCInst2_MC3_v3_2Inst_0_n2 ), .B(Red_MCInst2_MC3_v3_1[0] ), .ZN(
        Red_MCInst2_MC3_v3_2[0] ) );
  XNOR2_X1 Red_MCInst2_MC3_v3_2Inst_0_U3  ( .A(MCInst2_MC3_v3_2 [2]), .B(
        MCInst2_MC3_v3_0 [2]), .ZN(Red_MCInst2_MC3_v3_2Inst_0_n2 ) );
  XOR2_X1 Red_MCInst2_MC3_v3_3Inst_0_U3  ( .A(MCInst2_MC3_v3_2 [3]), .B(
        MCInst2_MC3_v3_2 [2]), .Z(Red_MCInst2_MC3_v3_3[0] ) );
  XNOR2_X1 Red_MCInst2_MC3_r0Inst_XORInst_0_0_U3  ( .A(
        Red_MCInst2_MC3_r0Inst_XORInst_0_0_n5 ), .B(
        Red_MCInst2_MC3_r0Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback2[12]) );
  XNOR2_X1 Red_MCInst2_MC3_r0Inst_XORInst_0_0_U2  ( .A(
        Red_MCInst2_MC3_v3_0[0] ), .B(Red_MCInst2_MC3_v2_0[0] ), .ZN(
        Red_MCInst2_MC3_r0Inst_XORInst_0_0_n4 ) );
  XOR2_X1 Red_MCInst2_MC3_r0Inst_XORInst_0_0_U1  ( .A(
        Red_MCInst2_MC3_v0_0[0] ), .B(Red_MCInst2_MC3_v1_0[0] ), .Z(
        Red_MCInst2_MC3_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 Red_MCInst2_MC3_r1Inst_XORInst_0_0_U3  ( .A(
        Red_MCInst2_MC3_r1Inst_XORInst_0_0_n5 ), .B(
        Red_MCInst2_MC3_r1Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback2[8]) );
  XNOR2_X1 Red_MCInst2_MC3_r1Inst_XORInst_0_0_U2  ( .A(
        Red_MCInst2_MC3_v3_1[0] ), .B(Red_MCInst2_MC3_v2_1[0] ), .ZN(
        Red_MCInst2_MC3_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 Red_MCInst2_MC3_r1Inst_XORInst_0_0_U1  ( .A(
        Red_MCInst2_MC3_v0_1[0] ), .B(Red_MCInst2_MC3_v1_1[0] ), .Z(
        Red_MCInst2_MC3_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 Red_MCInst2_MC3_r2Inst_XORInst_0_0_U3  ( .A(
        Red_MCInst2_MC3_r2Inst_XORInst_0_0_n5 ), .B(
        Red_MCInst2_MC3_r2Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback2[4]) );
  XNOR2_X1 Red_MCInst2_MC3_r2Inst_XORInst_0_0_U2  ( .A(
        Red_MCInst2_MC3_v3_2[0] ), .B(Red_MCInst2_MC3_v2_2[0] ), .ZN(
        Red_MCInst2_MC3_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 Red_MCInst2_MC3_r2Inst_XORInst_0_0_U1  ( .A(
        Red_MCInst2_MC3_v0_2[0] ), .B(Red_MCInst2_MC3_v1_2[0] ), .Z(
        Red_MCInst2_MC3_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 Red_MCInst2_MC3_r3Inst_XORInst_0_0_U3  ( .A(
        Red_MCInst2_MC3_r3Inst_XORInst_0_0_n5 ), .B(
        Red_MCInst2_MC3_r3Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback2[0]) );
  XNOR2_X1 Red_MCInst2_MC3_r3Inst_XORInst_0_0_U2  ( .A(
        Red_MCInst2_MC3_v3_3[0] ), .B(Red_MCInst2_MC3_v2_3[0] ), .ZN(
        Red_MCInst2_MC3_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 Red_MCInst2_MC3_r3Inst_XORInst_0_0_U1  ( .A(
        Red_MCInst2_MC3_v0_3[0] ), .B(Red_MCInst2_MC3_v1_3[0] ), .Z(
        Red_MCInst2_MC3_r3Inst_XORInst_0_0_n5 ) );
  DFF_X1 RedStateReg2_s_current_state_reg[0]  ( .D(Red_Feedback2[0]), .CK(clk), .Q(Red_SubCellInput2[0]) );
  DFF_X1 RedStateReg2_s_current_state_reg[1]  ( .D(Red_Feedback2[1]), .CK(clk), .Q(Red_SubCellInput2[1]) );
  DFF_X1 RedStateReg2_s_current_state_reg[2]  ( .D(Red_Feedback2[2]), .CK(clk), .Q(Red_SubCellInput2[2]) );
  DFF_X1 RedStateReg2_s_current_state_reg[3]  ( .D(Red_Feedback2[3]), .CK(clk), .Q(Red_SubCellInput2[3]) );
  DFF_X1 RedStateReg2_s_current_state_reg[4]  ( .D(Red_Feedback2[4]), .CK(clk), .Q(Red_SubCellInput2[4]) );
  DFF_X1 RedStateReg2_s_current_state_reg[5]  ( .D(Red_Feedback2[5]), .CK(clk), .Q(Red_SubCellInput2[5]) );
  DFF_X1 RedStateReg2_s_current_state_reg[6]  ( .D(Red_Feedback2[6]), .CK(clk), .Q(Red_SubCellInput2[6]) );
  DFF_X1 RedStateReg2_s_current_state_reg[7]  ( .D(Red_Feedback2[7]), .CK(clk), .Q(Red_SubCellInput2[7]) );
  DFF_X1 RedStateReg2_s_current_state_reg[8]  ( .D(Red_Feedback2[8]), .CK(clk), .Q(Red_SubCellInput2[8]) );
  DFF_X1 RedStateReg2_s_current_state_reg[9]  ( .D(Red_Feedback2[9]), .CK(clk), .Q(Red_SubCellInput2[9]) );
  DFF_X1 RedStateReg2_s_current_state_reg[10]  ( .D(Red_Feedback2[10]), .CK(
        clk), .Q(Red_SubCellInput2[10]) );
  DFF_X1 RedStateReg2_s_current_state_reg[11]  ( .D(Red_Feedback2[11]), .CK(
        clk), .Q(Red_SubCellInput2[11]) );
  DFF_X1 RedStateReg2_s_current_state_reg[12]  ( .D(Red_Feedback2[12]), .CK(
        clk), .Q(Red_SubCellInput2[12]) );
  DFF_X1 RedStateReg2_s_current_state_reg[13]  ( .D(Red_Feedback2[13]), .CK(
        clk), .Q(Red_SubCellInput2[13]) );
  DFF_X1 RedStateReg2_s_current_state_reg[14]  ( .D(Red_Feedback2[14]), .CK(
        clk), .Q(Red_SubCellInput2[14]) );
  DFF_X1 RedStateReg2_s_current_state_reg[15]  ( .D(Red_Feedback2[15]), .CK(
        clk), .Q(Red_SubCellInput2[15]) );
  NAND2_X1 Red_SubCellInst3_LFInst_0_LFInst_0_U6  ( .A1(
        Red_SubCellInst3_LFInst_0_LFInst_0_n6 ), .A2(
        Red_SubCellInst3_LFInst_0_LFInst_0_n5 ), .ZN(Red_ShiftRowsOutput3[3])
         );
  NAND2_X1 Red_SubCellInst3_LFInst_0_LFInst_0_U5  ( .A1(SubCellInput2[3]), 
        .A2(SubCellInput2[2]), .ZN(Red_SubCellInst3_LFInst_0_LFInst_0_n5 ) );
  NAND2_X1 Red_SubCellInst3_LFInst_0_LFInst_0_U4  ( .A1(SubCellInput2[0]), 
        .A2(Red_SubCellInst3_LFInst_0_LFInst_0_n4 ), .ZN(
        Red_SubCellInst3_LFInst_0_LFInst_0_n6 ) );
  OR2_X1 Red_SubCellInst3_LFInst_0_LFInst_0_U3  ( .A1(SubCellInput2[1]), .A2(
        SubCellInput2[3]), .ZN(Red_SubCellInst3_LFInst_0_LFInst_0_n4 ) );
  NAND2_X1 Red_SubCellInst3_LFInst_1_LFInst_0_U6  ( .A1(
        Red_SubCellInst3_LFInst_1_LFInst_0_n6 ), .A2(
        Red_SubCellInst3_LFInst_1_LFInst_0_n5 ), .ZN(Red_ShiftRowsOutput3[0])
         );
  NAND2_X1 Red_SubCellInst3_LFInst_1_LFInst_0_U5  ( .A1(SubCellInput2[7]), 
        .A2(SubCellInput2[6]), .ZN(Red_SubCellInst3_LFInst_1_LFInst_0_n5 ) );
  NAND2_X1 Red_SubCellInst3_LFInst_1_LFInst_0_U4  ( .A1(SubCellInput2[4]), 
        .A2(Red_SubCellInst3_LFInst_1_LFInst_0_n4 ), .ZN(
        Red_SubCellInst3_LFInst_1_LFInst_0_n6 ) );
  OR2_X1 Red_SubCellInst3_LFInst_1_LFInst_0_U3  ( .A1(SubCellInput2[5]), .A2(
        SubCellInput2[7]), .ZN(Red_SubCellInst3_LFInst_1_LFInst_0_n4 ) );
  NAND2_X1 Red_SubCellInst3_LFInst_2_LFInst_0_U6  ( .A1(
        Red_SubCellInst3_LFInst_2_LFInst_0_n6 ), .A2(
        Red_SubCellInst3_LFInst_2_LFInst_0_n5 ), .ZN(Red_ShiftRowsOutput3[1])
         );
  NAND2_X1 Red_SubCellInst3_LFInst_2_LFInst_0_U5  ( .A1(SubCellInput2[11]), 
        .A2(SubCellInput2[10]), .ZN(Red_SubCellInst3_LFInst_2_LFInst_0_n5 )
         );
  NAND2_X1 Red_SubCellInst3_LFInst_2_LFInst_0_U4  ( .A1(SubCellInput2[8]), 
        .A2(Red_SubCellInst3_LFInst_2_LFInst_0_n4 ), .ZN(
        Red_SubCellInst3_LFInst_2_LFInst_0_n6 ) );
  OR2_X1 Red_SubCellInst3_LFInst_2_LFInst_0_U3  ( .A1(SubCellInput2[9]), .A2(
        SubCellInput2[11]), .ZN(Red_SubCellInst3_LFInst_2_LFInst_0_n4 ) );
  NAND2_X1 Red_SubCellInst3_LFInst_3_LFInst_0_U6  ( .A1(
        Red_SubCellInst3_LFInst_3_LFInst_0_n6 ), .A2(
        Red_SubCellInst3_LFInst_3_LFInst_0_n5 ), .ZN(Red_ShiftRowsOutput3[2])
         );
  NAND2_X1 Red_SubCellInst3_LFInst_3_LFInst_0_U5  ( .A1(SubCellInput2[15]), 
        .A2(SubCellInput2[14]), .ZN(Red_SubCellInst3_LFInst_3_LFInst_0_n5 )
         );
  NAND2_X1 Red_SubCellInst3_LFInst_3_LFInst_0_U4  ( .A1(SubCellInput2[12]), 
        .A2(Red_SubCellInst3_LFInst_3_LFInst_0_n4 ), .ZN(
        Red_SubCellInst3_LFInst_3_LFInst_0_n6 ) );
  OR2_X1 Red_SubCellInst3_LFInst_3_LFInst_0_U3  ( .A1(SubCellInput2[13]), 
        .A2(SubCellInput2[15]), .ZN(Red_SubCellInst3_LFInst_3_LFInst_0_n4 )
         );
  NAND2_X1 Red_SubCellInst3_LFInst_4_LFInst_0_U6  ( .A1(
        Red_SubCellInst3_LFInst_4_LFInst_0_n6 ), .A2(
        Red_SubCellInst3_LFInst_4_LFInst_0_n5 ), .ZN(Red_ShiftRowsOutput3[6])
         );
  NAND2_X1 Red_SubCellInst3_LFInst_4_LFInst_0_U5  ( .A1(SubCellInput2[19]), 
        .A2(SubCellInput2[18]), .ZN(Red_SubCellInst3_LFInst_4_LFInst_0_n5 )
         );
  NAND2_X1 Red_SubCellInst3_LFInst_4_LFInst_0_U4  ( .A1(SubCellInput2[16]), 
        .A2(Red_SubCellInst3_LFInst_4_LFInst_0_n4 ), .ZN(
        Red_SubCellInst3_LFInst_4_LFInst_0_n6 ) );
  OR2_X1 Red_SubCellInst3_LFInst_4_LFInst_0_U3  ( .A1(SubCellInput2[17]), 
        .A2(SubCellInput2[19]), .ZN(Red_SubCellInst3_LFInst_4_LFInst_0_n4 )
         );
  NAND2_X1 Red_SubCellInst3_LFInst_5_LFInst_0_U6  ( .A1(
        Red_SubCellInst3_LFInst_5_LFInst_0_n6 ), .A2(
        Red_SubCellInst3_LFInst_5_LFInst_0_n5 ), .ZN(Red_ShiftRowsOutput3[7])
         );
  NAND2_X1 Red_SubCellInst3_LFInst_5_LFInst_0_U5  ( .A1(SubCellInput2[23]), 
        .A2(SubCellInput2[22]), .ZN(Red_SubCellInst3_LFInst_5_LFInst_0_n5 )
         );
  NAND2_X1 Red_SubCellInst3_LFInst_5_LFInst_0_U4  ( .A1(SubCellInput2[20]), 
        .A2(Red_SubCellInst3_LFInst_5_LFInst_0_n4 ), .ZN(
        Red_SubCellInst3_LFInst_5_LFInst_0_n6 ) );
  OR2_X1 Red_SubCellInst3_LFInst_5_LFInst_0_U3  ( .A1(SubCellInput2[21]), 
        .A2(SubCellInput2[23]), .ZN(Red_SubCellInst3_LFInst_5_LFInst_0_n4 )
         );
  NAND2_X1 Red_SubCellInst3_LFInst_6_LFInst_0_U6  ( .A1(
        Red_SubCellInst3_LFInst_6_LFInst_0_n6 ), .A2(
        Red_SubCellInst3_LFInst_6_LFInst_0_n5 ), .ZN(Red_ShiftRowsOutput3[4])
         );
  NAND2_X1 Red_SubCellInst3_LFInst_6_LFInst_0_U5  ( .A1(SubCellInput2[27]), 
        .A2(SubCellInput2[26]), .ZN(Red_SubCellInst3_LFInst_6_LFInst_0_n5 )
         );
  NAND2_X1 Red_SubCellInst3_LFInst_6_LFInst_0_U4  ( .A1(SubCellInput2[24]), 
        .A2(Red_SubCellInst3_LFInst_6_LFInst_0_n4 ), .ZN(
        Red_SubCellInst3_LFInst_6_LFInst_0_n6 ) );
  OR2_X1 Red_SubCellInst3_LFInst_6_LFInst_0_U3  ( .A1(SubCellInput2[25]), 
        .A2(SubCellInput2[27]), .ZN(Red_SubCellInst3_LFInst_6_LFInst_0_n4 )
         );
  NAND2_X1 Red_SubCellInst3_LFInst_7_LFInst_0_U6  ( .A1(
        Red_SubCellInst3_LFInst_7_LFInst_0_n6 ), .A2(
        Red_SubCellInst3_LFInst_7_LFInst_0_n5 ), .ZN(Red_ShiftRowsOutput3[5])
         );
  NAND2_X1 Red_SubCellInst3_LFInst_7_LFInst_0_U5  ( .A1(SubCellInput2[31]), 
        .A2(SubCellInput2[30]), .ZN(Red_SubCellInst3_LFInst_7_LFInst_0_n5 )
         );
  NAND2_X1 Red_SubCellInst3_LFInst_7_LFInst_0_U4  ( .A1(SubCellInput2[28]), 
        .A2(Red_SubCellInst3_LFInst_7_LFInst_0_n4 ), .ZN(
        Red_SubCellInst3_LFInst_7_LFInst_0_n6 ) );
  OR2_X1 Red_SubCellInst3_LFInst_7_LFInst_0_U3  ( .A1(SubCellInput2[29]), 
        .A2(SubCellInput2[31]), .ZN(Red_SubCellInst3_LFInst_7_LFInst_0_n4 )
         );
  NAND2_X1 Red_SubCellInst3_LFInst_8_LFInst_0_U6  ( .A1(
        Red_SubCellInst3_LFInst_8_LFInst_0_n6 ), .A2(
        Red_SubCellInst3_LFInst_8_LFInst_0_n5 ), .ZN(Red_ShiftRowsOutput3[9])
         );
  NAND2_X1 Red_SubCellInst3_LFInst_8_LFInst_0_U5  ( .A1(SubCellInput2[35]), 
        .A2(SubCellInput2[34]), .ZN(Red_SubCellInst3_LFInst_8_LFInst_0_n5 )
         );
  NAND2_X1 Red_SubCellInst3_LFInst_8_LFInst_0_U4  ( .A1(SubCellInput2[32]), 
        .A2(Red_SubCellInst3_LFInst_8_LFInst_0_n4 ), .ZN(
        Red_SubCellInst3_LFInst_8_LFInst_0_n6 ) );
  OR2_X1 Red_SubCellInst3_LFInst_8_LFInst_0_U3  ( .A1(SubCellInput2[33]), 
        .A2(SubCellInput2[35]), .ZN(Red_SubCellInst3_LFInst_8_LFInst_0_n4 )
         );
  NAND2_X1 Red_SubCellInst3_LFInst_9_LFInst_0_U6  ( .A1(
        Red_SubCellInst3_LFInst_9_LFInst_0_n6 ), .A2(
        Red_SubCellInst3_LFInst_9_LFInst_0_n5 ), .ZN(Red_ShiftRowsOutput3[10]) );
  NAND2_X1 Red_SubCellInst3_LFInst_9_LFInst_0_U5  ( .A1(SubCellInput2[39]), 
        .A2(SubCellInput2[38]), .ZN(Red_SubCellInst3_LFInst_9_LFInst_0_n5 )
         );
  NAND2_X1 Red_SubCellInst3_LFInst_9_LFInst_0_U4  ( .A1(SubCellInput2[36]), 
        .A2(Red_SubCellInst3_LFInst_9_LFInst_0_n4 ), .ZN(
        Red_SubCellInst3_LFInst_9_LFInst_0_n6 ) );
  OR2_X1 Red_SubCellInst3_LFInst_9_LFInst_0_U3  ( .A1(SubCellInput2[37]), 
        .A2(SubCellInput2[39]), .ZN(Red_SubCellInst3_LFInst_9_LFInst_0_n4 )
         );
  NAND2_X1 Red_SubCellInst3_LFInst_10_LFInst_0_U6  ( .A1(
        Red_SubCellInst3_LFInst_10_LFInst_0_n6 ), .A2(
        Red_SubCellInst3_LFInst_10_LFInst_0_n5 ), .ZN(
        Red_ShiftRowsOutput3[11]) );
  NAND2_X1 Red_SubCellInst3_LFInst_10_LFInst_0_U5  ( .A1(SubCellInput2[43]), 
        .A2(SubCellInput2[42]), .ZN(Red_SubCellInst3_LFInst_10_LFInst_0_n5 )
         );
  NAND2_X1 Red_SubCellInst3_LFInst_10_LFInst_0_U4  ( .A1(SubCellInput2[40]), 
        .A2(Red_SubCellInst3_LFInst_10_LFInst_0_n4 ), .ZN(
        Red_SubCellInst3_LFInst_10_LFInst_0_n6 ) );
  OR2_X1 Red_SubCellInst3_LFInst_10_LFInst_0_U3  ( .A1(SubCellInput2[41]), 
        .A2(SubCellInput2[43]), .ZN(Red_SubCellInst3_LFInst_10_LFInst_0_n4 )
         );
  NAND2_X1 Red_SubCellInst3_LFInst_11_LFInst_0_U6  ( .A1(
        Red_SubCellInst3_LFInst_11_LFInst_0_n6 ), .A2(
        Red_SubCellInst3_LFInst_11_LFInst_0_n5 ), .ZN(Red_ShiftRowsOutput3[8]) );
  NAND2_X1 Red_SubCellInst3_LFInst_11_LFInst_0_U5  ( .A1(SubCellInput2[47]), 
        .A2(SubCellInput2[46]), .ZN(Red_SubCellInst3_LFInst_11_LFInst_0_n5 )
         );
  NAND2_X1 Red_SubCellInst3_LFInst_11_LFInst_0_U4  ( .A1(SubCellInput2[44]), 
        .A2(Red_SubCellInst3_LFInst_11_LFInst_0_n4 ), .ZN(
        Red_SubCellInst3_LFInst_11_LFInst_0_n6 ) );
  OR2_X1 Red_SubCellInst3_LFInst_11_LFInst_0_U3  ( .A1(SubCellInput2[45]), 
        .A2(SubCellInput2[47]), .ZN(Red_SubCellInst3_LFInst_11_LFInst_0_n4 )
         );
  NAND2_X1 Red_SubCellInst3_LFInst_12_LFInst_0_U6  ( .A1(
        Red_SubCellInst3_LFInst_12_LFInst_0_n6 ), .A2(
        Red_SubCellInst3_LFInst_12_LFInst_0_n5 ), .ZN(
        Red_ShiftRowsOutput3[12]) );
  NAND2_X1 Red_SubCellInst3_LFInst_12_LFInst_0_U5  ( .A1(SubCellInput2[51]), 
        .A2(SubCellInput2[50]), .ZN(Red_SubCellInst3_LFInst_12_LFInst_0_n5 )
         );
  NAND2_X1 Red_SubCellInst3_LFInst_12_LFInst_0_U4  ( .A1(SubCellInput2[48]), 
        .A2(Red_SubCellInst3_LFInst_12_LFInst_0_n4 ), .ZN(
        Red_SubCellInst3_LFInst_12_LFInst_0_n6 ) );
  OR2_X1 Red_SubCellInst3_LFInst_12_LFInst_0_U3  ( .A1(SubCellInput2[49]), 
        .A2(SubCellInput2[51]), .ZN(Red_SubCellInst3_LFInst_12_LFInst_0_n4 )
         );
  NAND2_X1 Red_SubCellInst3_LFInst_13_LFInst_0_U6  ( .A1(
        Red_SubCellInst3_LFInst_13_LFInst_0_n6 ), .A2(
        Red_SubCellInst3_LFInst_13_LFInst_0_n5 ), .ZN(
        Red_ShiftRowsOutput3[13]) );
  NAND2_X1 Red_SubCellInst3_LFInst_13_LFInst_0_U5  ( .A1(SubCellInput2[55]), 
        .A2(SubCellInput2[54]), .ZN(Red_SubCellInst3_LFInst_13_LFInst_0_n5 )
         );
  NAND2_X1 Red_SubCellInst3_LFInst_13_LFInst_0_U4  ( .A1(SubCellInput2[52]), 
        .A2(Red_SubCellInst3_LFInst_13_LFInst_0_n4 ), .ZN(
        Red_SubCellInst3_LFInst_13_LFInst_0_n6 ) );
  OR2_X1 Red_SubCellInst3_LFInst_13_LFInst_0_U3  ( .A1(SubCellInput2[53]), 
        .A2(SubCellInput2[55]), .ZN(Red_SubCellInst3_LFInst_13_LFInst_0_n4 )
         );
  NAND2_X1 Red_SubCellInst3_LFInst_14_LFInst_0_U6  ( .A1(
        Red_SubCellInst3_LFInst_14_LFInst_0_n6 ), .A2(
        Red_SubCellInst3_LFInst_14_LFInst_0_n5 ), .ZN(
        Red_ShiftRowsOutput3[14]) );
  NAND2_X1 Red_SubCellInst3_LFInst_14_LFInst_0_U5  ( .A1(SubCellInput2[59]), 
        .A2(SubCellInput2[58]), .ZN(Red_SubCellInst3_LFInst_14_LFInst_0_n5 )
         );
  NAND2_X1 Red_SubCellInst3_LFInst_14_LFInst_0_U4  ( .A1(SubCellInput2[56]), 
        .A2(Red_SubCellInst3_LFInst_14_LFInst_0_n4 ), .ZN(
        Red_SubCellInst3_LFInst_14_LFInst_0_n6 ) );
  OR2_X1 Red_SubCellInst3_LFInst_14_LFInst_0_U3  ( .A1(SubCellInput2[57]), 
        .A2(SubCellInput2[59]), .ZN(Red_SubCellInst3_LFInst_14_LFInst_0_n4 )
         );
  NAND2_X1 Red_SubCellInst3_LFInst_15_LFInst_0_U6  ( .A1(
        Red_SubCellInst3_LFInst_15_LFInst_0_n6 ), .A2(
        Red_SubCellInst3_LFInst_15_LFInst_0_n5 ), .ZN(
        Red_ShiftRowsOutput3[15]) );
  NAND2_X1 Red_SubCellInst3_LFInst_15_LFInst_0_U5  ( .A1(SubCellInput2[63]), 
        .A2(SubCellInput2[62]), .ZN(Red_SubCellInst3_LFInst_15_LFInst_0_n5 )
         );
  NAND2_X1 Red_SubCellInst3_LFInst_15_LFInst_0_U4  ( .A1(SubCellInput2[60]), 
        .A2(Red_SubCellInst3_LFInst_15_LFInst_0_n4 ), .ZN(
        Red_SubCellInst3_LFInst_15_LFInst_0_n6 ) );
  OR2_X1 Red_SubCellInst3_LFInst_15_LFInst_0_U3  ( .A1(SubCellInput2[61]), 
        .A2(SubCellInput2[63]), .ZN(Red_SubCellInst3_LFInst_15_LFInst_0_n4 )
         );
  XOR2_X1 Red_MCInst3_MC0_v0_0Inst_0_U3  ( .A(Red_MCInst3_MC0_v0_1[0] ), .B(
        MCInst3_MC0_v0_0 [3]), .Z(Red_MCInst3_MC0_v0_0[0] ) );
  XOR2_X1 Red_MCInst3_MC0_v0_2Inst_0_U3  ( .A(Red_MCInst3_MC0_v0_1[0] ), .B(
        MCInst3_MC0_v0_3 [0]), .Z(Red_MCInst3_MC0_v0_2[0] ) );
  XNOR2_X1 Red_MCInst3_MC0_v0_3Inst_0_U4  ( .A(
        Red_MCInst3_MC0_v0_3Inst_0_n2 ), .B(MCInst3_MC0_v0_0 [3]), .ZN(
        Red_MCInst3_MC0_v0_3[0] ) );
  XNOR2_X1 Red_MCInst3_MC0_v0_3Inst_0_U3  ( .A(MCInst3_MC0_v0_3 [3]), .B(
        Red_MCInst3_MC0_v0_1[0] ), .ZN(Red_MCInst3_MC0_v0_3Inst_0_n2 ) );
  XNOR2_X1 Red_MCInst3_MC0_v1_0Inst_0_U5  ( .A(
        Red_MCInst3_MC0_v1_0Inst_0_n4 ), .B(Red_MCInst3_MC0_v1_0Inst_0_n3 ), 
        .ZN(Red_MCInst3_MC0_v1_0[0] ) );
  XNOR2_X1 Red_MCInst3_MC0_v1_0Inst_0_U4  ( .A(MCInst3_MC0_v1_3 [2]), .B(
        MCInst3_MC0_v1_0 [0]), .ZN(Red_MCInst3_MC0_v1_0Inst_0_n3 ) );
  XOR2_X1 Red_MCInst3_MC0_v1_0Inst_0_U3  ( .A(Red_MCInst3_MC0_v1_1[0] ), .B(
        MCInst3_MC0_v1_0 [3]), .Z(Red_MCInst3_MC0_v1_0Inst_0_n4 ) );
  XOR2_X1 Red_MCInst3_MC0_v1_2Inst_0_U3  ( .A(MCInst3_MC0_v1_0 [0]), .B(
        Red_MCInst3_MC0_v1_1[0] ), .Z(Red_MCInst3_MC0_v1_2[0] ) );
  XNOR2_X1 Red_MCInst3_MC0_v1_3Inst_0_U4  ( .A(
        Red_MCInst3_MC0_v1_3Inst_0_n2 ), .B(MCInst3_MC0_v1_3 [2]), .ZN(
        Red_MCInst3_MC0_v1_3[0] ) );
  XNOR2_X1 Red_MCInst3_MC0_v1_3Inst_0_U3  ( .A(Red_MCInst3_MC0_v1_1[0] ), 
        .B(MCInst3_MC0_v1_0 [0]), .ZN(Red_MCInst3_MC0_v1_3Inst_0_n2 ) );
  XNOR2_X1 Red_MCInst3_MC0_v2_0Inst_0_U4  ( .A(
        Red_MCInst3_MC0_v2_0Inst_0_n2 ), .B(MCInst3_MC0_v2_0 [2]), .ZN(
        Red_MCInst3_MC0_v2_0[0] ) );
  XNOR2_X1 Red_MCInst3_MC0_v2_0Inst_0_U3  ( .A(MCInst3_MC0_v2_0 [3]), .B(
        MCInst3_MC0_v2_3 [1]), .ZN(Red_MCInst3_MC0_v2_0Inst_0_n2 ) );
  XOR2_X1 Red_MCInst3_MC0_v2_1Inst_0_U3  ( .A(MCInst3_MC0_v2_0 [3]), .B(
        MCInst3_MC0_v2_0 [0]), .Z(Red_MCInst3_MC0_v2_1[0] ) );
  XOR2_X1 Red_MCInst3_MC0_v2_2Inst_0_U3  ( .A(MCInst3_MC0_v2_0 [2]), .B(
        MCInst3_MC0_v2_0 [3]), .Z(Red_MCInst3_MC0_v2_2[0] ) );
  XOR2_X1 Red_MCInst3_MC0_v2_3Inst_0_U3  ( .A(MCInst3_MC0_v2_0 [2]), .B(
        MCInst3_MC0_v2_0 [0]), .Z(Red_MCInst3_MC0_v2_3[0] ) );
  XNOR2_X1 Red_MCInst3_MC0_v3_0Inst_0_U4  ( .A(
        Red_MCInst3_MC0_v3_0Inst_0_n2 ), .B(MCInst3_MC0_v3_0 [2]), .ZN(
        Red_MCInst3_MC0_v3_0[0] ) );
  XNOR2_X1 Red_MCInst3_MC0_v3_0Inst_0_U3  ( .A(Red_MCInst3_MC0_v3_1[0] ), 
        .B(MCInst3_MC0_v3_2 [3]), .ZN(Red_MCInst3_MC0_v3_0Inst_0_n2 ) );
  XNOR2_X1 Red_MCInst3_MC0_v3_2Inst_0_U4  ( .A(
        Red_MCInst3_MC0_v3_2Inst_0_n2 ), .B(Red_MCInst3_MC0_v3_1[0] ), .ZN(
        Red_MCInst3_MC0_v3_2[0] ) );
  XNOR2_X1 Red_MCInst3_MC0_v3_2Inst_0_U3  ( .A(MCInst3_MC0_v3_2 [2]), .B(
        MCInst3_MC0_v3_0 [2]), .ZN(Red_MCInst3_MC0_v3_2Inst_0_n2 ) );
  XOR2_X1 Red_MCInst3_MC0_v3_3Inst_0_U3  ( .A(MCInst3_MC0_v3_2 [3]), .B(
        MCInst3_MC0_v3_2 [2]), .Z(Red_MCInst3_MC0_v3_3[0] ) );
  XNOR2_X1 Red_MCInst3_MC0_r0Inst_XORInst_0_0_U3  ( .A(
        Red_MCInst3_MC0_r0Inst_XORInst_0_0_n5 ), .B(
        Red_MCInst3_MC0_r0Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback3[15]) );
  XNOR2_X1 Red_MCInst3_MC0_r0Inst_XORInst_0_0_U2  ( .A(
        Red_MCInst3_MC0_v3_0[0] ), .B(Red_MCInst3_MC0_v2_0[0] ), .ZN(
        Red_MCInst3_MC0_r0Inst_XORInst_0_0_n4 ) );
  XOR2_X1 Red_MCInst3_MC0_r0Inst_XORInst_0_0_U1  ( .A(
        Red_MCInst3_MC0_v0_0[0] ), .B(Red_MCInst3_MC0_v1_0[0] ), .Z(
        Red_MCInst3_MC0_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 Red_MCInst3_MC0_r1Inst_XORInst_0_0_U3  ( .A(
        Red_MCInst3_MC0_r1Inst_XORInst_0_0_n5 ), .B(
        Red_MCInst3_MC0_r1Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback3[11]) );
  XNOR2_X1 Red_MCInst3_MC0_r1Inst_XORInst_0_0_U2  ( .A(
        Red_MCInst3_MC0_v3_1[0] ), .B(Red_MCInst3_MC0_v2_1[0] ), .ZN(
        Red_MCInst3_MC0_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 Red_MCInst3_MC0_r1Inst_XORInst_0_0_U1  ( .A(
        Red_MCInst3_MC0_v0_1[0] ), .B(Red_MCInst3_MC0_v1_1[0] ), .Z(
        Red_MCInst3_MC0_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 Red_MCInst3_MC0_r2Inst_XORInst_0_0_U3  ( .A(
        Red_MCInst3_MC0_r2Inst_XORInst_0_0_n5 ), .B(
        Red_MCInst3_MC0_r2Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback3[7]) );
  XNOR2_X1 Red_MCInst3_MC0_r2Inst_XORInst_0_0_U2  ( .A(
        Red_MCInst3_MC0_v3_2[0] ), .B(Red_MCInst3_MC0_v2_2[0] ), .ZN(
        Red_MCInst3_MC0_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 Red_MCInst3_MC0_r2Inst_XORInst_0_0_U1  ( .A(
        Red_MCInst3_MC0_v0_2[0] ), .B(Red_MCInst3_MC0_v1_2[0] ), .Z(
        Red_MCInst3_MC0_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 Red_MCInst3_MC0_r3Inst_XORInst_0_0_U3  ( .A(
        Red_MCInst3_MC0_r3Inst_XORInst_0_0_n5 ), .B(
        Red_MCInst3_MC0_r3Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback3[3]) );
  XNOR2_X1 Red_MCInst3_MC0_r3Inst_XORInst_0_0_U2  ( .A(
        Red_MCInst3_MC0_v3_3[0] ), .B(Red_MCInst3_MC0_v2_3[0] ), .ZN(
        Red_MCInst3_MC0_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 Red_MCInst3_MC0_r3Inst_XORInst_0_0_U1  ( .A(
        Red_MCInst3_MC0_v0_3[0] ), .B(Red_MCInst3_MC0_v1_3[0] ), .Z(
        Red_MCInst3_MC0_r3Inst_XORInst_0_0_n5 ) );
  XOR2_X1 Red_MCInst3_MC1_v0_0Inst_0_U3  ( .A(Red_MCInst3_MC1_v0_1[0] ), .B(
        MCInst3_MC1_v0_0 [3]), .Z(Red_MCInst3_MC1_v0_0[0] ) );
  XOR2_X1 Red_MCInst3_MC1_v0_2Inst_0_U3  ( .A(Red_MCInst3_MC1_v0_1[0] ), .B(
        MCInst3_MC1_v0_3 [0]), .Z(Red_MCInst3_MC1_v0_2[0] ) );
  XNOR2_X1 Red_MCInst3_MC1_v0_3Inst_0_U4  ( .A(
        Red_MCInst3_MC1_v0_3Inst_0_n2 ), .B(MCInst3_MC1_v0_0 [3]), .ZN(
        Red_MCInst3_MC1_v0_3[0] ) );
  XNOR2_X1 Red_MCInst3_MC1_v0_3Inst_0_U3  ( .A(MCInst3_MC1_v0_3 [3]), .B(
        Red_MCInst3_MC1_v0_1[0] ), .ZN(Red_MCInst3_MC1_v0_3Inst_0_n2 ) );
  XNOR2_X1 Red_MCInst3_MC1_v1_0Inst_0_U5  ( .A(
        Red_MCInst3_MC1_v1_0Inst_0_n4 ), .B(Red_MCInst3_MC1_v1_0Inst_0_n3 ), 
        .ZN(Red_MCInst3_MC1_v1_0[0] ) );
  XNOR2_X1 Red_MCInst3_MC1_v1_0Inst_0_U4  ( .A(MCInst3_MC1_v1_3 [2]), .B(
        MCInst3_MC1_v1_0 [0]), .ZN(Red_MCInst3_MC1_v1_0Inst_0_n3 ) );
  XOR2_X1 Red_MCInst3_MC1_v1_0Inst_0_U3  ( .A(Red_MCInst3_MC1_v1_1[0] ), .B(
        MCInst3_MC1_v1_0 [3]), .Z(Red_MCInst3_MC1_v1_0Inst_0_n4 ) );
  XOR2_X1 Red_MCInst3_MC1_v1_2Inst_0_U3  ( .A(MCInst3_MC1_v1_0 [0]), .B(
        Red_MCInst3_MC1_v1_1[0] ), .Z(Red_MCInst3_MC1_v1_2[0] ) );
  XNOR2_X1 Red_MCInst3_MC1_v1_3Inst_0_U4  ( .A(
        Red_MCInst3_MC1_v1_3Inst_0_n2 ), .B(MCInst3_MC1_v1_3 [2]), .ZN(
        Red_MCInst3_MC1_v1_3[0] ) );
  XNOR2_X1 Red_MCInst3_MC1_v1_3Inst_0_U3  ( .A(Red_MCInst3_MC1_v1_1[0] ), 
        .B(MCInst3_MC1_v1_0 [0]), .ZN(Red_MCInst3_MC1_v1_3Inst_0_n2 ) );
  XNOR2_X1 Red_MCInst3_MC1_v2_0Inst_0_U4  ( .A(
        Red_MCInst3_MC1_v2_0Inst_0_n2 ), .B(MCInst3_MC1_v2_0 [2]), .ZN(
        Red_MCInst3_MC1_v2_0[0] ) );
  XNOR2_X1 Red_MCInst3_MC1_v2_0Inst_0_U3  ( .A(MCInst3_MC1_v2_0 [3]), .B(
        MCInst3_MC1_v2_3 [1]), .ZN(Red_MCInst3_MC1_v2_0Inst_0_n2 ) );
  XOR2_X1 Red_MCInst3_MC1_v2_1Inst_0_U3  ( .A(MCInst3_MC1_v2_0 [3]), .B(
        MCInst3_MC1_v2_0 [0]), .Z(Red_MCInst3_MC1_v2_1[0] ) );
  XOR2_X1 Red_MCInst3_MC1_v2_2Inst_0_U3  ( .A(MCInst3_MC1_v2_0 [2]), .B(
        MCInst3_MC1_v2_0 [3]), .Z(Red_MCInst3_MC1_v2_2[0] ) );
  XOR2_X1 Red_MCInst3_MC1_v2_3Inst_0_U3  ( .A(MCInst3_MC1_v2_0 [2]), .B(
        MCInst3_MC1_v2_0 [0]), .Z(Red_MCInst3_MC1_v2_3[0] ) );
  XNOR2_X1 Red_MCInst3_MC1_v3_0Inst_0_U4  ( .A(
        Red_MCInst3_MC1_v3_0Inst_0_n2 ), .B(MCInst3_MC1_v3_0 [2]), .ZN(
        Red_MCInst3_MC1_v3_0[0] ) );
  XNOR2_X1 Red_MCInst3_MC1_v3_0Inst_0_U3  ( .A(Red_MCInst3_MC1_v3_1[0] ), 
        .B(MCInst3_MC1_v3_2 [3]), .ZN(Red_MCInst3_MC1_v3_0Inst_0_n2 ) );
  XNOR2_X1 Red_MCInst3_MC1_v3_2Inst_0_U4  ( .A(
        Red_MCInst3_MC1_v3_2Inst_0_n2 ), .B(Red_MCInst3_MC1_v3_1[0] ), .ZN(
        Red_MCInst3_MC1_v3_2[0] ) );
  XNOR2_X1 Red_MCInst3_MC1_v3_2Inst_0_U3  ( .A(MCInst3_MC1_v3_2 [2]), .B(
        MCInst3_MC1_v3_0 [2]), .ZN(Red_MCInst3_MC1_v3_2Inst_0_n2 ) );
  XOR2_X1 Red_MCInst3_MC1_v3_3Inst_0_U3  ( .A(MCInst3_MC1_v3_2 [3]), .B(
        MCInst3_MC1_v3_2 [2]), .Z(Red_MCInst3_MC1_v3_3[0] ) );
  XNOR2_X1 Red_MCInst3_MC1_r0Inst_XORInst_0_0_U3  ( .A(
        Red_MCInst3_MC1_r0Inst_XORInst_0_0_n5 ), .B(
        Red_MCInst3_MC1_r0Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback3[14]) );
  XNOR2_X1 Red_MCInst3_MC1_r0Inst_XORInst_0_0_U2  ( .A(
        Red_MCInst3_MC1_v3_0[0] ), .B(Red_MCInst3_MC1_v2_0[0] ), .ZN(
        Red_MCInst3_MC1_r0Inst_XORInst_0_0_n4 ) );
  XOR2_X1 Red_MCInst3_MC1_r0Inst_XORInst_0_0_U1  ( .A(
        Red_MCInst3_MC1_v0_0[0] ), .B(Red_MCInst3_MC1_v1_0[0] ), .Z(
        Red_MCInst3_MC1_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 Red_MCInst3_MC1_r1Inst_XORInst_0_0_U3  ( .A(
        Red_MCInst3_MC1_r1Inst_XORInst_0_0_n5 ), .B(
        Red_MCInst3_MC1_r1Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback3[10]) );
  XNOR2_X1 Red_MCInst3_MC1_r1Inst_XORInst_0_0_U2  ( .A(
        Red_MCInst3_MC1_v3_1[0] ), .B(Red_MCInst3_MC1_v2_1[0] ), .ZN(
        Red_MCInst3_MC1_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 Red_MCInst3_MC1_r1Inst_XORInst_0_0_U1  ( .A(
        Red_MCInst3_MC1_v0_1[0] ), .B(Red_MCInst3_MC1_v1_1[0] ), .Z(
        Red_MCInst3_MC1_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 Red_MCInst3_MC1_r2Inst_XORInst_0_0_U3  ( .A(
        Red_MCInst3_MC1_r2Inst_XORInst_0_0_n5 ), .B(
        Red_MCInst3_MC1_r2Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback3[6]) );
  XNOR2_X1 Red_MCInst3_MC1_r2Inst_XORInst_0_0_U2  ( .A(
        Red_MCInst3_MC1_v3_2[0] ), .B(Red_MCInst3_MC1_v2_2[0] ), .ZN(
        Red_MCInst3_MC1_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 Red_MCInst3_MC1_r2Inst_XORInst_0_0_U1  ( .A(
        Red_MCInst3_MC1_v0_2[0] ), .B(Red_MCInst3_MC1_v1_2[0] ), .Z(
        Red_MCInst3_MC1_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 Red_MCInst3_MC1_r3Inst_XORInst_0_0_U3  ( .A(
        Red_MCInst3_MC1_r3Inst_XORInst_0_0_n5 ), .B(
        Red_MCInst3_MC1_r3Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback3[2]) );
  XNOR2_X1 Red_MCInst3_MC1_r3Inst_XORInst_0_0_U2  ( .A(
        Red_MCInst3_MC1_v3_3[0] ), .B(Red_MCInst3_MC1_v2_3[0] ), .ZN(
        Red_MCInst3_MC1_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 Red_MCInst3_MC1_r3Inst_XORInst_0_0_U1  ( .A(
        Red_MCInst3_MC1_v0_3[0] ), .B(Red_MCInst3_MC1_v1_3[0] ), .Z(
        Red_MCInst3_MC1_r3Inst_XORInst_0_0_n5 ) );
  XOR2_X1 Red_MCInst3_MC2_v0_0Inst_0_U3  ( .A(Red_MCInst3_MC2_v0_1[0] ), .B(
        MCInst3_MC2_v0_0 [3]), .Z(Red_MCInst3_MC2_v0_0[0] ) );
  XOR2_X1 Red_MCInst3_MC2_v0_2Inst_0_U3  ( .A(Red_MCInst3_MC2_v0_1[0] ), .B(
        MCInst3_MC2_v0_3 [0]), .Z(Red_MCInst3_MC2_v0_2[0] ) );
  XNOR2_X1 Red_MCInst3_MC2_v0_3Inst_0_U4  ( .A(
        Red_MCInst3_MC2_v0_3Inst_0_n2 ), .B(MCInst3_MC2_v0_0 [3]), .ZN(
        Red_MCInst3_MC2_v0_3[0] ) );
  XNOR2_X1 Red_MCInst3_MC2_v0_3Inst_0_U3  ( .A(MCInst3_MC2_v0_3 [3]), .B(
        Red_MCInst3_MC2_v0_1[0] ), .ZN(Red_MCInst3_MC2_v0_3Inst_0_n2 ) );
  XNOR2_X1 Red_MCInst3_MC2_v1_0Inst_0_U5  ( .A(
        Red_MCInst3_MC2_v1_0Inst_0_n4 ), .B(Red_MCInst3_MC2_v1_0Inst_0_n3 ), 
        .ZN(Red_MCInst3_MC2_v1_0[0] ) );
  XNOR2_X1 Red_MCInst3_MC2_v1_0Inst_0_U4  ( .A(MCInst3_MC2_v1_3 [2]), .B(
        MCInst3_MC2_v1_0 [0]), .ZN(Red_MCInst3_MC2_v1_0Inst_0_n3 ) );
  XOR2_X1 Red_MCInst3_MC2_v1_0Inst_0_U3  ( .A(Red_MCInst3_MC2_v1_1[0] ), .B(
        MCInst3_MC2_v1_0 [3]), .Z(Red_MCInst3_MC2_v1_0Inst_0_n4 ) );
  XOR2_X1 Red_MCInst3_MC2_v1_2Inst_0_U3  ( .A(MCInst3_MC2_v1_0 [0]), .B(
        Red_MCInst3_MC2_v1_1[0] ), .Z(Red_MCInst3_MC2_v1_2[0] ) );
  XNOR2_X1 Red_MCInst3_MC2_v1_3Inst_0_U4  ( .A(
        Red_MCInst3_MC2_v1_3Inst_0_n2 ), .B(MCInst3_MC2_v1_3 [2]), .ZN(
        Red_MCInst3_MC2_v1_3[0] ) );
  XNOR2_X1 Red_MCInst3_MC2_v1_3Inst_0_U3  ( .A(Red_MCInst3_MC2_v1_1[0] ), 
        .B(MCInst3_MC2_v1_0 [0]), .ZN(Red_MCInst3_MC2_v1_3Inst_0_n2 ) );
  XNOR2_X1 Red_MCInst3_MC2_v2_0Inst_0_U4  ( .A(
        Red_MCInst3_MC2_v2_0Inst_0_n2 ), .B(MCInst3_MC2_v2_0 [2]), .ZN(
        Red_MCInst3_MC2_v2_0[0] ) );
  XNOR2_X1 Red_MCInst3_MC2_v2_0Inst_0_U3  ( .A(MCInst3_MC2_v2_0 [3]), .B(
        MCInst3_MC2_v2_3 [1]), .ZN(Red_MCInst3_MC2_v2_0Inst_0_n2 ) );
  XOR2_X1 Red_MCInst3_MC2_v2_1Inst_0_U3  ( .A(MCInst3_MC2_v2_0 [3]), .B(
        MCInst3_MC2_v2_0 [0]), .Z(Red_MCInst3_MC2_v2_1[0] ) );
  XOR2_X1 Red_MCInst3_MC2_v2_2Inst_0_U3  ( .A(MCInst3_MC2_v2_0 [2]), .B(
        MCInst3_MC2_v2_0 [3]), .Z(Red_MCInst3_MC2_v2_2[0] ) );
  XOR2_X1 Red_MCInst3_MC2_v2_3Inst_0_U3  ( .A(MCInst3_MC2_v2_0 [2]), .B(
        MCInst3_MC2_v2_0 [0]), .Z(Red_MCInst3_MC2_v2_3[0] ) );
  XNOR2_X1 Red_MCInst3_MC2_v3_0Inst_0_U4  ( .A(
        Red_MCInst3_MC2_v3_0Inst_0_n2 ), .B(MCInst3_MC2_v3_0 [2]), .ZN(
        Red_MCInst3_MC2_v3_0[0] ) );
  XNOR2_X1 Red_MCInst3_MC2_v3_0Inst_0_U3  ( .A(Red_MCInst3_MC2_v3_1[0] ), 
        .B(MCInst3_MC2_v3_2 [3]), .ZN(Red_MCInst3_MC2_v3_0Inst_0_n2 ) );
  XNOR2_X1 Red_MCInst3_MC2_v3_2Inst_0_U4  ( .A(
        Red_MCInst3_MC2_v3_2Inst_0_n2 ), .B(Red_MCInst3_MC2_v3_1[0] ), .ZN(
        Red_MCInst3_MC2_v3_2[0] ) );
  XNOR2_X1 Red_MCInst3_MC2_v3_2Inst_0_U3  ( .A(MCInst3_MC2_v3_2 [2]), .B(
        MCInst3_MC2_v3_0 [2]), .ZN(Red_MCInst3_MC2_v3_2Inst_0_n2 ) );
  XOR2_X1 Red_MCInst3_MC2_v3_3Inst_0_U3  ( .A(MCInst3_MC2_v3_2 [3]), .B(
        MCInst3_MC2_v3_2 [2]), .Z(Red_MCInst3_MC2_v3_3[0] ) );
  XNOR2_X1 Red_MCInst3_MC2_r0Inst_XORInst_0_0_U3  ( .A(
        Red_MCInst3_MC2_r0Inst_XORInst_0_0_n5 ), .B(
        Red_MCInst3_MC2_r0Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback3[13]) );
  XNOR2_X1 Red_MCInst3_MC2_r0Inst_XORInst_0_0_U2  ( .A(
        Red_MCInst3_MC2_v3_0[0] ), .B(Red_MCInst3_MC2_v2_0[0] ), .ZN(
        Red_MCInst3_MC2_r0Inst_XORInst_0_0_n4 ) );
  XOR2_X1 Red_MCInst3_MC2_r0Inst_XORInst_0_0_U1  ( .A(
        Red_MCInst3_MC2_v0_0[0] ), .B(Red_MCInst3_MC2_v1_0[0] ), .Z(
        Red_MCInst3_MC2_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 Red_MCInst3_MC2_r1Inst_XORInst_0_0_U3  ( .A(
        Red_MCInst3_MC2_r1Inst_XORInst_0_0_n5 ), .B(
        Red_MCInst3_MC2_r1Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback3[9]) );
  XNOR2_X1 Red_MCInst3_MC2_r1Inst_XORInst_0_0_U2  ( .A(
        Red_MCInst3_MC2_v3_1[0] ), .B(Red_MCInst3_MC2_v2_1[0] ), .ZN(
        Red_MCInst3_MC2_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 Red_MCInst3_MC2_r1Inst_XORInst_0_0_U1  ( .A(
        Red_MCInst3_MC2_v0_1[0] ), .B(Red_MCInst3_MC2_v1_1[0] ), .Z(
        Red_MCInst3_MC2_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 Red_MCInst3_MC2_r2Inst_XORInst_0_0_U3  ( .A(
        Red_MCInst3_MC2_r2Inst_XORInst_0_0_n5 ), .B(
        Red_MCInst3_MC2_r2Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback3[5]) );
  XNOR2_X1 Red_MCInst3_MC2_r2Inst_XORInst_0_0_U2  ( .A(
        Red_MCInst3_MC2_v3_2[0] ), .B(Red_MCInst3_MC2_v2_2[0] ), .ZN(
        Red_MCInst3_MC2_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 Red_MCInst3_MC2_r2Inst_XORInst_0_0_U1  ( .A(
        Red_MCInst3_MC2_v0_2[0] ), .B(Red_MCInst3_MC2_v1_2[0] ), .Z(
        Red_MCInst3_MC2_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 Red_MCInst3_MC2_r3Inst_XORInst_0_0_U3  ( .A(
        Red_MCInst3_MC2_r3Inst_XORInst_0_0_n5 ), .B(
        Red_MCInst3_MC2_r3Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback3[1]) );
  XNOR2_X1 Red_MCInst3_MC2_r3Inst_XORInst_0_0_U2  ( .A(
        Red_MCInst3_MC2_v3_3[0] ), .B(Red_MCInst3_MC2_v2_3[0] ), .ZN(
        Red_MCInst3_MC2_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 Red_MCInst3_MC2_r3Inst_XORInst_0_0_U1  ( .A(
        Red_MCInst3_MC2_v0_3[0] ), .B(Red_MCInst3_MC2_v1_3[0] ), .Z(
        Red_MCInst3_MC2_r3Inst_XORInst_0_0_n5 ) );
  XOR2_X1 Red_MCInst3_MC3_v0_0Inst_0_U3  ( .A(Red_MCInst3_MC3_v0_1[0] ), .B(
        MCInst3_MC3_v0_0 [3]), .Z(Red_MCInst3_MC3_v0_0[0] ) );
  XOR2_X1 Red_MCInst3_MC3_v0_2Inst_0_U3  ( .A(Red_MCInst3_MC3_v0_1[0] ), .B(
        MCInst3_MC3_v0_3 [0]), .Z(Red_MCInst3_MC3_v0_2[0] ) );
  XNOR2_X1 Red_MCInst3_MC3_v0_3Inst_0_U4  ( .A(
        Red_MCInst3_MC3_v0_3Inst_0_n2 ), .B(MCInst3_MC3_v0_0 [3]), .ZN(
        Red_MCInst3_MC3_v0_3[0] ) );
  XNOR2_X1 Red_MCInst3_MC3_v0_3Inst_0_U3  ( .A(MCInst3_MC3_v0_3 [3]), .B(
        Red_MCInst3_MC3_v0_1[0] ), .ZN(Red_MCInst3_MC3_v0_3Inst_0_n2 ) );
  XNOR2_X1 Red_MCInst3_MC3_v1_0Inst_0_U5  ( .A(
        Red_MCInst3_MC3_v1_0Inst_0_n4 ), .B(Red_MCInst3_MC3_v1_0Inst_0_n3 ), 
        .ZN(Red_MCInst3_MC3_v1_0[0] ) );
  XNOR2_X1 Red_MCInst3_MC3_v1_0Inst_0_U4  ( .A(MCInst3_MC3_v1_3 [2]), .B(
        MCInst3_MC3_v1_0 [0]), .ZN(Red_MCInst3_MC3_v1_0Inst_0_n3 ) );
  XOR2_X1 Red_MCInst3_MC3_v1_0Inst_0_U3  ( .A(Red_MCInst3_MC3_v1_1[0] ), .B(
        MCInst3_MC3_v1_0 [3]), .Z(Red_MCInst3_MC3_v1_0Inst_0_n4 ) );
  XOR2_X1 Red_MCInst3_MC3_v1_2Inst_0_U3  ( .A(MCInst3_MC3_v1_0 [0]), .B(
        Red_MCInst3_MC3_v1_1[0] ), .Z(Red_MCInst3_MC3_v1_2[0] ) );
  XNOR2_X1 Red_MCInst3_MC3_v1_3Inst_0_U4  ( .A(
        Red_MCInst3_MC3_v1_3Inst_0_n2 ), .B(MCInst3_MC3_v1_3 [2]), .ZN(
        Red_MCInst3_MC3_v1_3[0] ) );
  XNOR2_X1 Red_MCInst3_MC3_v1_3Inst_0_U3  ( .A(Red_MCInst3_MC3_v1_1[0] ), 
        .B(MCInst3_MC3_v1_0 [0]), .ZN(Red_MCInst3_MC3_v1_3Inst_0_n2 ) );
  XNOR2_X1 Red_MCInst3_MC3_v2_0Inst_0_U4  ( .A(
        Red_MCInst3_MC3_v2_0Inst_0_n2 ), .B(MCInst3_MC3_v2_0 [2]), .ZN(
        Red_MCInst3_MC3_v2_0[0] ) );
  XNOR2_X1 Red_MCInst3_MC3_v2_0Inst_0_U3  ( .A(MCInst3_MC3_v2_0 [3]), .B(
        MCInst3_MC3_v2_3 [1]), .ZN(Red_MCInst3_MC3_v2_0Inst_0_n2 ) );
  XOR2_X1 Red_MCInst3_MC3_v2_1Inst_0_U3  ( .A(MCInst3_MC3_v2_0 [3]), .B(
        MCInst3_MC3_v2_0 [0]), .Z(Red_MCInst3_MC3_v2_1[0] ) );
  XOR2_X1 Red_MCInst3_MC3_v2_2Inst_0_U3  ( .A(MCInst3_MC3_v2_0 [2]), .B(
        MCInst3_MC3_v2_0 [3]), .Z(Red_MCInst3_MC3_v2_2[0] ) );
  XOR2_X1 Red_MCInst3_MC3_v2_3Inst_0_U3  ( .A(MCInst3_MC3_v2_0 [2]), .B(
        MCInst3_MC3_v2_0 [0]), .Z(Red_MCInst3_MC3_v2_3[0] ) );
  XNOR2_X1 Red_MCInst3_MC3_v3_0Inst_0_U4  ( .A(
        Red_MCInst3_MC3_v3_0Inst_0_n2 ), .B(MCInst3_MC3_v3_0 [2]), .ZN(
        Red_MCInst3_MC3_v3_0[0] ) );
  XNOR2_X1 Red_MCInst3_MC3_v3_0Inst_0_U3  ( .A(Red_MCInst3_MC3_v3_1[0] ), 
        .B(MCInst3_MC3_v3_2 [3]), .ZN(Red_MCInst3_MC3_v3_0Inst_0_n2 ) );
  XNOR2_X1 Red_MCInst3_MC3_v3_2Inst_0_U4  ( .A(
        Red_MCInst3_MC3_v3_2Inst_0_n2 ), .B(Red_MCInst3_MC3_v3_1[0] ), .ZN(
        Red_MCInst3_MC3_v3_2[0] ) );
  XNOR2_X1 Red_MCInst3_MC3_v3_2Inst_0_U3  ( .A(MCInst3_MC3_v3_2 [2]), .B(
        MCInst3_MC3_v3_0 [2]), .ZN(Red_MCInst3_MC3_v3_2Inst_0_n2 ) );
  XOR2_X1 Red_MCInst3_MC3_v3_3Inst_0_U3  ( .A(MCInst3_MC3_v3_2 [3]), .B(
        MCInst3_MC3_v3_2 [2]), .Z(Red_MCInst3_MC3_v3_3[0] ) );
  XNOR2_X1 Red_MCInst3_MC3_r0Inst_XORInst_0_0_U3  ( .A(
        Red_MCInst3_MC3_r0Inst_XORInst_0_0_n5 ), .B(
        Red_MCInst3_MC3_r0Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback3[12]) );
  XNOR2_X1 Red_MCInst3_MC3_r0Inst_XORInst_0_0_U2  ( .A(
        Red_MCInst3_MC3_v3_0[0] ), .B(Red_MCInst3_MC3_v2_0[0] ), .ZN(
        Red_MCInst3_MC3_r0Inst_XORInst_0_0_n4 ) );
  XOR2_X1 Red_MCInst3_MC3_r0Inst_XORInst_0_0_U1  ( .A(
        Red_MCInst3_MC3_v0_0[0] ), .B(Red_MCInst3_MC3_v1_0[0] ), .Z(
        Red_MCInst3_MC3_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 Red_MCInst3_MC3_r1Inst_XORInst_0_0_U3  ( .A(
        Red_MCInst3_MC3_r1Inst_XORInst_0_0_n5 ), .B(
        Red_MCInst3_MC3_r1Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback3[8]) );
  XNOR2_X1 Red_MCInst3_MC3_r1Inst_XORInst_0_0_U2  ( .A(
        Red_MCInst3_MC3_v3_1[0] ), .B(Red_MCInst3_MC3_v2_1[0] ), .ZN(
        Red_MCInst3_MC3_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 Red_MCInst3_MC3_r1Inst_XORInst_0_0_U1  ( .A(
        Red_MCInst3_MC3_v0_1[0] ), .B(Red_MCInst3_MC3_v1_1[0] ), .Z(
        Red_MCInst3_MC3_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 Red_MCInst3_MC3_r2Inst_XORInst_0_0_U3  ( .A(
        Red_MCInst3_MC3_r2Inst_XORInst_0_0_n5 ), .B(
        Red_MCInst3_MC3_r2Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback3[4]) );
  XNOR2_X1 Red_MCInst3_MC3_r2Inst_XORInst_0_0_U2  ( .A(
        Red_MCInst3_MC3_v3_2[0] ), .B(Red_MCInst3_MC3_v2_2[0] ), .ZN(
        Red_MCInst3_MC3_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 Red_MCInst3_MC3_r2Inst_XORInst_0_0_U1  ( .A(
        Red_MCInst3_MC3_v0_2[0] ), .B(Red_MCInst3_MC3_v1_2[0] ), .Z(
        Red_MCInst3_MC3_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 Red_MCInst3_MC3_r3Inst_XORInst_0_0_U3  ( .A(
        Red_MCInst3_MC3_r3Inst_XORInst_0_0_n5 ), .B(
        Red_MCInst3_MC3_r3Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback3[0]) );
  XNOR2_X1 Red_MCInst3_MC3_r3Inst_XORInst_0_0_U2  ( .A(
        Red_MCInst3_MC3_v3_3[0] ), .B(Red_MCInst3_MC3_v2_3[0] ), .ZN(
        Red_MCInst3_MC3_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 Red_MCInst3_MC3_r3Inst_XORInst_0_0_U1  ( .A(
        Red_MCInst3_MC3_v0_3[0] ), .B(Red_MCInst3_MC3_v1_3[0] ), .Z(
        Red_MCInst3_MC3_r3Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 Red_KeyInst_LFInst_0_LFInst_0_U5  ( .A(
        Red_KeyInst_LFInst_0_LFInst_0_n4 ), .B(
        Red_KeyInst_LFInst_0_LFInst_0_n3 ), .ZN(Red_RoundKey[0]) );
  XNOR2_X1 Red_KeyInst_LFInst_0_LFInst_0_U4  ( .A(Key[1]), .B(Key[0]), .ZN(
        Red_KeyInst_LFInst_0_LFInst_0_n3 ) );
  XOR2_X1 Red_KeyInst_LFInst_0_LFInst_0_U3  ( .A(Key[2]), .B(Key[3]), .Z(
        Red_KeyInst_LFInst_0_LFInst_0_n4 ) );
  XNOR2_X1 Red_KeyInst_LFInst_1_LFInst_0_U5  ( .A(
        Red_KeyInst_LFInst_1_LFInst_0_n4 ), .B(
        Red_KeyInst_LFInst_1_LFInst_0_n3 ), .ZN(Red_RoundKey[1]) );
  XNOR2_X1 Red_KeyInst_LFInst_1_LFInst_0_U4  ( .A(Key[5]), .B(Key[4]), .ZN(
        Red_KeyInst_LFInst_1_LFInst_0_n3 ) );
  XOR2_X1 Red_KeyInst_LFInst_1_LFInst_0_U3  ( .A(Key[6]), .B(Key[7]), .Z(
        Red_KeyInst_LFInst_1_LFInst_0_n4 ) );
  XNOR2_X1 Red_KeyInst_LFInst_2_LFInst_0_U5  ( .A(
        Red_KeyInst_LFInst_2_LFInst_0_n4 ), .B(
        Red_KeyInst_LFInst_2_LFInst_0_n3 ), .ZN(Red_RoundKey[2]) );
  XNOR2_X1 Red_KeyInst_LFInst_2_LFInst_0_U4  ( .A(Key[9]), .B(Key[8]), .ZN(
        Red_KeyInst_LFInst_2_LFInst_0_n3 ) );
  XOR2_X1 Red_KeyInst_LFInst_2_LFInst_0_U3  ( .A(Key[10]), .B(Key[11]), .Z(
        Red_KeyInst_LFInst_2_LFInst_0_n4 ) );
  XNOR2_X1 Red_KeyInst_LFInst_3_LFInst_0_U5  ( .A(
        Red_KeyInst_LFInst_3_LFInst_0_n4 ), .B(
        Red_KeyInst_LFInst_3_LFInst_0_n3 ), .ZN(Red_RoundKey[3]) );
  XNOR2_X1 Red_KeyInst_LFInst_3_LFInst_0_U4  ( .A(Key[13]), .B(Key[12]), .ZN(
        Red_KeyInst_LFInst_3_LFInst_0_n3 ) );
  XOR2_X1 Red_KeyInst_LFInst_3_LFInst_0_U3  ( .A(Key[14]), .B(Key[15]), .Z(
        Red_KeyInst_LFInst_3_LFInst_0_n4 ) );
  XNOR2_X1 Red_KeyInst_LFInst_4_LFInst_0_U5  ( .A(
        Red_KeyInst_LFInst_4_LFInst_0_n4 ), .B(
        Red_KeyInst_LFInst_4_LFInst_0_n3 ), .ZN(Red_RoundKey[4]) );
  XNOR2_X1 Red_KeyInst_LFInst_4_LFInst_0_U4  ( .A(Key[17]), .B(Key[16]), .ZN(
        Red_KeyInst_LFInst_4_LFInst_0_n3 ) );
  XOR2_X1 Red_KeyInst_LFInst_4_LFInst_0_U3  ( .A(Key[18]), .B(Key[19]), .Z(
        Red_KeyInst_LFInst_4_LFInst_0_n4 ) );
  XNOR2_X1 Red_KeyInst_LFInst_5_LFInst_0_U5  ( .A(
        Red_KeyInst_LFInst_5_LFInst_0_n4 ), .B(
        Red_KeyInst_LFInst_5_LFInst_0_n3 ), .ZN(Red_RoundKey[5]) );
  XNOR2_X1 Red_KeyInst_LFInst_5_LFInst_0_U4  ( .A(Key[21]), .B(Key[20]), .ZN(
        Red_KeyInst_LFInst_5_LFInst_0_n3 ) );
  XOR2_X1 Red_KeyInst_LFInst_5_LFInst_0_U3  ( .A(Key[22]), .B(Key[23]), .Z(
        Red_KeyInst_LFInst_5_LFInst_0_n4 ) );
  XNOR2_X1 Red_KeyInst_LFInst_6_LFInst_0_U5  ( .A(
        Red_KeyInst_LFInst_6_LFInst_0_n4 ), .B(
        Red_KeyInst_LFInst_6_LFInst_0_n3 ), .ZN(Red_RoundKey[6]) );
  XNOR2_X1 Red_KeyInst_LFInst_6_LFInst_0_U4  ( .A(Key[25]), .B(Key[24]), .ZN(
        Red_KeyInst_LFInst_6_LFInst_0_n3 ) );
  XOR2_X1 Red_KeyInst_LFInst_6_LFInst_0_U3  ( .A(Key[26]), .B(Key[27]), .Z(
        Red_KeyInst_LFInst_6_LFInst_0_n4 ) );
  XNOR2_X1 Red_KeyInst_LFInst_7_LFInst_0_U5  ( .A(
        Red_KeyInst_LFInst_7_LFInst_0_n4 ), .B(
        Red_KeyInst_LFInst_7_LFInst_0_n3 ), .ZN(Red_RoundKey[7]) );
  XNOR2_X1 Red_KeyInst_LFInst_7_LFInst_0_U4  ( .A(Key[29]), .B(Key[28]), .ZN(
        Red_KeyInst_LFInst_7_LFInst_0_n3 ) );
  XOR2_X1 Red_KeyInst_LFInst_7_LFInst_0_U3  ( .A(Key[30]), .B(Key[31]), .Z(
        Red_KeyInst_LFInst_7_LFInst_0_n4 ) );
  XNOR2_X1 Red_KeyInst_LFInst_8_LFInst_0_U5  ( .A(
        Red_KeyInst_LFInst_8_LFInst_0_n4 ), .B(
        Red_KeyInst_LFInst_8_LFInst_0_n3 ), .ZN(Red_RoundKey[8]) );
  XNOR2_X1 Red_KeyInst_LFInst_8_LFInst_0_U4  ( .A(Key[33]), .B(Key[32]), .ZN(
        Red_KeyInst_LFInst_8_LFInst_0_n3 ) );
  XOR2_X1 Red_KeyInst_LFInst_8_LFInst_0_U3  ( .A(Key[34]), .B(Key[35]), .Z(
        Red_KeyInst_LFInst_8_LFInst_0_n4 ) );
  XNOR2_X1 Red_KeyInst_LFInst_9_LFInst_0_U5  ( .A(
        Red_KeyInst_LFInst_9_LFInst_0_n4 ), .B(
        Red_KeyInst_LFInst_9_LFInst_0_n3 ), .ZN(Red_RoundKey[9]) );
  XNOR2_X1 Red_KeyInst_LFInst_9_LFInst_0_U4  ( .A(Key[37]), .B(Key[36]), .ZN(
        Red_KeyInst_LFInst_9_LFInst_0_n3 ) );
  XOR2_X1 Red_KeyInst_LFInst_9_LFInst_0_U3  ( .A(Key[38]), .B(Key[39]), .Z(
        Red_KeyInst_LFInst_9_LFInst_0_n4 ) );
  XNOR2_X1 Red_KeyInst_LFInst_10_LFInst_0_U5  ( .A(
        Red_KeyInst_LFInst_10_LFInst_0_n4 ), .B(
        Red_KeyInst_LFInst_10_LFInst_0_n3 ), .ZN(Red_RoundKey[10]) );
  XNOR2_X1 Red_KeyInst_LFInst_10_LFInst_0_U4  ( .A(Key[41]), .B(Key[40]), 
        .ZN(Red_KeyInst_LFInst_10_LFInst_0_n3 ) );
  XOR2_X1 Red_KeyInst_LFInst_10_LFInst_0_U3  ( .A(Key[42]), .B(Key[43]), .Z(
        Red_KeyInst_LFInst_10_LFInst_0_n4 ) );
  XNOR2_X1 Red_KeyInst_LFInst_11_LFInst_0_U5  ( .A(
        Red_KeyInst_LFInst_11_LFInst_0_n4 ), .B(
        Red_KeyInst_LFInst_11_LFInst_0_n3 ), .ZN(Red_RoundKey[11]) );
  XNOR2_X1 Red_KeyInst_LFInst_11_LFInst_0_U4  ( .A(Key[45]), .B(Key[44]), 
        .ZN(Red_KeyInst_LFInst_11_LFInst_0_n3 ) );
  XOR2_X1 Red_KeyInst_LFInst_11_LFInst_0_U3  ( .A(Key[46]), .B(Key[47]), .Z(
        Red_KeyInst_LFInst_11_LFInst_0_n4 ) );
  XNOR2_X1 Red_KeyInst_LFInst_12_LFInst_0_U5  ( .A(
        Red_KeyInst_LFInst_12_LFInst_0_n4 ), .B(
        Red_KeyInst_LFInst_12_LFInst_0_n3 ), .ZN(Red_RoundKey[12]) );
  XNOR2_X1 Red_KeyInst_LFInst_12_LFInst_0_U4  ( .A(Key[49]), .B(Key[48]), 
        .ZN(Red_KeyInst_LFInst_12_LFInst_0_n3 ) );
  XOR2_X1 Red_KeyInst_LFInst_12_LFInst_0_U3  ( .A(Key[50]), .B(Key[51]), .Z(
        Red_KeyInst_LFInst_12_LFInst_0_n4 ) );
  XNOR2_X1 Red_KeyInst_LFInst_13_LFInst_0_U5  ( .A(
        Red_KeyInst_LFInst_13_LFInst_0_n4 ), .B(
        Red_KeyInst_LFInst_13_LFInst_0_n3 ), .ZN(Red_RoundKey[13]) );
  XNOR2_X1 Red_KeyInst_LFInst_13_LFInst_0_U4  ( .A(Key[53]), .B(Key[52]), 
        .ZN(Red_KeyInst_LFInst_13_LFInst_0_n3 ) );
  XOR2_X1 Red_KeyInst_LFInst_13_LFInst_0_U3  ( .A(Key[54]), .B(Key[55]), .Z(
        Red_KeyInst_LFInst_13_LFInst_0_n4 ) );
  XNOR2_X1 Red_KeyInst_LFInst_14_LFInst_0_U5  ( .A(
        Red_KeyInst_LFInst_14_LFInst_0_n4 ), .B(
        Red_KeyInst_LFInst_14_LFInst_0_n3 ), .ZN(Red_RoundKey[14]) );
  XNOR2_X1 Red_KeyInst_LFInst_14_LFInst_0_U4  ( .A(Key[57]), .B(Key[56]), 
        .ZN(Red_KeyInst_LFInst_14_LFInst_0_n3 ) );
  XOR2_X1 Red_KeyInst_LFInst_14_LFInst_0_U3  ( .A(Key[58]), .B(Key[59]), .Z(
        Red_KeyInst_LFInst_14_LFInst_0_n4 ) );
  XNOR2_X1 Red_KeyInst_LFInst_15_LFInst_0_U5  ( .A(
        Red_KeyInst_LFInst_15_LFInst_0_n4 ), .B(
        Red_KeyInst_LFInst_15_LFInst_0_n3 ), .ZN(Red_RoundKey[15]) );
  XNOR2_X1 Red_KeyInst_LFInst_15_LFInst_0_U4  ( .A(Key[61]), .B(Key[60]), 
        .ZN(Red_KeyInst_LFInst_15_LFInst_0_n3 ) );
  XOR2_X1 Red_KeyInst_LFInst_15_LFInst_0_U3  ( .A(Key[62]), .B(Key[63]), .Z(
        Red_KeyInst_LFInst_15_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_0_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_0_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_0_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[0]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_0_LFInst_0_U4  ( .A(AddRoundKeyOutput[1]), 
        .B(AddRoundKeyOutput[0]), .ZN(Red_ToCheckInst_LFInst_0_LFInst_0_n3 )
         );
  XOR2_X1 Red_ToCheckInst_LFInst_0_LFInst_0_U3  ( .A(AddRoundKeyOutput[2]), 
        .B(AddRoundKeyOutput[3]), .Z(Red_ToCheckInst_LFInst_0_LFInst_0_n4 )
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_1_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_1_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_1_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[1]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_1_LFInst_0_U4  ( .A(AddRoundKeyOutput[5]), 
        .B(AddRoundKeyOutput[4]), .ZN(Red_ToCheckInst_LFInst_1_LFInst_0_n3 )
         );
  XOR2_X1 Red_ToCheckInst_LFInst_1_LFInst_0_U3  ( .A(AddRoundKeyOutput[6]), 
        .B(AddRoundKeyOutput[7]), .Z(Red_ToCheckInst_LFInst_1_LFInst_0_n4 )
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_2_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_2_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_2_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[2]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_2_LFInst_0_U4  ( .A(AddRoundKeyOutput[9]), 
        .B(AddRoundKeyOutput[8]), .ZN(Red_ToCheckInst_LFInst_2_LFInst_0_n3 )
         );
  XOR2_X1 Red_ToCheckInst_LFInst_2_LFInst_0_U3  ( .A(AddRoundKeyOutput[10]), 
        .B(AddRoundKeyOutput[11]), .Z(Red_ToCheckInst_LFInst_2_LFInst_0_n4 )
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_3_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_3_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_3_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[3]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_3_LFInst_0_U4  ( .A(AddRoundKeyOutput[13]), 
        .B(AddRoundKeyOutput[12]), .ZN(Red_ToCheckInst_LFInst_3_LFInst_0_n3 )
         );
  XOR2_X1 Red_ToCheckInst_LFInst_3_LFInst_0_U3  ( .A(AddRoundKeyOutput[14]), 
        .B(AddRoundKeyOutput[15]), .Z(Red_ToCheckInst_LFInst_3_LFInst_0_n4 )
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_4_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_4_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_4_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[4]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_4_LFInst_0_U4  ( .A(AddRoundKeyOutput[17]), 
        .B(AddRoundKeyOutput[16]), .ZN(Red_ToCheckInst_LFInst_4_LFInst_0_n3 )
         );
  XOR2_X1 Red_ToCheckInst_LFInst_4_LFInst_0_U3  ( .A(AddRoundKeyOutput[18]), 
        .B(AddRoundKeyOutput[19]), .Z(Red_ToCheckInst_LFInst_4_LFInst_0_n4 )
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_5_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_5_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_5_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[5]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_5_LFInst_0_U4  ( .A(AddRoundKeyOutput[21]), 
        .B(AddRoundKeyOutput[20]), .ZN(Red_ToCheckInst_LFInst_5_LFInst_0_n3 )
         );
  XOR2_X1 Red_ToCheckInst_LFInst_5_LFInst_0_U3  ( .A(AddRoundKeyOutput[22]), 
        .B(AddRoundKeyOutput[23]), .Z(Red_ToCheckInst_LFInst_5_LFInst_0_n4 )
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_6_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_6_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_6_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[6]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_6_LFInst_0_U4  ( .A(AddRoundKeyOutput[25]), 
        .B(AddRoundKeyOutput[24]), .ZN(Red_ToCheckInst_LFInst_6_LFInst_0_n3 )
         );
  XOR2_X1 Red_ToCheckInst_LFInst_6_LFInst_0_U3  ( .A(AddRoundKeyOutput[26]), 
        .B(AddRoundKeyOutput[27]), .Z(Red_ToCheckInst_LFInst_6_LFInst_0_n4 )
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_7_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_7_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_7_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[7]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_7_LFInst_0_U4  ( .A(AddRoundKeyOutput[29]), 
        .B(AddRoundKeyOutput[28]), .ZN(Red_ToCheckInst_LFInst_7_LFInst_0_n3 )
         );
  XOR2_X1 Red_ToCheckInst_LFInst_7_LFInst_0_U3  ( .A(AddRoundKeyOutput[30]), 
        .B(AddRoundKeyOutput[31]), .Z(Red_ToCheckInst_LFInst_7_LFInst_0_n4 )
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_8_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_8_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_8_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[8]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_8_LFInst_0_U4  ( .A(AddRoundKeyOutput[33]), 
        .B(AddRoundKeyOutput[32]), .ZN(Red_ToCheckInst_LFInst_8_LFInst_0_n3 )
         );
  XOR2_X1 Red_ToCheckInst_LFInst_8_LFInst_0_U3  ( .A(AddRoundKeyOutput[34]), 
        .B(AddRoundKeyOutput[35]), .Z(Red_ToCheckInst_LFInst_8_LFInst_0_n4 )
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_9_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_9_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_9_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[9]) );
  XNOR2_X1 Red_ToCheckInst_LFInst_9_LFInst_0_U4  ( .A(AddRoundKeyOutput[37]), 
        .B(AddRoundKeyOutput[36]), .ZN(Red_ToCheckInst_LFInst_9_LFInst_0_n3 )
         );
  XOR2_X1 Red_ToCheckInst_LFInst_9_LFInst_0_U3  ( .A(AddRoundKeyOutput[38]), 
        .B(AddRoundKeyOutput[39]), .Z(Red_ToCheckInst_LFInst_9_LFInst_0_n4 )
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_10_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_10_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_10_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[10])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_10_LFInst_0_U4  ( .A(AddRoundKeyOutput[41]), 
        .B(AddRoundKeyOutput[40]), .ZN(Red_ToCheckInst_LFInst_10_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_10_LFInst_0_U3  ( .A(AddRoundKeyOutput[42]), 
        .B(AddRoundKeyOutput[43]), .Z(Red_ToCheckInst_LFInst_10_LFInst_0_n4 )
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_11_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_11_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_11_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[11])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_11_LFInst_0_U4  ( .A(AddRoundKeyOutput[45]), 
        .B(AddRoundKeyOutput[44]), .ZN(Red_ToCheckInst_LFInst_11_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_11_LFInst_0_U3  ( .A(AddRoundKeyOutput[46]), 
        .B(AddRoundKeyOutput[47]), .Z(Red_ToCheckInst_LFInst_11_LFInst_0_n4 )
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_12_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_12_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_12_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[12])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_12_LFInst_0_U4  ( .A(AddRoundKeyOutput[49]), 
        .B(AddRoundKeyOutput[48]), .ZN(Red_ToCheckInst_LFInst_12_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_12_LFInst_0_U3  ( .A(AddRoundKeyOutput[50]), 
        .B(AddRoundKeyOutput[51]), .Z(Red_ToCheckInst_LFInst_12_LFInst_0_n4 )
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_13_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_13_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_13_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[13])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_13_LFInst_0_U4  ( .A(AddRoundKeyOutput[53]), 
        .B(AddRoundKeyOutput[52]), .ZN(Red_ToCheckInst_LFInst_13_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_13_LFInst_0_U3  ( .A(AddRoundKeyOutput[54]), 
        .B(AddRoundKeyOutput[55]), .Z(Red_ToCheckInst_LFInst_13_LFInst_0_n4 )
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_14_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_14_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_14_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[14])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_14_LFInst_0_U4  ( .A(AddRoundKeyOutput[57]), 
        .B(AddRoundKeyOutput[56]), .ZN(Red_ToCheckInst_LFInst_14_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_14_LFInst_0_U3  ( .A(AddRoundKeyOutput[58]), 
        .B(AddRoundKeyOutput[59]), .Z(Red_ToCheckInst_LFInst_14_LFInst_0_n4 )
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_15_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_15_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_15_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[15])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_15_LFInst_0_U4  ( .A(AddRoundKeyOutput[61]), 
        .B(AddRoundKeyOutput[60]), .ZN(Red_ToCheckInst_LFInst_15_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_15_LFInst_0_U3  ( .A(AddRoundKeyOutput[62]), 
        .B(AddRoundKeyOutput[63]), .Z(Red_ToCheckInst_LFInst_15_LFInst_0_n4 )
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_16_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_16_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_16_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[16])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_16_LFInst_0_U4  ( .A(Ciphertext[1]), .B(
        Ciphertext[0]), .ZN(Red_ToCheckInst_LFInst_16_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_16_LFInst_0_U3  ( .A(Ciphertext[2]), .B(
        Ciphertext[3]), .Z(Red_ToCheckInst_LFInst_16_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_17_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_17_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_17_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[17])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_17_LFInst_0_U4  ( .A(Ciphertext[5]), .B(
        Ciphertext[4]), .ZN(Red_ToCheckInst_LFInst_17_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_17_LFInst_0_U3  ( .A(Ciphertext[6]), .B(
        Ciphertext[7]), .Z(Red_ToCheckInst_LFInst_17_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_18_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_18_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_18_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[18])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_18_LFInst_0_U4  ( .A(Ciphertext[9]), .B(
        Ciphertext[8]), .ZN(Red_ToCheckInst_LFInst_18_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_18_LFInst_0_U3  ( .A(Ciphertext[10]), .B(
        Ciphertext[11]), .Z(Red_ToCheckInst_LFInst_18_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_19_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_19_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_19_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[19])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_19_LFInst_0_U4  ( .A(Ciphertext[13]), .B(
        Ciphertext[12]), .ZN(Red_ToCheckInst_LFInst_19_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_19_LFInst_0_U3  ( .A(Ciphertext[14]), .B(
        Ciphertext[15]), .Z(Red_ToCheckInst_LFInst_19_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_20_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_20_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_20_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[20])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_20_LFInst_0_U4  ( .A(Ciphertext[17]), .B(
        Ciphertext[16]), .ZN(Red_ToCheckInst_LFInst_20_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_20_LFInst_0_U3  ( .A(Ciphertext[18]), .B(
        Ciphertext[19]), .Z(Red_ToCheckInst_LFInst_20_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_21_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_21_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_21_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[21])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_21_LFInst_0_U4  ( .A(Ciphertext[21]), .B(
        Ciphertext[20]), .ZN(Red_ToCheckInst_LFInst_21_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_21_LFInst_0_U3  ( .A(Ciphertext[22]), .B(
        Ciphertext[23]), .Z(Red_ToCheckInst_LFInst_21_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_22_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_22_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_22_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[22])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_22_LFInst_0_U4  ( .A(Ciphertext[25]), .B(
        Ciphertext[24]), .ZN(Red_ToCheckInst_LFInst_22_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_22_LFInst_0_U3  ( .A(Ciphertext[26]), .B(
        Ciphertext[27]), .Z(Red_ToCheckInst_LFInst_22_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_23_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_23_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_23_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[23])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_23_LFInst_0_U4  ( .A(Ciphertext[29]), .B(
        Ciphertext[28]), .ZN(Red_ToCheckInst_LFInst_23_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_23_LFInst_0_U3  ( .A(Ciphertext[30]), .B(
        Ciphertext[31]), .Z(Red_ToCheckInst_LFInst_23_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_24_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_24_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_24_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[24])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_24_LFInst_0_U4  ( .A(Ciphertext[33]), .B(
        Ciphertext[32]), .ZN(Red_ToCheckInst_LFInst_24_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_24_LFInst_0_U3  ( .A(Ciphertext[34]), .B(
        Ciphertext[35]), .Z(Red_ToCheckInst_LFInst_24_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_25_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_25_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_25_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[25])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_25_LFInst_0_U4  ( .A(Ciphertext[37]), .B(
        Ciphertext[36]), .ZN(Red_ToCheckInst_LFInst_25_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_25_LFInst_0_U3  ( .A(Ciphertext[38]), .B(
        Ciphertext[39]), .Z(Red_ToCheckInst_LFInst_25_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_26_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_26_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_26_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[26])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_26_LFInst_0_U4  ( .A(Ciphertext[41]), .B(
        Ciphertext[40]), .ZN(Red_ToCheckInst_LFInst_26_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_26_LFInst_0_U3  ( .A(Ciphertext[42]), .B(
        Ciphertext[43]), .Z(Red_ToCheckInst_LFInst_26_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_27_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_27_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_27_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[27])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_27_LFInst_0_U4  ( .A(Ciphertext[45]), .B(
        Ciphertext[44]), .ZN(Red_ToCheckInst_LFInst_27_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_27_LFInst_0_U3  ( .A(Ciphertext[46]), .B(
        Ciphertext[47]), .Z(Red_ToCheckInst_LFInst_27_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_28_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_28_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_28_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[28])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_28_LFInst_0_U4  ( .A(Ciphertext[49]), .B(
        Ciphertext[48]), .ZN(Red_ToCheckInst_LFInst_28_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_28_LFInst_0_U3  ( .A(Ciphertext[50]), .B(
        Ciphertext[51]), .Z(Red_ToCheckInst_LFInst_28_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_29_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_29_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_29_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[29])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_29_LFInst_0_U4  ( .A(Ciphertext[53]), .B(
        Ciphertext[52]), .ZN(Red_ToCheckInst_LFInst_29_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_29_LFInst_0_U3  ( .A(Ciphertext[54]), .B(
        Ciphertext[55]), .Z(Red_ToCheckInst_LFInst_29_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_30_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_30_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_30_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[30])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_30_LFInst_0_U4  ( .A(Ciphertext[57]), .B(
        Ciphertext[56]), .ZN(Red_ToCheckInst_LFInst_30_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_30_LFInst_0_U3  ( .A(Ciphertext[58]), .B(
        Ciphertext[59]), .Z(Red_ToCheckInst_LFInst_30_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_31_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_31_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_31_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[31])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_31_LFInst_0_U4  ( .A(Ciphertext[61]), .B(
        Ciphertext[60]), .ZN(Red_ToCheckInst_LFInst_31_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_31_LFInst_0_U3  ( .A(Ciphertext[62]), .B(
        Ciphertext[63]), .Z(Red_ToCheckInst_LFInst_31_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_32_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_32_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_32_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[32])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_32_LFInst_0_U4  ( .A(MCInst3_MC3_v3_0 [2]), 
        .B(MCInst3_MC3_v3_2 [3]), .ZN(Red_ToCheckInst_LFInst_32_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_32_LFInst_0_U3  ( .A(
        Red_MCInst3_MC3_v3_1[0] ), .B(MCInst3_MC3_v3_2 [2]), .Z(
        Red_ToCheckInst_LFInst_32_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_33_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_33_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_33_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[33])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_33_LFInst_0_U4  ( .A(MCInst3_MC2_v3_0 [2]), 
        .B(MCInst3_MC2_v3_2 [3]), .ZN(Red_ToCheckInst_LFInst_33_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_33_LFInst_0_U3  ( .A(
        Red_MCInst3_MC2_v3_1[0] ), .B(MCInst3_MC2_v3_2 [2]), .Z(
        Red_ToCheckInst_LFInst_33_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_34_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_34_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_34_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[34])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_34_LFInst_0_U4  ( .A(MCInst3_MC1_v3_0 [2]), 
        .B(MCInst3_MC1_v3_2 [3]), .ZN(Red_ToCheckInst_LFInst_34_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_34_LFInst_0_U3  ( .A(
        Red_MCInst3_MC1_v3_1[0] ), .B(MCInst3_MC1_v3_2 [2]), .Z(
        Red_ToCheckInst_LFInst_34_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_35_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_35_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_35_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[35])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_35_LFInst_0_U4  ( .A(MCInst3_MC0_v3_0 [2]), 
        .B(MCInst3_MC0_v3_2 [3]), .ZN(Red_ToCheckInst_LFInst_35_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_35_LFInst_0_U3  ( .A(
        Red_MCInst3_MC0_v3_1[0] ), .B(MCInst3_MC0_v3_2 [2]), .Z(
        Red_ToCheckInst_LFInst_35_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_36_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_36_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_36_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[36])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_36_LFInst_0_U4  ( .A(MCInst3_MC3_v2_0 [2]), 
        .B(MCInst3_MC3_v2_3 [1]), .ZN(Red_ToCheckInst_LFInst_36_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_36_LFInst_0_U3  ( .A(MCInst3_MC3_v2_0 [3]), 
        .B(MCInst3_MC3_v2_0 [0]), .Z(Red_ToCheckInst_LFInst_36_LFInst_0_n4 )
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_37_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_37_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_37_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[37])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_37_LFInst_0_U4  ( .A(MCInst3_MC2_v2_0 [2]), 
        .B(MCInst3_MC2_v2_3 [1]), .ZN(Red_ToCheckInst_LFInst_37_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_37_LFInst_0_U3  ( .A(MCInst3_MC2_v2_0 [3]), 
        .B(MCInst3_MC2_v2_0 [0]), .Z(Red_ToCheckInst_LFInst_37_LFInst_0_n4 )
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_38_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_38_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_38_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[38])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_38_LFInst_0_U4  ( .A(MCInst3_MC1_v2_0 [2]), 
        .B(MCInst3_MC1_v2_3 [1]), .ZN(Red_ToCheckInst_LFInst_38_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_38_LFInst_0_U3  ( .A(MCInst3_MC1_v2_0 [3]), 
        .B(MCInst3_MC1_v2_0 [0]), .Z(Red_ToCheckInst_LFInst_38_LFInst_0_n4 )
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_39_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_39_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_39_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[39])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_39_LFInst_0_U4  ( .A(MCInst3_MC0_v2_0 [2]), 
        .B(MCInst3_MC0_v2_3 [1]), .ZN(Red_ToCheckInst_LFInst_39_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_39_LFInst_0_U3  ( .A(MCInst3_MC0_v2_0 [3]), 
        .B(MCInst3_MC0_v2_0 [0]), .Z(Red_ToCheckInst_LFInst_39_LFInst_0_n4 )
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_40_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_40_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_40_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[40])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_40_LFInst_0_U4  ( .A(MCInst3_MC3_v1_3 [2]), 
        .B(MCInst3_MC3_v1_0 [0]), .ZN(Red_ToCheckInst_LFInst_40_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_40_LFInst_0_U3  ( .A(
        Red_MCInst3_MC3_v1_1[0] ), .B(MCInst3_MC3_v1_0 [3]), .Z(
        Red_ToCheckInst_LFInst_40_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_41_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_41_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_41_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[41])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_41_LFInst_0_U4  ( .A(MCInst3_MC2_v1_3 [2]), 
        .B(MCInst3_MC2_v1_0 [0]), .ZN(Red_ToCheckInst_LFInst_41_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_41_LFInst_0_U3  ( .A(
        Red_MCInst3_MC2_v1_1[0] ), .B(MCInst3_MC2_v1_0 [3]), .Z(
        Red_ToCheckInst_LFInst_41_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_42_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_42_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_42_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[42])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_42_LFInst_0_U4  ( .A(MCInst3_MC1_v1_3 [2]), 
        .B(MCInst3_MC1_v1_0 [0]), .ZN(Red_ToCheckInst_LFInst_42_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_42_LFInst_0_U3  ( .A(
        Red_MCInst3_MC1_v1_1[0] ), .B(MCInst3_MC1_v1_0 [3]), .Z(
        Red_ToCheckInst_LFInst_42_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_43_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_43_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_43_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[43])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_43_LFInst_0_U4  ( .A(MCInst3_MC0_v1_3 [2]), 
        .B(MCInst3_MC0_v1_0 [0]), .ZN(Red_ToCheckInst_LFInst_43_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_43_LFInst_0_U3  ( .A(
        Red_MCInst3_MC0_v1_1[0] ), .B(MCInst3_MC0_v1_0 [3]), .Z(
        Red_ToCheckInst_LFInst_43_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_44_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_44_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_44_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[44])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_44_LFInst_0_U4  ( .A(MCInst3_MC3_v0_0 [3]), 
        .B(Red_MCInst3_MC3_v0_1[0] ), .ZN(
        Red_ToCheckInst_LFInst_44_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_44_LFInst_0_U3  ( .A(MCInst3_MC3_v0_3 [3]), 
        .B(MCInst3_MC3_v0_3 [0]), .Z(Red_ToCheckInst_LFInst_44_LFInst_0_n4 )
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_45_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_45_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_45_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[45])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_45_LFInst_0_U4  ( .A(MCInst3_MC2_v0_0 [3]), 
        .B(Red_MCInst3_MC2_v0_1[0] ), .ZN(
        Red_ToCheckInst_LFInst_45_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_45_LFInst_0_U3  ( .A(MCInst3_MC2_v0_3 [3]), 
        .B(MCInst3_MC2_v0_3 [0]), .Z(Red_ToCheckInst_LFInst_45_LFInst_0_n4 )
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_46_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_46_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_46_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[46])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_46_LFInst_0_U4  ( .A(MCInst3_MC1_v0_0 [3]), 
        .B(Red_MCInst3_MC1_v0_1[0] ), .ZN(
        Red_ToCheckInst_LFInst_46_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_46_LFInst_0_U3  ( .A(MCInst3_MC1_v0_3 [3]), 
        .B(MCInst3_MC1_v0_3 [0]), .Z(Red_ToCheckInst_LFInst_46_LFInst_0_n4 )
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_47_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_47_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_47_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[47])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_47_LFInst_0_U4  ( .A(MCInst3_MC0_v0_0 [3]), 
        .B(Red_MCInst3_MC0_v0_1[0] ), .ZN(
        Red_ToCheckInst_LFInst_47_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_47_LFInst_0_U3  ( .A(MCInst3_MC0_v0_3 [3]), 
        .B(MCInst3_MC0_v0_3 [0]), .Z(Red_ToCheckInst_LFInst_47_LFInst_0_n4 )
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_48_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_48_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_48_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[48])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_48_LFInst_0_U4  ( .A(SubCellInput2[1]), .B(
        SubCellInput2[0]), .ZN(Red_ToCheckInst_LFInst_48_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_48_LFInst_0_U3  ( .A(SubCellInput2[2]), .B(
        SubCellInput2[3]), .Z(Red_ToCheckInst_LFInst_48_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_49_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_49_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_49_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[49])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_49_LFInst_0_U4  ( .A(SubCellInput2[5]), .B(
        SubCellInput2[4]), .ZN(Red_ToCheckInst_LFInst_49_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_49_LFInst_0_U3  ( .A(SubCellInput2[6]), .B(
        SubCellInput2[7]), .Z(Red_ToCheckInst_LFInst_49_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_50_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_50_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_50_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[50])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_50_LFInst_0_U4  ( .A(SubCellInput2[9]), .B(
        SubCellInput2[8]), .ZN(Red_ToCheckInst_LFInst_50_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_50_LFInst_0_U3  ( .A(SubCellInput2[10]), .B(
        SubCellInput2[11]), .Z(Red_ToCheckInst_LFInst_50_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_51_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_51_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_51_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[51])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_51_LFInst_0_U4  ( .A(SubCellInput2[13]), 
        .B(SubCellInput2[12]), .ZN(Red_ToCheckInst_LFInst_51_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_51_LFInst_0_U3  ( .A(SubCellInput2[14]), .B(
        SubCellInput2[15]), .Z(Red_ToCheckInst_LFInst_51_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_52_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_52_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_52_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[52])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_52_LFInst_0_U4  ( .A(SubCellInput2[17]), 
        .B(SubCellInput2[16]), .ZN(Red_ToCheckInst_LFInst_52_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_52_LFInst_0_U3  ( .A(SubCellInput2[18]), .B(
        SubCellInput2[19]), .Z(Red_ToCheckInst_LFInst_52_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_53_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_53_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_53_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[53])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_53_LFInst_0_U4  ( .A(SubCellInput2[21]), 
        .B(SubCellInput2[20]), .ZN(Red_ToCheckInst_LFInst_53_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_53_LFInst_0_U3  ( .A(SubCellInput2[22]), .B(
        SubCellInput2[23]), .Z(Red_ToCheckInst_LFInst_53_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_54_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_54_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_54_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[54])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_54_LFInst_0_U4  ( .A(SubCellInput2[25]), 
        .B(SubCellInput2[24]), .ZN(Red_ToCheckInst_LFInst_54_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_54_LFInst_0_U3  ( .A(SubCellInput2[26]), .B(
        SubCellInput2[27]), .Z(Red_ToCheckInst_LFInst_54_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_55_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_55_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_55_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[55])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_55_LFInst_0_U4  ( .A(SubCellInput2[29]), 
        .B(SubCellInput2[28]), .ZN(Red_ToCheckInst_LFInst_55_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_55_LFInst_0_U3  ( .A(SubCellInput2[30]), .B(
        SubCellInput2[31]), .Z(Red_ToCheckInst_LFInst_55_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_56_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_56_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_56_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[56])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_56_LFInst_0_U4  ( .A(SubCellInput2[33]), 
        .B(SubCellInput2[32]), .ZN(Red_ToCheckInst_LFInst_56_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_56_LFInst_0_U3  ( .A(SubCellInput2[34]), .B(
        SubCellInput2[35]), .Z(Red_ToCheckInst_LFInst_56_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_57_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_57_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_57_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[57])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_57_LFInst_0_U4  ( .A(SubCellInput2[37]), 
        .B(SubCellInput2[36]), .ZN(Red_ToCheckInst_LFInst_57_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_57_LFInst_0_U3  ( .A(SubCellInput2[38]), .B(
        SubCellInput2[39]), .Z(Red_ToCheckInst_LFInst_57_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_58_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_58_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_58_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[58])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_58_LFInst_0_U4  ( .A(SubCellInput2[41]), 
        .B(SubCellInput2[40]), .ZN(Red_ToCheckInst_LFInst_58_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_58_LFInst_0_U3  ( .A(SubCellInput2[42]), .B(
        SubCellInput2[43]), .Z(Red_ToCheckInst_LFInst_58_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_59_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_59_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_59_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[59])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_59_LFInst_0_U4  ( .A(SubCellInput2[45]), 
        .B(SubCellInput2[44]), .ZN(Red_ToCheckInst_LFInst_59_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_59_LFInst_0_U3  ( .A(SubCellInput2[46]), .B(
        SubCellInput2[47]), .Z(Red_ToCheckInst_LFInst_59_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_60_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_60_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_60_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[60])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_60_LFInst_0_U4  ( .A(SubCellInput2[49]), 
        .B(SubCellInput2[48]), .ZN(Red_ToCheckInst_LFInst_60_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_60_LFInst_0_U3  ( .A(SubCellInput2[50]), .B(
        SubCellInput2[51]), .Z(Red_ToCheckInst_LFInst_60_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_61_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_61_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_61_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[61])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_61_LFInst_0_U4  ( .A(SubCellInput2[53]), 
        .B(SubCellInput2[52]), .ZN(Red_ToCheckInst_LFInst_61_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_61_LFInst_0_U3  ( .A(SubCellInput2[54]), .B(
        SubCellInput2[55]), .Z(Red_ToCheckInst_LFInst_61_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_62_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_62_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_62_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[62])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_62_LFInst_0_U4  ( .A(SubCellInput2[57]), 
        .B(SubCellInput2[56]), .ZN(Red_ToCheckInst_LFInst_62_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_62_LFInst_0_U3  ( .A(SubCellInput2[58]), .B(
        SubCellInput2[59]), .Z(Red_ToCheckInst_LFInst_62_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_63_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_63_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_63_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[63])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_63_LFInst_0_U4  ( .A(SubCellInput2[61]), 
        .B(SubCellInput2[60]), .ZN(Red_ToCheckInst_LFInst_63_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_63_LFInst_0_U3  ( .A(SubCellInput2[62]), .B(
        SubCellInput2[63]), .Z(Red_ToCheckInst_LFInst_63_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_64_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_64_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_64_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[64])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_64_LFInst_0_U4  ( .A(Feedback2[1]), .B(
        Feedback2[0]), .ZN(Red_ToCheckInst_LFInst_64_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_64_LFInst_0_U3  ( .A(Feedback2[2]), .B(
        Feedback2[3]), .Z(Red_ToCheckInst_LFInst_64_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_65_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_65_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_65_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[65])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_65_LFInst_0_U4  ( .A(Feedback2[5]), .B(
        Feedback2[4]), .ZN(Red_ToCheckInst_LFInst_65_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_65_LFInst_0_U3  ( .A(Feedback2[6]), .B(
        Feedback2[7]), .Z(Red_ToCheckInst_LFInst_65_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_66_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_66_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_66_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[66])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_66_LFInst_0_U4  ( .A(Feedback2[9]), .B(
        Feedback2[8]), .ZN(Red_ToCheckInst_LFInst_66_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_66_LFInst_0_U3  ( .A(Feedback2[10]), .B(
        Feedback2[11]), .Z(Red_ToCheckInst_LFInst_66_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_67_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_67_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_67_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[67])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_67_LFInst_0_U4  ( .A(Feedback2[13]), .B(
        Feedback2[12]), .ZN(Red_ToCheckInst_LFInst_67_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_67_LFInst_0_U3  ( .A(Feedback2[14]), .B(
        Feedback2[15]), .Z(Red_ToCheckInst_LFInst_67_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_68_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_68_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_68_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[68])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_68_LFInst_0_U4  ( .A(Feedback2[17]), .B(
        Feedback2[16]), .ZN(Red_ToCheckInst_LFInst_68_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_68_LFInst_0_U3  ( .A(Feedback2[18]), .B(
        Feedback2[19]), .Z(Red_ToCheckInst_LFInst_68_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_69_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_69_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_69_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[69])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_69_LFInst_0_U4  ( .A(Feedback2[21]), .B(
        Feedback2[20]), .ZN(Red_ToCheckInst_LFInst_69_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_69_LFInst_0_U3  ( .A(Feedback2[22]), .B(
        Feedback2[23]), .Z(Red_ToCheckInst_LFInst_69_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_70_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_70_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_70_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[70])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_70_LFInst_0_U4  ( .A(Feedback2[25]), .B(
        Feedback2[24]), .ZN(Red_ToCheckInst_LFInst_70_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_70_LFInst_0_U3  ( .A(Feedback2[26]), .B(
        Feedback2[27]), .Z(Red_ToCheckInst_LFInst_70_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_71_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_71_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_71_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[71])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_71_LFInst_0_U4  ( .A(Feedback2[29]), .B(
        Feedback2[28]), .ZN(Red_ToCheckInst_LFInst_71_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_71_LFInst_0_U3  ( .A(Feedback2[30]), .B(
        Feedback2[31]), .Z(Red_ToCheckInst_LFInst_71_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_72_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_72_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_72_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[72])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_72_LFInst_0_U4  ( .A(Feedback2[33]), .B(
        Feedback2[32]), .ZN(Red_ToCheckInst_LFInst_72_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_72_LFInst_0_U3  ( .A(Feedback2[34]), .B(
        Feedback2[35]), .Z(Red_ToCheckInst_LFInst_72_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_73_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_73_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_73_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[73])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_73_LFInst_0_U4  ( .A(Feedback2[37]), .B(
        Feedback2[36]), .ZN(Red_ToCheckInst_LFInst_73_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_73_LFInst_0_U3  ( .A(Feedback2[38]), .B(
        Feedback2[39]), .Z(Red_ToCheckInst_LFInst_73_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_74_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_74_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_74_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[74])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_74_LFInst_0_U4  ( .A(Feedback2[41]), .B(
        Feedback2[40]), .ZN(Red_ToCheckInst_LFInst_74_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_74_LFInst_0_U3  ( .A(Feedback2[42]), .B(
        Feedback2[43]), .Z(Red_ToCheckInst_LFInst_74_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_75_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_75_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_75_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[75])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_75_LFInst_0_U4  ( .A(Feedback2[45]), .B(
        Feedback2[44]), .ZN(Red_ToCheckInst_LFInst_75_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_75_LFInst_0_U3  ( .A(Feedback2[46]), .B(
        Feedback2[47]), .Z(Red_ToCheckInst_LFInst_75_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_76_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_76_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_76_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[76])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_76_LFInst_0_U4  ( .A(Feedback2[49]), .B(
        Feedback2[48]), .ZN(Red_ToCheckInst_LFInst_76_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_76_LFInst_0_U3  ( .A(Feedback2[50]), .B(
        Feedback2[51]), .Z(Red_ToCheckInst_LFInst_76_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_77_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_77_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_77_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[77])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_77_LFInst_0_U4  ( .A(Feedback2[53]), .B(
        Feedback2[52]), .ZN(Red_ToCheckInst_LFInst_77_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_77_LFInst_0_U3  ( .A(Feedback2[54]), .B(
        Feedback2[55]), .Z(Red_ToCheckInst_LFInst_77_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_78_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_78_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_78_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[78])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_78_LFInst_0_U4  ( .A(Feedback2[57]), .B(
        Feedback2[56]), .ZN(Red_ToCheckInst_LFInst_78_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_78_LFInst_0_U3  ( .A(Feedback2[58]), .B(
        Feedback2[59]), .Z(Red_ToCheckInst_LFInst_78_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_79_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_79_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_79_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[79])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_79_LFInst_0_U4  ( .A(Feedback2[61]), .B(
        Feedback2[60]), .ZN(Red_ToCheckInst_LFInst_79_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_79_LFInst_0_U3  ( .A(Feedback2[62]), .B(
        Feedback2[63]), .Z(Red_ToCheckInst_LFInst_79_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_80_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_80_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_80_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[80])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_80_LFInst_0_U4  ( .A(MCInst2_MC3_v3_0 [2]), 
        .B(MCInst2_MC3_v3_2 [3]), .ZN(Red_ToCheckInst_LFInst_80_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_80_LFInst_0_U3  ( .A(
        Red_MCInst2_MC3_v3_1[0] ), .B(MCInst2_MC3_v3_2 [2]), .Z(
        Red_ToCheckInst_LFInst_80_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_81_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_81_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_81_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[81])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_81_LFInst_0_U4  ( .A(MCInst2_MC2_v3_0 [2]), 
        .B(MCInst2_MC2_v3_2 [3]), .ZN(Red_ToCheckInst_LFInst_81_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_81_LFInst_0_U3  ( .A(
        Red_MCInst2_MC2_v3_1[0] ), .B(MCInst2_MC2_v3_2 [2]), .Z(
        Red_ToCheckInst_LFInst_81_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_82_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_82_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_82_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[82])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_82_LFInst_0_U4  ( .A(MCInst2_MC1_v3_0 [2]), 
        .B(MCInst2_MC1_v3_2 [3]), .ZN(Red_ToCheckInst_LFInst_82_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_82_LFInst_0_U3  ( .A(
        Red_MCInst2_MC1_v3_1[0] ), .B(MCInst2_MC1_v3_2 [2]), .Z(
        Red_ToCheckInst_LFInst_82_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_83_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_83_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_83_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[83])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_83_LFInst_0_U4  ( .A(MCInst2_MC0_v3_0 [2]), 
        .B(MCInst2_MC0_v3_2 [3]), .ZN(Red_ToCheckInst_LFInst_83_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_83_LFInst_0_U3  ( .A(
        Red_MCInst2_MC0_v3_1[0] ), .B(MCInst2_MC0_v3_2 [2]), .Z(
        Red_ToCheckInst_LFInst_83_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_84_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_84_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_84_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[84])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_84_LFInst_0_U4  ( .A(MCInst2_MC3_v2_0 [2]), 
        .B(MCInst2_MC3_v2_3 [1]), .ZN(Red_ToCheckInst_LFInst_84_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_84_LFInst_0_U3  ( .A(MCInst2_MC3_v2_0 [3]), 
        .B(MCInst2_MC3_v2_0 [0]), .Z(Red_ToCheckInst_LFInst_84_LFInst_0_n4 )
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_85_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_85_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_85_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[85])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_85_LFInst_0_U4  ( .A(MCInst2_MC2_v2_0 [2]), 
        .B(MCInst2_MC2_v2_3 [1]), .ZN(Red_ToCheckInst_LFInst_85_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_85_LFInst_0_U3  ( .A(MCInst2_MC2_v2_0 [3]), 
        .B(MCInst2_MC2_v2_0 [0]), .Z(Red_ToCheckInst_LFInst_85_LFInst_0_n4 )
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_86_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_86_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_86_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[86])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_86_LFInst_0_U4  ( .A(MCInst2_MC1_v2_0 [2]), 
        .B(MCInst2_MC1_v2_3 [1]), .ZN(Red_ToCheckInst_LFInst_86_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_86_LFInst_0_U3  ( .A(MCInst2_MC1_v2_0 [3]), 
        .B(MCInst2_MC1_v2_0 [0]), .Z(Red_ToCheckInst_LFInst_86_LFInst_0_n4 )
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_87_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_87_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_87_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[87])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_87_LFInst_0_U4  ( .A(MCInst2_MC0_v2_0 [2]), 
        .B(MCInst2_MC0_v2_3 [1]), .ZN(Red_ToCheckInst_LFInst_87_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_87_LFInst_0_U3  ( .A(MCInst2_MC0_v2_0 [3]), 
        .B(MCInst2_MC0_v2_0 [0]), .Z(Red_ToCheckInst_LFInst_87_LFInst_0_n4 )
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_88_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_88_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_88_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[88])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_88_LFInst_0_U4  ( .A(MCInst2_MC3_v1_3 [2]), 
        .B(MCInst2_MC3_v1_0 [0]), .ZN(Red_ToCheckInst_LFInst_88_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_88_LFInst_0_U3  ( .A(
        Red_MCInst2_MC3_v1_1[0] ), .B(MCInst2_MC3_v1_0 [3]), .Z(
        Red_ToCheckInst_LFInst_88_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_89_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_89_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_89_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[89])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_89_LFInst_0_U4  ( .A(MCInst2_MC2_v1_3 [2]), 
        .B(MCInst2_MC2_v1_0 [0]), .ZN(Red_ToCheckInst_LFInst_89_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_89_LFInst_0_U3  ( .A(
        Red_MCInst2_MC2_v1_1[0] ), .B(MCInst2_MC2_v1_0 [3]), .Z(
        Red_ToCheckInst_LFInst_89_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_90_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_90_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_90_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[90])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_90_LFInst_0_U4  ( .A(MCInst2_MC1_v1_3 [2]), 
        .B(MCInst2_MC1_v1_0 [0]), .ZN(Red_ToCheckInst_LFInst_90_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_90_LFInst_0_U3  ( .A(
        Red_MCInst2_MC1_v1_1[0] ), .B(MCInst2_MC1_v1_0 [3]), .Z(
        Red_ToCheckInst_LFInst_90_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_91_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_91_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_91_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[91])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_91_LFInst_0_U4  ( .A(MCInst2_MC0_v1_3 [2]), 
        .B(MCInst2_MC0_v1_0 [0]), .ZN(Red_ToCheckInst_LFInst_91_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_91_LFInst_0_U3  ( .A(
        Red_MCInst2_MC0_v1_1[0] ), .B(MCInst2_MC0_v1_0 [3]), .Z(
        Red_ToCheckInst_LFInst_91_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_92_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_92_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_92_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[92])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_92_LFInst_0_U4  ( .A(MCInst2_MC3_v0_0 [3]), 
        .B(Red_MCInst2_MC3_v0_1[0] ), .ZN(
        Red_ToCheckInst_LFInst_92_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_92_LFInst_0_U3  ( .A(MCInst2_MC3_v0_3 [3]), 
        .B(MCInst2_MC3_v0_3 [0]), .Z(Red_ToCheckInst_LFInst_92_LFInst_0_n4 )
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_93_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_93_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_93_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[93])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_93_LFInst_0_U4  ( .A(MCInst2_MC2_v0_0 [3]), 
        .B(Red_MCInst2_MC2_v0_1[0] ), .ZN(
        Red_ToCheckInst_LFInst_93_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_93_LFInst_0_U3  ( .A(MCInst2_MC2_v0_3 [3]), 
        .B(MCInst2_MC2_v0_3 [0]), .Z(Red_ToCheckInst_LFInst_93_LFInst_0_n4 )
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_94_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_94_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_94_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[94])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_94_LFInst_0_U4  ( .A(MCInst2_MC1_v0_0 [3]), 
        .B(Red_MCInst2_MC1_v0_1[0] ), .ZN(
        Red_ToCheckInst_LFInst_94_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_94_LFInst_0_U3  ( .A(MCInst2_MC1_v0_3 [3]), 
        .B(MCInst2_MC1_v0_3 [0]), .Z(Red_ToCheckInst_LFInst_94_LFInst_0_n4 )
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_95_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_95_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_95_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[95])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_95_LFInst_0_U4  ( .A(MCInst2_MC0_v0_0 [3]), 
        .B(Red_MCInst2_MC0_v0_1[0] ), .ZN(
        Red_ToCheckInst_LFInst_95_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_95_LFInst_0_U3  ( .A(MCInst2_MC0_v0_3 [3]), 
        .B(MCInst2_MC0_v0_3 [0]), .Z(Red_ToCheckInst_LFInst_95_LFInst_0_n4 )
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_96_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_96_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_96_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[96])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_96_LFInst_0_U4  ( .A(SubCellInput[1]), .B(
        SubCellInput[0]), .ZN(Red_ToCheckInst_LFInst_96_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_96_LFInst_0_U3  ( .A(SubCellInput[2]), .B(
        SubCellInput[3]), .Z(Red_ToCheckInst_LFInst_96_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_97_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_97_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_97_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[97])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_97_LFInst_0_U4  ( .A(SubCellInput[5]), .B(
        SubCellInput[4]), .ZN(Red_ToCheckInst_LFInst_97_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_97_LFInst_0_U3  ( .A(SubCellInput[6]), .B(
        SubCellInput[7]), .Z(Red_ToCheckInst_LFInst_97_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_98_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_98_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_98_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[98])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_98_LFInst_0_U4  ( .A(SubCellInput[9]), .B(
        SubCellInput[8]), .ZN(Red_ToCheckInst_LFInst_98_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_98_LFInst_0_U3  ( .A(SubCellInput[10]), .B(
        SubCellInput[11]), .Z(Red_ToCheckInst_LFInst_98_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_99_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_99_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_99_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[99])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_99_LFInst_0_U4  ( .A(SubCellInput[13]), .B(
        SubCellInput[12]), .ZN(Red_ToCheckInst_LFInst_99_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_99_LFInst_0_U3  ( .A(SubCellInput[14]), .B(
        SubCellInput[15]), .Z(Red_ToCheckInst_LFInst_99_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_100_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_100_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_100_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[100])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_100_LFInst_0_U4  ( .A(SubCellInput[17]), 
        .B(SubCellInput[16]), .ZN(Red_ToCheckInst_LFInst_100_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_100_LFInst_0_U3  ( .A(SubCellInput[18]), .B(
        SubCellInput[19]), .Z(Red_ToCheckInst_LFInst_100_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_101_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_101_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_101_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[101])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_101_LFInst_0_U4  ( .A(SubCellInput[21]), 
        .B(SubCellInput[20]), .ZN(Red_ToCheckInst_LFInst_101_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_101_LFInst_0_U3  ( .A(SubCellInput[22]), .B(
        SubCellInput[23]), .Z(Red_ToCheckInst_LFInst_101_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_102_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_102_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_102_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[102])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_102_LFInst_0_U4  ( .A(SubCellInput[25]), 
        .B(SubCellInput[24]), .ZN(Red_ToCheckInst_LFInst_102_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_102_LFInst_0_U3  ( .A(SubCellInput[26]), .B(
        SubCellInput[27]), .Z(Red_ToCheckInst_LFInst_102_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_103_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_103_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_103_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[103])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_103_LFInst_0_U4  ( .A(SubCellInput[29]), 
        .B(SubCellInput[28]), .ZN(Red_ToCheckInst_LFInst_103_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_103_LFInst_0_U3  ( .A(SubCellInput[30]), .B(
        SubCellInput[31]), .Z(Red_ToCheckInst_LFInst_103_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_104_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_104_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_104_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[104])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_104_LFInst_0_U4  ( .A(SubCellInput[33]), 
        .B(SubCellInput[32]), .ZN(Red_ToCheckInst_LFInst_104_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_104_LFInst_0_U3  ( .A(SubCellInput[34]), .B(
        SubCellInput[35]), .Z(Red_ToCheckInst_LFInst_104_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_105_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_105_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_105_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[105])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_105_LFInst_0_U4  ( .A(SubCellInput[37]), 
        .B(SubCellInput[36]), .ZN(Red_ToCheckInst_LFInst_105_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_105_LFInst_0_U3  ( .A(SubCellInput[38]), .B(
        SubCellInput[39]), .Z(Red_ToCheckInst_LFInst_105_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_106_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_106_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_106_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[106])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_106_LFInst_0_U4  ( .A(SubCellInput[41]), 
        .B(SubCellInput[40]), .ZN(Red_ToCheckInst_LFInst_106_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_106_LFInst_0_U3  ( .A(SubCellInput[42]), .B(
        SubCellInput[43]), .Z(Red_ToCheckInst_LFInst_106_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_107_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_107_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_107_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[107])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_107_LFInst_0_U4  ( .A(SubCellInput[45]), 
        .B(SubCellInput[44]), .ZN(Red_ToCheckInst_LFInst_107_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_107_LFInst_0_U3  ( .A(SubCellInput[46]), .B(
        SubCellInput[47]), .Z(Red_ToCheckInst_LFInst_107_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_108_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_108_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_108_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[108])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_108_LFInst_0_U4  ( .A(SubCellInput[49]), 
        .B(SubCellInput[48]), .ZN(Red_ToCheckInst_LFInst_108_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_108_LFInst_0_U3  ( .A(SubCellInput[50]), .B(
        SubCellInput[51]), .Z(Red_ToCheckInst_LFInst_108_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_109_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_109_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_109_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[109])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_109_LFInst_0_U4  ( .A(SubCellInput[53]), 
        .B(SubCellInput[52]), .ZN(Red_ToCheckInst_LFInst_109_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_109_LFInst_0_U3  ( .A(SubCellInput[54]), .B(
        SubCellInput[55]), .Z(Red_ToCheckInst_LFInst_109_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_110_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_110_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_110_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[110])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_110_LFInst_0_U4  ( .A(SubCellInput[57]), 
        .B(SubCellInput[56]), .ZN(Red_ToCheckInst_LFInst_110_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_110_LFInst_0_U3  ( .A(SubCellInput[58]), .B(
        SubCellInput[59]), .Z(Red_ToCheckInst_LFInst_110_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_111_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_111_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_111_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[111])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_111_LFInst_0_U4  ( .A(SubCellInput[61]), 
        .B(SubCellInput[60]), .ZN(Red_ToCheckInst_LFInst_111_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_111_LFInst_0_U3  ( .A(SubCellInput[62]), .B(
        SubCellInput[63]), .Z(Red_ToCheckInst_LFInst_111_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_112_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_112_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_112_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[112])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_112_LFInst_0_U4  ( .A(Feedback[1]), .B(
        Feedback[0]), .ZN(Red_ToCheckInst_LFInst_112_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_112_LFInst_0_U3  ( .A(Feedback[2]), .B(
        Feedback[3]), .Z(Red_ToCheckInst_LFInst_112_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_113_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_113_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_113_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[113])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_113_LFInst_0_U4  ( .A(Feedback[5]), .B(
        Feedback[4]), .ZN(Red_ToCheckInst_LFInst_113_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_113_LFInst_0_U3  ( .A(Feedback[6]), .B(
        Feedback[7]), .Z(Red_ToCheckInst_LFInst_113_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_114_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_114_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_114_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[114])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_114_LFInst_0_U4  ( .A(Feedback[9]), .B(
        Feedback[8]), .ZN(Red_ToCheckInst_LFInst_114_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_114_LFInst_0_U3  ( .A(Feedback[10]), .B(
        Feedback[11]), .Z(Red_ToCheckInst_LFInst_114_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_115_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_115_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_115_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[115])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_115_LFInst_0_U4  ( .A(Feedback[13]), .B(
        Feedback[12]), .ZN(Red_ToCheckInst_LFInst_115_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_115_LFInst_0_U3  ( .A(Feedback[14]), .B(
        Feedback[15]), .Z(Red_ToCheckInst_LFInst_115_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_116_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_116_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_116_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[116])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_116_LFInst_0_U4  ( .A(Feedback[17]), .B(
        Feedback[16]), .ZN(Red_ToCheckInst_LFInst_116_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_116_LFInst_0_U3  ( .A(Feedback[18]), .B(
        Feedback[19]), .Z(Red_ToCheckInst_LFInst_116_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_117_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_117_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_117_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[117])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_117_LFInst_0_U4  ( .A(Feedback[21]), .B(
        Feedback[20]), .ZN(Red_ToCheckInst_LFInst_117_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_117_LFInst_0_U3  ( .A(Feedback[22]), .B(
        Feedback[23]), .Z(Red_ToCheckInst_LFInst_117_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_118_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_118_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_118_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[118])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_118_LFInst_0_U4  ( .A(Feedback[25]), .B(
        Feedback[24]), .ZN(Red_ToCheckInst_LFInst_118_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_118_LFInst_0_U3  ( .A(Feedback[26]), .B(
        Feedback[27]), .Z(Red_ToCheckInst_LFInst_118_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_119_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_119_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_119_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[119])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_119_LFInst_0_U4  ( .A(Feedback[29]), .B(
        Feedback[28]), .ZN(Red_ToCheckInst_LFInst_119_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_119_LFInst_0_U3  ( .A(Feedback[30]), .B(
        Feedback[31]), .Z(Red_ToCheckInst_LFInst_119_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_120_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_120_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_120_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[120])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_120_LFInst_0_U4  ( .A(Feedback[33]), .B(
        Feedback[32]), .ZN(Red_ToCheckInst_LFInst_120_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_120_LFInst_0_U3  ( .A(Feedback[34]), .B(
        Feedback[35]), .Z(Red_ToCheckInst_LFInst_120_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_121_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_121_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_121_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[121])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_121_LFInst_0_U4  ( .A(Feedback[37]), .B(
        Feedback[36]), .ZN(Red_ToCheckInst_LFInst_121_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_121_LFInst_0_U3  ( .A(Feedback[38]), .B(
        Feedback[39]), .Z(Red_ToCheckInst_LFInst_121_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_122_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_122_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_122_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[122])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_122_LFInst_0_U4  ( .A(Feedback[41]), .B(
        Feedback[40]), .ZN(Red_ToCheckInst_LFInst_122_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_122_LFInst_0_U3  ( .A(Feedback[42]), .B(
        Feedback[43]), .Z(Red_ToCheckInst_LFInst_122_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_123_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_123_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_123_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[123])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_123_LFInst_0_U4  ( .A(Feedback[45]), .B(
        Feedback[44]), .ZN(Red_ToCheckInst_LFInst_123_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_123_LFInst_0_U3  ( .A(Feedback[46]), .B(
        Feedback[47]), .Z(Red_ToCheckInst_LFInst_123_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_124_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_124_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_124_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[124])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_124_LFInst_0_U4  ( .A(Feedback[49]), .B(
        Feedback[48]), .ZN(Red_ToCheckInst_LFInst_124_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_124_LFInst_0_U3  ( .A(Feedback[50]), .B(
        Feedback[51]), .Z(Red_ToCheckInst_LFInst_124_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_125_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_125_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_125_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[125])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_125_LFInst_0_U4  ( .A(Feedback[53]), .B(
        Feedback[52]), .ZN(Red_ToCheckInst_LFInst_125_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_125_LFInst_0_U3  ( .A(Feedback[54]), .B(
        Feedback[55]), .Z(Red_ToCheckInst_LFInst_125_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_126_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_126_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_126_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[126])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_126_LFInst_0_U4  ( .A(Feedback[57]), .B(
        Feedback[56]), .ZN(Red_ToCheckInst_LFInst_126_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_126_LFInst_0_U3  ( .A(Feedback[58]), .B(
        Feedback[59]), .Z(Red_ToCheckInst_LFInst_126_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_127_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_127_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_127_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[127])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_127_LFInst_0_U4  ( .A(Feedback[61]), .B(
        Feedback[60]), .ZN(Red_ToCheckInst_LFInst_127_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_127_LFInst_0_U3  ( .A(Feedback[62]), .B(
        Feedback[63]), .Z(Red_ToCheckInst_LFInst_127_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_128_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_128_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_128_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[128])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_128_LFInst_0_U4  ( .A(MCInst_MC3_v3_0 [2]), 
        .B(MCInst_MC3_v3_2 [3]), .ZN(Red_ToCheckInst_LFInst_128_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_128_LFInst_0_U3  ( .A(
        Red_MCInst_MC3_v3_1[0] ), .B(MCInst_MC3_v3_2 [2]), .Z(
        Red_ToCheckInst_LFInst_128_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_129_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_129_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_129_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[129])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_129_LFInst_0_U4  ( .A(MCInst_MC2_v3_0 [2]), 
        .B(MCInst_MC2_v3_2 [3]), .ZN(Red_ToCheckInst_LFInst_129_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_129_LFInst_0_U3  ( .A(
        Red_MCInst_MC2_v3_1[0] ), .B(MCInst_MC2_v3_2 [2]), .Z(
        Red_ToCheckInst_LFInst_129_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_130_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_130_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_130_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[130])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_130_LFInst_0_U4  ( .A(MCInst_MC1_v3_0 [2]), 
        .B(MCInst_MC1_v3_2 [3]), .ZN(Red_ToCheckInst_LFInst_130_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_130_LFInst_0_U3  ( .A(
        Red_MCInst_MC1_v3_1[0] ), .B(MCInst_MC1_v3_2 [2]), .Z(
        Red_ToCheckInst_LFInst_130_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_131_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_131_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_131_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[131])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_131_LFInst_0_U4  ( .A(MCInst_MC0_v3_0 [2]), 
        .B(MCInst_MC0_v3_2 [3]), .ZN(Red_ToCheckInst_LFInst_131_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_131_LFInst_0_U3  ( .A(
        Red_MCInst_MC0_v3_1[0] ), .B(MCInst_MC0_v3_2 [2]), .Z(
        Red_ToCheckInst_LFInst_131_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_132_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_132_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_132_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[132])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_132_LFInst_0_U4  ( .A(MCInst_MC3_v2_0 [2]), 
        .B(MCInst_MC3_v2_3 [1]), .ZN(Red_ToCheckInst_LFInst_132_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_132_LFInst_0_U3  ( .A(MCInst_MC3_v2_0 [3]), 
        .B(MCInst_MC3_v2_0 [0]), .Z(Red_ToCheckInst_LFInst_132_LFInst_0_n4 )
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_133_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_133_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_133_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[133])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_133_LFInst_0_U4  ( .A(MCInst_MC2_v2_0 [2]), 
        .B(MCInst_MC2_v2_3 [1]), .ZN(Red_ToCheckInst_LFInst_133_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_133_LFInst_0_U3  ( .A(MCInst_MC2_v2_0 [3]), 
        .B(MCInst_MC2_v2_0 [0]), .Z(Red_ToCheckInst_LFInst_133_LFInst_0_n4 )
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_134_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_134_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_134_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[134])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_134_LFInst_0_U4  ( .A(MCInst_MC1_v2_0 [2]), 
        .B(MCInst_MC1_v2_3 [1]), .ZN(Red_ToCheckInst_LFInst_134_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_134_LFInst_0_U3  ( .A(MCInst_MC1_v2_0 [3]), 
        .B(MCInst_MC1_v2_0 [0]), .Z(Red_ToCheckInst_LFInst_134_LFInst_0_n4 )
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_135_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_135_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_135_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[135])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_135_LFInst_0_U4  ( .A(MCInst_MC0_v2_0 [2]), 
        .B(MCInst_MC0_v2_3 [1]), .ZN(Red_ToCheckInst_LFInst_135_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_135_LFInst_0_U3  ( .A(MCInst_MC0_v2_0 [3]), 
        .B(MCInst_MC0_v2_0 [0]), .Z(Red_ToCheckInst_LFInst_135_LFInst_0_n4 )
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_136_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_136_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_136_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[136])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_136_LFInst_0_U4  ( .A(MCInst_MC3_v1_3 [2]), 
        .B(MCInst_MC3_v1_0 [0]), .ZN(Red_ToCheckInst_LFInst_136_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_136_LFInst_0_U3  ( .A(
        Red_MCInst_MC3_v1_1[0] ), .B(MCInst_MC3_v1_0 [3]), .Z(
        Red_ToCheckInst_LFInst_136_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_137_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_137_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_137_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[137])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_137_LFInst_0_U4  ( .A(MCInst_MC2_v1_3 [2]), 
        .B(MCInst_MC2_v1_0 [0]), .ZN(Red_ToCheckInst_LFInst_137_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_137_LFInst_0_U3  ( .A(
        Red_MCInst_MC2_v1_1[0] ), .B(MCInst_MC2_v1_0 [3]), .Z(
        Red_ToCheckInst_LFInst_137_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_138_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_138_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_138_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[138])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_138_LFInst_0_U4  ( .A(MCInst_MC1_v1_3 [2]), 
        .B(MCInst_MC1_v1_0 [0]), .ZN(Red_ToCheckInst_LFInst_138_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_138_LFInst_0_U3  ( .A(
        Red_MCInst_MC1_v1_1[0] ), .B(MCInst_MC1_v1_0 [3]), .Z(
        Red_ToCheckInst_LFInst_138_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_139_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_139_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_139_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[139])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_139_LFInst_0_U4  ( .A(MCInst_MC0_v1_3 [2]), 
        .B(MCInst_MC0_v1_0 [0]), .ZN(Red_ToCheckInst_LFInst_139_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_139_LFInst_0_U3  ( .A(
        Red_MCInst_MC0_v1_1[0] ), .B(MCInst_MC0_v1_0 [3]), .Z(
        Red_ToCheckInst_LFInst_139_LFInst_0_n4 ) );
  XNOR2_X1 Red_ToCheckInst_LFInst_140_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_140_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_140_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[140])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_140_LFInst_0_U4  ( .A(MCInst_MC3_v0_0 [3]), 
        .B(Red_MCInst_MC3_v0_1[0] ), .ZN(
        Red_ToCheckInst_LFInst_140_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_140_LFInst_0_U3  ( .A(MCInst_MC3_v0_3 [3]), 
        .B(MCInst_MC3_v0_3 [0]), .Z(Red_ToCheckInst_LFInst_140_LFInst_0_n4 )
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_141_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_141_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_141_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[141])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_141_LFInst_0_U4  ( .A(MCInst_MC2_v0_0 [3]), 
        .B(Red_MCInst_MC2_v0_1[0] ), .ZN(
        Red_ToCheckInst_LFInst_141_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_141_LFInst_0_U3  ( .A(MCInst_MC2_v0_3 [3]), 
        .B(MCInst_MC2_v0_3 [0]), .Z(Red_ToCheckInst_LFInst_141_LFInst_0_n4 )
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_142_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_142_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_142_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[142])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_142_LFInst_0_U4  ( .A(MCInst_MC1_v0_0 [3]), 
        .B(Red_MCInst_MC1_v0_1[0] ), .ZN(
        Red_ToCheckInst_LFInst_142_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_142_LFInst_0_U3  ( .A(MCInst_MC1_v0_3 [3]), 
        .B(MCInst_MC1_v0_3 [0]), .Z(Red_ToCheckInst_LFInst_142_LFInst_0_n4 )
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_143_LFInst_0_U5  ( .A(
        Red_ToCheckInst_LFInst_143_LFInst_0_n4 ), .B(
        Red_ToCheckInst_LFInst_143_LFInst_0_n3 ), .ZN(Red_SignaltoCheck[143])
         );
  XNOR2_X1 Red_ToCheckInst_LFInst_143_LFInst_0_U4  ( .A(MCInst_MC0_v0_0 [3]), 
        .B(Red_MCInst_MC0_v0_1[0] ), .ZN(
        Red_ToCheckInst_LFInst_143_LFInst_0_n3 ) );
  XOR2_X1 Red_ToCheckInst_LFInst_143_LFInst_0_U3  ( .A(MCInst_MC0_v0_3 [3]), 
        .B(MCInst_MC0_v0_3 [0]), .Z(Red_ToCheckInst_LFInst_143_LFInst_0_n4 )
         );
  NOR2_X1 Check1_CheckInst_0_U287  ( .A1(Check1_CheckInst_0_n286 ), .A2(
        Check1_CheckInst_0_n285 ), .ZN(Error[0] ) );
  NAND2_X1 Check1_CheckInst_0_U286  ( .A1(Check1_CheckInst_0_n284 ), .A2(
        Check1_CheckInst_0_n283 ), .ZN(Check1_CheckInst_0_n285 ) );
  NOR2_X1 Check1_CheckInst_0_U285  ( .A1(Check1_CheckInst_0_n282 ), .A2(
        Check1_CheckInst_0_n281 ), .ZN(Check1_CheckInst_0_n283 ) );
  NAND2_X1 Check1_CheckInst_0_U284  ( .A1(Check1_CheckInst_0_n280 ), .A2(
        Check1_CheckInst_0_n279 ), .ZN(Check1_CheckInst_0_n281 ) );
  NOR2_X1 Check1_CheckInst_0_U283  ( .A1(Check1_CheckInst_0_n278 ), .A2(
        Check1_CheckInst_0_n277 ), .ZN(Check1_CheckInst_0_n279 ) );
  NAND2_X1 Check1_CheckInst_0_U282  ( .A1(Check1_CheckInst_0_n276 ), .A2(
        Check1_CheckInst_0_n275 ), .ZN(Check1_CheckInst_0_n277 ) );
  NOR2_X1 Check1_CheckInst_0_U281  ( .A1(Check1_CheckInst_0_n274 ), .A2(
        Check1_CheckInst_0_n273 ), .ZN(Check1_CheckInst_0_n275 ) );
  NAND2_X1 Check1_CheckInst_0_U280  ( .A1(Check1_CheckInst_0_n272 ), .A2(
        Check1_CheckInst_0_n271 ), .ZN(Check1_CheckInst_0_n273 ) );
  NOR2_X1 Check1_CheckInst_0_U279  ( .A1(Check1_CheckInst_0_n270 ), .A2(
        Check1_CheckInst_0_n269 ), .ZN(Check1_CheckInst_0_n271 ) );
  NAND2_X1 Check1_CheckInst_0_U278  ( .A1(Check1_CheckInst_0_n268 ), .A2(
        Check1_CheckInst_0_n267 ), .ZN(Check1_CheckInst_0_n269 ) );
  NOR2_X1 Check1_CheckInst_0_U277  ( .A1(Check1_CheckInst_0_n266 ), .A2(
        Check1_CheckInst_0_n265 ), .ZN(Check1_CheckInst_0_n267 ) );
  XOR2_X1 Check1_CheckInst_0_U276  ( .A(Red_SubCellInput2[5]), .B(
        Red_SignaltoCheck[53]), .Z(Check1_CheckInst_0_n265 ) );
  XOR2_X1 Check1_CheckInst_0_U275  ( .A(Red_SubCellInput2[6]), .B(
        Red_SignaltoCheck[54]), .Z(Check1_CheckInst_0_n266 ) );
  NOR2_X1 Check1_CheckInst_0_U274  ( .A1(Check1_CheckInst_0_n264 ), .A2(
        Check1_CheckInst_0_n263 ), .ZN(Check1_CheckInst_0_n268 ) );
  XOR2_X1 Check1_CheckInst_0_U273  ( .A(Red_SubCellInput2[9]), .B(
        Red_SignaltoCheck[57]), .Z(Check1_CheckInst_0_n263 ) );
  XOR2_X1 Check1_CheckInst_0_U272  ( .A(Red_SubCellInput2[8]), .B(
        Red_SignaltoCheck[56]), .Z(Check1_CheckInst_0_n264 ) );
  NAND2_X1 Check1_CheckInst_0_U271  ( .A1(Check1_CheckInst_0_n262 ), .A2(
        Check1_CheckInst_0_n261 ), .ZN(Check1_CheckInst_0_n270 ) );
  NOR2_X1 Check1_CheckInst_0_U270  ( .A1(Check1_CheckInst_0_n260 ), .A2(
        Check1_CheckInst_0_n259 ), .ZN(Check1_CheckInst_0_n261 ) );
  XOR2_X1 Check1_CheckInst_0_U269  ( .A(Red_Feedback2[3]), .B(
        Red_SignaltoCheck[67]), .Z(Check1_CheckInst_0_n259 ) );
  XOR2_X1 Check1_CheckInst_0_U268  ( .A(Red_Feedback2[6]), .B(
        Red_SignaltoCheck[70]), .Z(Check1_CheckInst_0_n260 ) );
  NOR2_X1 Check1_CheckInst_0_U267  ( .A1(Check1_CheckInst_0_n258 ), .A2(
        Check1_CheckInst_0_n257 ), .ZN(Check1_CheckInst_0_n262 ) );
  XOR2_X1 Check1_CheckInst_0_U266  ( .A(Red_Feedback2[5]), .B(
        Red_SignaltoCheck[69]), .Z(Check1_CheckInst_0_n257 ) );
  XOR2_X1 Check1_CheckInst_0_U265  ( .A(Red_SubCellInput2[7]), .B(
        Red_SignaltoCheck[55]), .Z(Check1_CheckInst_0_n258 ) );
  NOR2_X1 Check1_CheckInst_0_U264  ( .A1(Check1_CheckInst_0_n256 ), .A2(
        Check1_CheckInst_0_n255 ), .ZN(Check1_CheckInst_0_n272 ) );
  NAND2_X1 Check1_CheckInst_0_U263  ( .A1(Check1_CheckInst_0_n254 ), .A2(
        Check1_CheckInst_0_n253 ), .ZN(Check1_CheckInst_0_n255 ) );
  XNOR2_X1 Check1_CheckInst_0_U262  ( .A(Red_SubCellInput2[15]), .B(
        Red_SignaltoCheck[63]), .ZN(Check1_CheckInst_0_n253 ) );
  XNOR2_X1 Check1_CheckInst_0_U261  ( .A(Red_Feedback2[2]), .B(
        Red_SignaltoCheck[66]), .ZN(Check1_CheckInst_0_n254 ) );
  NAND2_X1 Check1_CheckInst_0_U260  ( .A1(Check1_CheckInst_0_n252 ), .A2(
        Check1_CheckInst_0_n251 ), .ZN(Check1_CheckInst_0_n256 ) );
  XNOR2_X1 Check1_CheckInst_0_U259  ( .A(Red_Feedback2[1]), .B(
        Red_SignaltoCheck[65]), .ZN(Check1_CheckInst_0_n251 ) );
  XNOR2_X1 Check1_CheckInst_0_U258  ( .A(Red_Feedback2[4]), .B(
        Red_SignaltoCheck[68]), .ZN(Check1_CheckInst_0_n252 ) );
  NAND2_X1 Check1_CheckInst_0_U257  ( .A1(Check1_CheckInst_0_n250 ), .A2(
        Check1_CheckInst_0_n249 ), .ZN(Check1_CheckInst_0_n274 ) );
  NOR2_X1 Check1_CheckInst_0_U256  ( .A1(Check1_CheckInst_0_n248 ), .A2(
        Check1_CheckInst_0_n247 ), .ZN(Check1_CheckInst_0_n249 ) );
  XOR2_X1 Check1_CheckInst_0_U255  ( .A(Red_ShiftRowsOutput3[11]), .B(
        Red_SignaltoCheck[43]), .Z(Check1_CheckInst_0_n247 ) );
  XOR2_X1 Check1_CheckInst_0_U254  ( .A(Red_ShiftRowsOutput3[10]), .B(
        Red_SignaltoCheck[42]), .Z(Check1_CheckInst_0_n248 ) );
  NOR2_X1 Check1_CheckInst_0_U253  ( .A1(Check1_CheckInst_0_n246 ), .A2(
        Check1_CheckInst_0_n245 ), .ZN(Check1_CheckInst_0_n250 ) );
  XOR2_X1 Check1_CheckInst_0_U252  ( .A(Red_Feedback2[0]), .B(
        Red_SignaltoCheck[64]), .Z(Check1_CheckInst_0_n245 ) );
  XOR2_X1 Check1_CheckInst_0_U251  ( .A(Red_SubCellInput2[14]), .B(
        Red_SignaltoCheck[62]), .Z(Check1_CheckInst_0_n246 ) );
  NOR2_X1 Check1_CheckInst_0_U250  ( .A1(Check1_CheckInst_0_n244 ), .A2(
        Check1_CheckInst_0_n243 ), .ZN(Check1_CheckInst_0_n276 ) );
  NAND2_X1 Check1_CheckInst_0_U249  ( .A1(Check1_CheckInst_0_n242 ), .A2(
        Check1_CheckInst_0_n241 ), .ZN(Check1_CheckInst_0_n243 ) );
  NOR2_X1 Check1_CheckInst_0_U248  ( .A1(Check1_CheckInst_0_n240 ), .A2(
        Check1_CheckInst_0_n239 ), .ZN(Check1_CheckInst_0_n241 ) );
  NAND2_X1 Check1_CheckInst_0_U247  ( .A1(Check1_CheckInst_0_n238 ), .A2(
        Check1_CheckInst_0_n237 ), .ZN(Check1_CheckInst_0_n239 ) );
  NOR2_X1 Check1_CheckInst_0_U246  ( .A1(Check1_CheckInst_0_n236 ), .A2(
        Check1_CheckInst_0_n235 ), .ZN(Check1_CheckInst_0_n237 ) );
  XOR2_X1 Check1_CheckInst_0_U245  ( .A(Red_ShiftRowsOutput3[7]), .B(
        Red_SignaltoCheck[39]), .Z(Check1_CheckInst_0_n235 ) );
  XOR2_X1 Check1_CheckInst_0_U244  ( .A(Red_ShiftRowsOutput3[6]), .B(
        Red_SignaltoCheck[38]), .Z(Check1_CheckInst_0_n236 ) );
  NOR2_X1 Check1_CheckInst_0_U243  ( .A1(Check1_CheckInst_0_n234 ), .A2(
        Check1_CheckInst_0_n233 ), .ZN(Check1_CheckInst_0_n238 ) );
  XOR2_X1 Check1_CheckInst_0_U242  ( .A(Red_ShiftRowsOutput3[9]), .B(
        Red_SignaltoCheck[41]), .Z(Check1_CheckInst_0_n233 ) );
  XOR2_X1 Check1_CheckInst_0_U241  ( .A(Red_ShiftRowsOutput3[8]), .B(
        Red_SignaltoCheck[40]), .Z(Check1_CheckInst_0_n234 ) );
  NAND2_X1 Check1_CheckInst_0_U240  ( .A1(Check1_CheckInst_0_n232 ), .A2(
        Check1_CheckInst_0_n231 ), .ZN(Check1_CheckInst_0_n240 ) );
  NOR2_X1 Check1_CheckInst_0_U239  ( .A1(Check1_CheckInst_0_n230 ), .A2(
        Check1_CheckInst_0_n229 ), .ZN(Check1_CheckInst_0_n231 ) );
  XOR2_X1 Check1_CheckInst_0_U238  ( .A(Red_SubCellInput2[3]), .B(
        Red_SignaltoCheck[51]), .Z(Check1_CheckInst_0_n229 ) );
  XOR2_X1 Check1_CheckInst_0_U237  ( .A(Red_ShiftRowsOutput3[5]), .B(
        Red_SignaltoCheck[37]), .Z(Check1_CheckInst_0_n230 ) );
  NOR2_X1 Check1_CheckInst_0_U236  ( .A1(Check1_CheckInst_0_n228 ), .A2(
        Check1_CheckInst_0_n227 ), .ZN(Check1_CheckInst_0_n232 ) );
  XOR2_X1 Check1_CheckInst_0_U235  ( .A(Red_ShiftRowsOutput3[3]), .B(
        Red_SignaltoCheck[35]), .Z(Check1_CheckInst_0_n227 ) );
  XOR2_X1 Check1_CheckInst_0_U234  ( .A(Red_ShiftRowsOutput3[4]), .B(
        Red_SignaltoCheck[36]), .Z(Check1_CheckInst_0_n228 ) );
  NOR2_X1 Check1_CheckInst_0_U233  ( .A1(Check1_CheckInst_0_n226 ), .A2(
        Check1_CheckInst_0_n225 ), .ZN(Check1_CheckInst_0_n242 ) );
  NAND2_X1 Check1_CheckInst_0_U232  ( .A1(Check1_CheckInst_0_n224 ), .A2(
        Check1_CheckInst_0_n223 ), .ZN(Check1_CheckInst_0_n225 ) );
  XNOR2_X1 Check1_CheckInst_0_U231  ( .A(Red_ShiftRowsOutput3[15]), .B(
        Red_SignaltoCheck[47]), .ZN(Check1_CheckInst_0_n223 ) );
  XNOR2_X1 Check1_CheckInst_0_U230  ( .A(Red_SubCellInput2[2]), .B(
        Red_SignaltoCheck[50]), .ZN(Check1_CheckInst_0_n224 ) );
  NAND2_X1 Check1_CheckInst_0_U229  ( .A1(Check1_CheckInst_0_n222 ), .A2(
        Check1_CheckInst_0_n221 ), .ZN(Check1_CheckInst_0_n226 ) );
  XNOR2_X1 Check1_CheckInst_0_U228  ( .A(Red_SubCellInput2[1]), .B(
        Red_SignaltoCheck[49]), .ZN(Check1_CheckInst_0_n221 ) );
  XNOR2_X1 Check1_CheckInst_0_U227  ( .A(Red_SubCellInput2[4]), .B(
        Red_SignaltoCheck[52]), .ZN(Check1_CheckInst_0_n222 ) );
  NAND2_X1 Check1_CheckInst_0_U226  ( .A1(Check1_CheckInst_0_n220 ), .A2(
        Check1_CheckInst_0_n219 ), .ZN(Check1_CheckInst_0_n244 ) );
  NOR2_X1 Check1_CheckInst_0_U225  ( .A1(Check1_CheckInst_0_n218 ), .A2(
        Check1_CheckInst_0_n217 ), .ZN(Check1_CheckInst_0_n219 ) );
  XOR2_X1 Check1_CheckInst_0_U224  ( .A(Red_ShiftRowsOutput3[14]), .B(
        Red_SignaltoCheck[46]), .Z(Check1_CheckInst_0_n217 ) );
  XOR2_X1 Check1_CheckInst_0_U223  ( .A(Red_ShiftRowsOutput3[12]), .B(
        Red_SignaltoCheck[44]), .Z(Check1_CheckInst_0_n218 ) );
  NOR2_X1 Check1_CheckInst_0_U222  ( .A1(Check1_CheckInst_0_n216 ), .A2(
        Check1_CheckInst_0_n215 ), .ZN(Check1_CheckInst_0_n220 ) );
  XOR2_X1 Check1_CheckInst_0_U221  ( .A(Red_ShiftRowsOutput3[13]), .B(
        Red_SignaltoCheck[45]), .Z(Check1_CheckInst_0_n215 ) );
  XOR2_X1 Check1_CheckInst_0_U220  ( .A(Red_SubCellInput2[0]), .B(
        Red_SignaltoCheck[48]), .Z(Check1_CheckInst_0_n216 ) );
  NAND2_X1 Check1_CheckInst_0_U219  ( .A1(Check1_CheckInst_0_n214 ), .A2(
        Check1_CheckInst_0_n213 ), .ZN(Check1_CheckInst_0_n278 ) );
  NOR2_X1 Check1_CheckInst_0_U218  ( .A1(Check1_CheckInst_0_n212 ), .A2(
        Check1_CheckInst_0_n211 ), .ZN(Check1_CheckInst_0_n213 ) );
  NAND2_X1 Check1_CheckInst_0_U217  ( .A1(Check1_CheckInst_0_n210 ), .A2(
        Check1_CheckInst_0_n209 ), .ZN(Check1_CheckInst_0_n211 ) );
  NOR2_X1 Check1_CheckInst_0_U216  ( .A1(Check1_CheckInst_0_n208 ), .A2(
        Check1_CheckInst_0_n207 ), .ZN(Check1_CheckInst_0_n209 ) );
  XOR2_X1 Check1_CheckInst_0_U215  ( .A(Red_SubCellInput[1]), .B(
        Red_SignaltoCheck[97]), .Z(Check1_CheckInst_0_n207 ) );
  XOR2_X1 Check1_CheckInst_0_U214  ( .A(Red_SubCellInput[0]), .B(
        Red_SignaltoCheck[96]), .Z(Check1_CheckInst_0_n208 ) );
  NOR2_X1 Check1_CheckInst_0_U213  ( .A1(Check1_CheckInst_0_n206 ), .A2(
        Check1_CheckInst_0_n205 ), .ZN(Check1_CheckInst_0_n210 ) );
  XOR2_X1 Check1_CheckInst_0_U212  ( .A(Red_ShiftRowsOutput2[15]), .B(
        Red_SignaltoCheck[95]), .Z(Check1_CheckInst_0_n205 ) );
  XOR2_X1 Check1_CheckInst_0_U211  ( .A(Red_ShiftRowsOutput2[14]), .B(
        Red_SignaltoCheck[94]), .Z(Check1_CheckInst_0_n206 ) );
  NAND2_X1 Check1_CheckInst_0_U210  ( .A1(Check1_CheckInst_0_n204 ), .A2(
        Check1_CheckInst_0_n203 ), .ZN(Check1_CheckInst_0_n212 ) );
  XNOR2_X1 Check1_CheckInst_0_U209  ( .A(Red_ShiftRowsOutput2[13]), .B(
        Red_SignaltoCheck[93]), .ZN(Check1_CheckInst_0_n203 ) );
  XNOR2_X1 Check1_CheckInst_0_U208  ( .A(Red_ShiftRowsOutput2[12]), .B(
        Red_SignaltoCheck[92]), .ZN(Check1_CheckInst_0_n204 ) );
  NOR2_X1 Check1_CheckInst_0_U207  ( .A1(Check1_CheckInst_0_n202 ), .A2(
        Check1_CheckInst_0_n201 ), .ZN(Check1_CheckInst_0_n214 ) );
  XOR2_X1 Check1_CheckInst_0_U206  ( .A(Red_ShiftRowsOutput2[9]), .B(
        Red_SignaltoCheck[89]), .Z(Check1_CheckInst_0_n201 ) );
  XOR2_X1 Check1_CheckInst_0_U205  ( .A(Red_ShiftRowsOutput2[10]), .B(
        Red_SignaltoCheck[90]), .Z(Check1_CheckInst_0_n202 ) );
  NOR2_X1 Check1_CheckInst_0_U204  ( .A1(Check1_CheckInst_0_n200 ), .A2(
        Check1_CheckInst_0_n199 ), .ZN(Check1_CheckInst_0_n280 ) );
  NAND2_X1 Check1_CheckInst_0_U203  ( .A1(Check1_CheckInst_0_n198 ), .A2(
        Check1_CheckInst_0_n197 ), .ZN(Check1_CheckInst_0_n199 ) );
  NOR2_X1 Check1_CheckInst_0_U202  ( .A1(Check1_CheckInst_0_n196 ), .A2(
        Check1_CheckInst_0_n195 ), .ZN(Check1_CheckInst_0_n197 ) );
  NAND2_X1 Check1_CheckInst_0_U201  ( .A1(Check1_CheckInst_0_n194 ), .A2(
        Check1_CheckInst_0_n193 ), .ZN(Check1_CheckInst_0_n195 ) );
  XNOR2_X1 Check1_CheckInst_0_U200  ( .A(Red_SubCellInput[9]), .B(
        Red_SignaltoCheck[105]), .ZN(Check1_CheckInst_0_n193 ) );
  XNOR2_X1 Check1_CheckInst_0_U199  ( .A(Red_ShiftRowsOutput2[11]), .B(
        Red_SignaltoCheck[91]), .ZN(Check1_CheckInst_0_n194 ) );
  NAND2_X1 Check1_CheckInst_0_U198  ( .A1(Check1_CheckInst_0_n192 ), .A2(
        Check1_CheckInst_0_n191 ), .ZN(Check1_CheckInst_0_n196 ) );
  XNOR2_X1 Check1_CheckInst_0_U197  ( .A(Red_SubCellInput[7]), .B(
        Red_SignaltoCheck[103]), .ZN(Check1_CheckInst_0_n191 ) );
  XNOR2_X1 Check1_CheckInst_0_U196  ( .A(Red_SubCellInput[10]), .B(
        Red_SignaltoCheck[106]), .ZN(Check1_CheckInst_0_n192 ) );
  NOR2_X1 Check1_CheckInst_0_U195  ( .A1(Check1_CheckInst_0_n190 ), .A2(
        Check1_CheckInst_0_n189 ), .ZN(Check1_CheckInst_0_n198 ) );
  XOR2_X1 Check1_CheckInst_0_U194  ( .A(Red_SubCellInput[5]), .B(
        Red_SignaltoCheck[101]), .Z(Check1_CheckInst_0_n189 ) );
  XOR2_X1 Check1_CheckInst_0_U193  ( .A(Red_SubCellInput[8]), .B(
        Red_SignaltoCheck[104]), .Z(Check1_CheckInst_0_n190 ) );
  NAND2_X1 Check1_CheckInst_0_U192  ( .A1(Check1_CheckInst_0_n188 ), .A2(
        Check1_CheckInst_0_n187 ), .ZN(Check1_CheckInst_0_n200 ) );
  XNOR2_X1 Check1_CheckInst_0_U191  ( .A(Red_SubCellInput[3]), .B(
        Red_SignaltoCheck[99]), .ZN(Check1_CheckInst_0_n187 ) );
  XNOR2_X1 Check1_CheckInst_0_U190  ( .A(Red_SubCellInput[6]), .B(
        Red_SignaltoCheck[102]), .ZN(Check1_CheckInst_0_n188 ) );
  NAND2_X1 Check1_CheckInst_0_U189  ( .A1(Check1_CheckInst_0_n186 ), .A2(
        Check1_CheckInst_0_n185 ), .ZN(Check1_CheckInst_0_n282 ) );
  NOR2_X1 Check1_CheckInst_0_U188  ( .A1(Check1_CheckInst_0_n184 ), .A2(
        Check1_CheckInst_0_n183 ), .ZN(Check1_CheckInst_0_n185 ) );
  NAND2_X1 Check1_CheckInst_0_U187  ( .A1(Check1_CheckInst_0_n182 ), .A2(
        Check1_CheckInst_0_n181 ), .ZN(Check1_CheckInst_0_n183 ) );
  NOR2_X1 Check1_CheckInst_0_U186  ( .A1(Check1_CheckInst_0_n180 ), .A2(
        Check1_CheckInst_0_n179 ), .ZN(Check1_CheckInst_0_n181 ) );
  NAND2_X1 Check1_CheckInst_0_U185  ( .A1(Check1_CheckInst_0_n178 ), .A2(
        Check1_CheckInst_0_n177 ), .ZN(Check1_CheckInst_0_n179 ) );
  NOR2_X1 Check1_CheckInst_0_U184  ( .A1(Check1_CheckInst_0_n176 ), .A2(
        Check1_CheckInst_0_n175 ), .ZN(Check1_CheckInst_0_n177 ) );
  NAND2_X1 Check1_CheckInst_0_U183  ( .A1(Check1_CheckInst_0_n174 ), .A2(
        Check1_CheckInst_0_n173 ), .ZN(Check1_CheckInst_0_n175 ) );
  XNOR2_X1 Check1_CheckInst_0_U182  ( .A(Red_SubCellInput[4]), .B(
        Red_SignaltoCheck[100]), .ZN(Check1_CheckInst_0_n173 ) );
  XNOR2_X1 Check1_CheckInst_0_U181  ( .A(Red_SubCellInput[2]), .B(
        Red_SignaltoCheck[98]), .ZN(Check1_CheckInst_0_n174 ) );
  NAND2_X1 Check1_CheckInst_0_U180  ( .A1(Check1_CheckInst_0_n172 ), .A2(
        Check1_CheckInst_0_n171 ), .ZN(Check1_CheckInst_0_n176 ) );
  XNOR2_X1 Check1_CheckInst_0_U179  ( .A(Red_Feedback2[15]), .B(
        Red_SignaltoCheck[79]), .ZN(Check1_CheckInst_0_n171 ) );
  XNOR2_X1 Check1_CheckInst_0_U178  ( .A(Red_Feedback2[14]), .B(
        Red_SignaltoCheck[78]), .ZN(Check1_CheckInst_0_n172 ) );
  NOR2_X1 Check1_CheckInst_0_U177  ( .A1(Check1_CheckInst_0_n170 ), .A2(
        Check1_CheckInst_0_n169 ), .ZN(Check1_CheckInst_0_n178 ) );
  XOR2_X1 Check1_CheckInst_0_U176  ( .A(Red_Feedback2[13]), .B(
        Red_SignaltoCheck[77]), .Z(Check1_CheckInst_0_n169 ) );
  XOR2_X1 Check1_CheckInst_0_U175  ( .A(Red_Feedback2[12]), .B(
        Red_SignaltoCheck[76]), .Z(Check1_CheckInst_0_n170 ) );
  NAND2_X1 Check1_CheckInst_0_U174  ( .A1(Check1_CheckInst_0_n168 ), .A2(
        Check1_CheckInst_0_n167 ), .ZN(Check1_CheckInst_0_n180 ) );
  XNOR2_X1 Check1_CheckInst_0_U173  ( .A(Red_Feedback2[11]), .B(
        Red_SignaltoCheck[75]), .ZN(Check1_CheckInst_0_n167 ) );
  XNOR2_X1 Check1_CheckInst_0_U172  ( .A(Red_Feedback2[10]), .B(
        Red_SignaltoCheck[74]), .ZN(Check1_CheckInst_0_n168 ) );
  NOR2_X1 Check1_CheckInst_0_U171  ( .A1(Check1_CheckInst_0_n166 ), .A2(
        Check1_CheckInst_0_n165 ), .ZN(Check1_CheckInst_0_n182 ) );
  NAND2_X1 Check1_CheckInst_0_U170  ( .A1(Check1_CheckInst_0_n164 ), .A2(
        Check1_CheckInst_0_n163 ), .ZN(Check1_CheckInst_0_n165 ) );
  NOR2_X1 Check1_CheckInst_0_U169  ( .A1(Check1_CheckInst_0_n162 ), .A2(
        Check1_CheckInst_0_n161 ), .ZN(Check1_CheckInst_0_n163 ) );
  NAND2_X1 Check1_CheckInst_0_U168  ( .A1(Check1_CheckInst_0_n160 ), .A2(
        Check1_CheckInst_0_n159 ), .ZN(Check1_CheckInst_0_n161 ) );
  XNOR2_X1 Check1_CheckInst_0_U167  ( .A(Red_Feedback2[7]), .B(
        Red_SignaltoCheck[71]), .ZN(Check1_CheckInst_0_n159 ) );
  XNOR2_X1 Check1_CheckInst_0_U166  ( .A(Red_Feedback2[8]), .B(
        Red_SignaltoCheck[72]), .ZN(Check1_CheckInst_0_n160 ) );
  NAND2_X1 Check1_CheckInst_0_U165  ( .A1(Check1_CheckInst_0_n158 ), .A2(
        Check1_CheckInst_0_n157 ), .ZN(Check1_CheckInst_0_n162 ) );
  XNOR2_X1 Check1_CheckInst_0_U164  ( .A(Red_ShiftRowsOutput2[7]), .B(
        Red_SignaltoCheck[87]), .ZN(Check1_CheckInst_0_n157 ) );
  XNOR2_X1 Check1_CheckInst_0_U163  ( .A(Red_Feedback2[9]), .B(
        Red_SignaltoCheck[73]), .ZN(Check1_CheckInst_0_n158 ) );
  NOR2_X1 Check1_CheckInst_0_U162  ( .A1(Check1_CheckInst_0_n156 ), .A2(
        Check1_CheckInst_0_n155 ), .ZN(Check1_CheckInst_0_n164 ) );
  XOR2_X1 Check1_CheckInst_0_U161  ( .A(Red_ShiftRowsOutput2[5]), .B(
        Red_SignaltoCheck[85]), .Z(Check1_CheckInst_0_n155 ) );
  XOR2_X1 Check1_CheckInst_0_U160  ( .A(Red_ShiftRowsOutput2[8]), .B(
        Red_SignaltoCheck[88]), .Z(Check1_CheckInst_0_n156 ) );
  NAND2_X1 Check1_CheckInst_0_U159  ( .A1(Check1_CheckInst_0_n154 ), .A2(
        Check1_CheckInst_0_n153 ), .ZN(Check1_CheckInst_0_n166 ) );
  XNOR2_X1 Check1_CheckInst_0_U158  ( .A(Red_ShiftRowsOutput2[3]), .B(
        Red_SignaltoCheck[83]), .ZN(Check1_CheckInst_0_n153 ) );
  XNOR2_X1 Check1_CheckInst_0_U157  ( .A(Red_ShiftRowsOutput2[6]), .B(
        Red_SignaltoCheck[86]), .ZN(Check1_CheckInst_0_n154 ) );
  NAND2_X1 Check1_CheckInst_0_U156  ( .A1(Check1_CheckInst_0_n152 ), .A2(
        Check1_CheckInst_0_n151 ), .ZN(Check1_CheckInst_0_n184 ) );
  NOR2_X1 Check1_CheckInst_0_U155  ( .A1(Check1_CheckInst_0_n150 ), .A2(
        Check1_CheckInst_0_n149 ), .ZN(Check1_CheckInst_0_n151 ) );
  NAND2_X1 Check1_CheckInst_0_U154  ( .A1(Check1_CheckInst_0_n148 ), .A2(
        Check1_CheckInst_0_n147 ), .ZN(Check1_CheckInst_0_n149 ) );
  NOR2_X1 Check1_CheckInst_0_U153  ( .A1(Check1_CheckInst_0_n146 ), .A2(
        Check1_CheckInst_0_n145 ), .ZN(Check1_CheckInst_0_n147 ) );
  XOR2_X1 Check1_CheckInst_0_U152  ( .A(Red_ShiftRowsOutput2[1]), .B(
        Red_SignaltoCheck[81]), .Z(Check1_CheckInst_0_n145 ) );
  XOR2_X1 Check1_CheckInst_0_U151  ( .A(Red_ShiftRowsOutput2[4]), .B(
        Red_SignaltoCheck[84]), .Z(Check1_CheckInst_0_n146 ) );
  NOR2_X1 Check1_CheckInst_0_U150  ( .A1(Check1_CheckInst_0_n144 ), .A2(
        Check1_CheckInst_0_n143 ), .ZN(Check1_CheckInst_0_n148 ) );
  XOR2_X1 Check1_CheckInst_0_U149  ( .A(Red_ShiftRowsOutput2[2]), .B(
        Red_SignaltoCheck[82]), .Z(Check1_CheckInst_0_n143 ) );
  XOR2_X1 Check1_CheckInst_0_U148  ( .A(Red_ShiftRowsOutput2[0]), .B(
        Red_SignaltoCheck[80]), .Z(Check1_CheckInst_0_n144 ) );
  NAND2_X1 Check1_CheckInst_0_U147  ( .A1(Check1_CheckInst_0_n142 ), .A2(
        Check1_CheckInst_0_n141 ), .ZN(Check1_CheckInst_0_n150 ) );
  XNOR2_X1 Check1_CheckInst_0_U146  ( .A(Red_ShiftRowsOutput[5]), .B(
        Red_SignaltoCheck[133]), .ZN(Check1_CheckInst_0_n141 ) );
  XNOR2_X1 Check1_CheckInst_0_U145  ( .A(Red_ShiftRowsOutput[4]), .B(
        Red_SignaltoCheck[132]), .ZN(Check1_CheckInst_0_n142 ) );
  NOR2_X1 Check1_CheckInst_0_U144  ( .A1(Check1_CheckInst_0_n140 ), .A2(
        Check1_CheckInst_0_n139 ), .ZN(Check1_CheckInst_0_n152 ) );
  XOR2_X1 Check1_CheckInst_0_U143  ( .A(Red_ShiftRowsOutput[3]), .B(
        Red_SignaltoCheck[131]), .Z(Check1_CheckInst_0_n139 ) );
  XOR2_X1 Check1_CheckInst_0_U142  ( .A(Red_ShiftRowsOutput[2]), .B(
        Red_SignaltoCheck[130]), .Z(Check1_CheckInst_0_n140 ) );
  NOR2_X1 Check1_CheckInst_0_U141  ( .A1(Check1_CheckInst_0_n138 ), .A2(
        Check1_CheckInst_0_n137 ), .ZN(Check1_CheckInst_0_n186 ) );
  NAND2_X1 Check1_CheckInst_0_U140  ( .A1(Check1_CheckInst_0_n136 ), .A2(
        Check1_CheckInst_0_n135 ), .ZN(Check1_CheckInst_0_n137 ) );
  NOR2_X1 Check1_CheckInst_0_U139  ( .A1(Check1_CheckInst_0_n134 ), .A2(
        Check1_CheckInst_0_n133 ), .ZN(Check1_CheckInst_0_n135 ) );
  NAND2_X1 Check1_CheckInst_0_U138  ( .A1(Check1_CheckInst_0_n132 ), .A2(
        Check1_CheckInst_0_n131 ), .ZN(Check1_CheckInst_0_n133 ) );
  XNOR2_X1 Check1_CheckInst_0_U137  ( .A(Red_ShiftRowsOutput[1]), .B(
        Red_SignaltoCheck[129]), .ZN(Check1_CheckInst_0_n131 ) );
  XNOR2_X1 Check1_CheckInst_0_U136  ( .A(Red_ShiftRowsOutput[0]), .B(
        Red_SignaltoCheck[128]), .ZN(Check1_CheckInst_0_n132 ) );
  NAND2_X1 Check1_CheckInst_0_U135  ( .A1(Check1_CheckInst_0_n130 ), .A2(
        Check1_CheckInst_0_n129 ), .ZN(Check1_CheckInst_0_n134 ) );
  XNOR2_X1 Check1_CheckInst_0_U134  ( .A(Red_Feedback[13]), .B(
        Red_SignaltoCheck[125]), .ZN(Check1_CheckInst_0_n129 ) );
  XNOR2_X1 Check1_CheckInst_0_U133  ( .A(Red_Feedback[14]), .B(
        Red_SignaltoCheck[126]), .ZN(Check1_CheckInst_0_n130 ) );
  NOR2_X1 Check1_CheckInst_0_U132  ( .A1(Check1_CheckInst_0_n128 ), .A2(
        Check1_CheckInst_0_n127 ), .ZN(Check1_CheckInst_0_n136 ) );
  XOR2_X1 Check1_CheckInst_0_U131  ( .A(Red_ShiftRowsOutput[13]), .B(
        Red_SignaltoCheck[141]), .Z(Check1_CheckInst_0_n127 ) );
  XOR2_X1 Check1_CheckInst_0_U130  ( .A(Red_Feedback[15]), .B(
        Red_SignaltoCheck[127]), .Z(Check1_CheckInst_0_n128 ) );
  NAND2_X1 Check1_CheckInst_0_U129  ( .A1(Check1_CheckInst_0_n126 ), .A2(
        Check1_CheckInst_0_n125 ), .ZN(Check1_CheckInst_0_n138 ) );
  XNOR2_X1 Check1_CheckInst_0_U128  ( .A(Red_ShiftRowsOutput[11]), .B(
        Red_SignaltoCheck[139]), .ZN(Check1_CheckInst_0_n125 ) );
  XNOR2_X1 Check1_CheckInst_0_U127  ( .A(Red_ShiftRowsOutput[14]), .B(
        Red_SignaltoCheck[142]), .ZN(Check1_CheckInst_0_n126 ) );
  NOR2_X1 Check1_CheckInst_0_U126  ( .A1(Check1_CheckInst_0_n124 ), .A2(
        Check1_CheckInst_0_n123 ), .ZN(Check1_CheckInst_0_n284 ) );
  NAND2_X1 Check1_CheckInst_0_U125  ( .A1(Check1_CheckInst_0_n122 ), .A2(
        Check1_CheckInst_0_n121 ), .ZN(Check1_CheckInst_0_n123 ) );
  NOR2_X1 Check1_CheckInst_0_U124  ( .A1(Check1_CheckInst_0_n120 ), .A2(
        Check1_CheckInst_0_n119 ), .ZN(Check1_CheckInst_0_n121 ) );
  NAND2_X1 Check1_CheckInst_0_U123  ( .A1(Check1_CheckInst_0_n118 ), .A2(
        Check1_CheckInst_0_n117 ), .ZN(Check1_CheckInst_0_n119 ) );
  NOR2_X1 Check1_CheckInst_0_U122  ( .A1(Check1_CheckInst_0_n116 ), .A2(
        Check1_CheckInst_0_n115 ), .ZN(Check1_CheckInst_0_n117 ) );
  NAND2_X1 Check1_CheckInst_0_U121  ( .A1(Check1_CheckInst_0_n114 ), .A2(
        Check1_CheckInst_0_n113 ), .ZN(Check1_CheckInst_0_n115 ) );
  NOR2_X1 Check1_CheckInst_0_U120  ( .A1(Check1_CheckInst_0_n112 ), .A2(
        Check1_CheckInst_0_n111 ), .ZN(Check1_CheckInst_0_n113 ) );
  XOR2_X1 Check1_CheckInst_0_U119  ( .A(Red_ShiftRowsOutput[9]), .B(
        Red_SignaltoCheck[137]), .Z(Check1_CheckInst_0_n111 ) );
  XOR2_X1 Check1_CheckInst_0_U118  ( .A(Red_ShiftRowsOutput[12]), .B(
        Red_SignaltoCheck[140]), .Z(Check1_CheckInst_0_n112 ) );
  NOR2_X1 Check1_CheckInst_0_U117  ( .A1(Check1_CheckInst_0_n110 ), .A2(
        Check1_CheckInst_0_n109 ), .ZN(Check1_CheckInst_0_n114 ) );
  XOR2_X1 Check1_CheckInst_0_U116  ( .A(Red_ShiftRowsOutput[7]), .B(
        Red_SignaltoCheck[135]), .Z(Check1_CheckInst_0_n109 ) );
  XOR2_X1 Check1_CheckInst_0_U115  ( .A(Red_ShiftRowsOutput[10]), .B(
        Red_SignaltoCheck[138]), .Z(Check1_CheckInst_0_n110 ) );
  NAND2_X1 Check1_CheckInst_0_U114  ( .A1(Check1_CheckInst_0_n108 ), .A2(
        Check1_CheckInst_0_n107 ), .ZN(Check1_CheckInst_0_n116 ) );
  XNOR2_X1 Check1_CheckInst_0_U113  ( .A(Red_ShiftRowsOutput[8]), .B(
        Red_SignaltoCheck[136]), .ZN(Check1_CheckInst_0_n107 ) );
  XNOR2_X1 Check1_CheckInst_0_U112  ( .A(Red_ShiftRowsOutput[6]), .B(
        Red_SignaltoCheck[134]), .ZN(Check1_CheckInst_0_n108 ) );
  NOR2_X1 Check1_CheckInst_0_U111  ( .A1(Check1_CheckInst_0_n106 ), .A2(
        Check1_CheckInst_0_n105 ), .ZN(Check1_CheckInst_0_n118 ) );
  XOR2_X1 Check1_CheckInst_0_U110  ( .A(Red_Feedback[3]), .B(
        Red_SignaltoCheck[115]), .Z(Check1_CheckInst_0_n105 ) );
  XOR2_X1 Check1_CheckInst_0_U109  ( .A(Red_Feedback[2]), .B(
        Red_SignaltoCheck[114]), .Z(Check1_CheckInst_0_n106 ) );
  NAND2_X1 Check1_CheckInst_0_U108  ( .A1(Check1_CheckInst_0_n104 ), .A2(
        Check1_CheckInst_0_n103 ), .ZN(Check1_CheckInst_0_n120 ) );
  NOR2_X1 Check1_CheckInst_0_U107  ( .A1(Check1_CheckInst_0_n102 ), .A2(
        Check1_CheckInst_0_n101 ), .ZN(Check1_CheckInst_0_n103 ) );
  NAND2_X1 Check1_CheckInst_0_U106  ( .A1(Check1_CheckInst_0_n100 ), .A2(
        Check1_CheckInst_0_n99 ), .ZN(Check1_CheckInst_0_n101 ) );
  NOR2_X1 Check1_CheckInst_0_U105  ( .A1(Check1_CheckInst_0_n98 ), .A2(
        Check1_CheckInst_0_n97 ), .ZN(Check1_CheckInst_0_n99 ) );
  XOR2_X1 Check1_CheckInst_0_U104  ( .A(Red_Feedback[1]), .B(
        Red_SignaltoCheck[113]), .Z(Check1_CheckInst_0_n97 ) );
  XOR2_X1 Check1_CheckInst_0_U103  ( .A(Red_Feedback[0]), .B(
        Red_SignaltoCheck[112]), .Z(Check1_CheckInst_0_n98 ) );
  NOR2_X1 Check1_CheckInst_0_U102  ( .A1(Check1_CheckInst_0_n96 ), .A2(
        Check1_CheckInst_0_n95 ), .ZN(Check1_CheckInst_0_n100 ) );
  XOR2_X1 Check1_CheckInst_0_U101  ( .A(Red_SubCellInput[15]), .B(
        Red_SignaltoCheck[111]), .Z(Check1_CheckInst_0_n95 ) );
  XOR2_X1 Check1_CheckInst_0_U100  ( .A(Red_SubCellInput[14]), .B(
        Red_SignaltoCheck[110]), .Z(Check1_CheckInst_0_n96 ) );
  NAND2_X1 Check1_CheckInst_0_U99  ( .A1(Check1_CheckInst_0_n94 ), .A2(
        Check1_CheckInst_0_n93 ), .ZN(Check1_CheckInst_0_n102 ) );
  XNOR2_X1 Check1_CheckInst_0_U98  ( .A(Red_SubCellInput[11]), .B(
        Red_SignaltoCheck[107]), .ZN(Check1_CheckInst_0_n93 ) );
  XNOR2_X1 Check1_CheckInst_0_U97  ( .A(Red_SubCellInput[12]), .B(
        Red_SignaltoCheck[108]), .ZN(Check1_CheckInst_0_n94 ) );
  NOR2_X1 Check1_CheckInst_0_U96  ( .A1(Check1_CheckInst_0_n92 ), .A2(
        Check1_CheckInst_0_n91 ), .ZN(Check1_CheckInst_0_n104 ) );
  XOR2_X1 Check1_CheckInst_0_U95  ( .A(Red_Feedback[11]), .B(
        Red_SignaltoCheck[123]), .Z(Check1_CheckInst_0_n91 ) );
  XOR2_X1 Check1_CheckInst_0_U94  ( .A(Red_SubCellInput[13]), .B(
        Red_SignaltoCheck[109]), .Z(Check1_CheckInst_0_n92 ) );
  NOR2_X1 Check1_CheckInst_0_U93  ( .A1(Check1_CheckInst_0_n90 ), .A2(
        Check1_CheckInst_0_n89 ), .ZN(Check1_CheckInst_0_n122 ) );
  NAND2_X1 Check1_CheckInst_0_U92  ( .A1(Check1_CheckInst_0_n88 ), .A2(
        Check1_CheckInst_0_n87 ), .ZN(Check1_CheckInst_0_n89 ) );
  NOR2_X1 Check1_CheckInst_0_U91  ( .A1(Check1_CheckInst_0_n86 ), .A2(
        Check1_CheckInst_0_n85 ), .ZN(Check1_CheckInst_0_n87 ) );
  NAND2_X1 Check1_CheckInst_0_U90  ( .A1(Check1_CheckInst_0_n84 ), .A2(
        Check1_CheckInst_0_n83 ), .ZN(Check1_CheckInst_0_n85 ) );
  XNOR2_X1 Check1_CheckInst_0_U89  ( .A(Red_Feedback[9]), .B(
        Red_SignaltoCheck[121]), .ZN(Check1_CheckInst_0_n83 ) );
  XNOR2_X1 Check1_CheckInst_0_U88  ( .A(Red_Feedback[12]), .B(
        Red_SignaltoCheck[124]), .ZN(Check1_CheckInst_0_n84 ) );
  NAND2_X1 Check1_CheckInst_0_U87  ( .A1(Check1_CheckInst_0_n82 ), .A2(
        Check1_CheckInst_0_n81 ), .ZN(Check1_CheckInst_0_n86 ) );
  XNOR2_X1 Check1_CheckInst_0_U86  ( .A(Red_Feedback[7]), .B(
        Red_SignaltoCheck[119]), .ZN(Check1_CheckInst_0_n81 ) );
  XNOR2_X1 Check1_CheckInst_0_U85  ( .A(Red_Feedback[10]), .B(
        Red_SignaltoCheck[122]), .ZN(Check1_CheckInst_0_n82 ) );
  NOR2_X1 Check1_CheckInst_0_U84  ( .A1(Check1_CheckInst_0_n80 ), .A2(
        Check1_CheckInst_0_n79 ), .ZN(Check1_CheckInst_0_n88 ) );
  XOR2_X1 Check1_CheckInst_0_U83  ( .A(Red_Feedback[5]), .B(
        Red_SignaltoCheck[117]), .Z(Check1_CheckInst_0_n79 ) );
  XOR2_X1 Check1_CheckInst_0_U82  ( .A(Red_Feedback[8]), .B(
        Red_SignaltoCheck[120]), .Z(Check1_CheckInst_0_n80 ) );
  NAND2_X1 Check1_CheckInst_0_U81  ( .A1(Check1_CheckInst_0_n78 ), .A2(
        Check1_CheckInst_0_n77 ), .ZN(Check1_CheckInst_0_n90 ) );
  XNOR2_X1 Check1_CheckInst_0_U80  ( .A(Red_Feedback[6]), .B(
        Red_SignaltoCheck[118]), .ZN(Check1_CheckInst_0_n77 ) );
  XNOR2_X1 Check1_CheckInst_0_U79  ( .A(Red_Feedback[4]), .B(
        Red_SignaltoCheck[116]), .ZN(Check1_CheckInst_0_n78 ) );
  NAND2_X1 Check1_CheckInst_0_U78  ( .A1(Check1_CheckInst_0_n76 ), .A2(
        Check1_CheckInst_0_n75 ), .ZN(Check1_CheckInst_0_n124 ) );
  NOR2_X1 Check1_CheckInst_0_U77  ( .A1(Check1_CheckInst_0_n74 ), .A2(
        Check1_CheckInst_0_n73 ), .ZN(Check1_CheckInst_0_n75 ) );
  NAND2_X1 Check1_CheckInst_0_U76  ( .A1(Check1_CheckInst_0_n72 ), .A2(
        Check1_CheckInst_0_n71 ), .ZN(Check1_CheckInst_0_n73 ) );
  NOR2_X1 Check1_CheckInst_0_U75  ( .A1(Check1_CheckInst_0_n70 ), .A2(
        Check1_CheckInst_0_n69 ), .ZN(Check1_CheckInst_0_n71 ) );
  XOR2_X1 Check1_CheckInst_0_U74  ( .A(Red_Feedback3[9]), .B(
        Red_SignaltoCheck[25]), .Z(Check1_CheckInst_0_n69 ) );
  XOR2_X1 Check1_CheckInst_0_U73  ( .A(Red_Feedback3[8]), .B(
        Red_SignaltoCheck[24]), .Z(Check1_CheckInst_0_n70 ) );
  NOR2_X1 Check1_CheckInst_0_U72  ( .A1(Check1_CheckInst_0_n68 ), .A2(
        Check1_CheckInst_0_n67 ), .ZN(Check1_CheckInst_0_n72 ) );
  XOR2_X1 Check1_CheckInst_0_U71  ( .A(Red_Feedback3[7]), .B(
        Red_SignaltoCheck[23]), .Z(Check1_CheckInst_0_n67 ) );
  XOR2_X1 Check1_CheckInst_0_U70  ( .A(Red_Feedback3[6]), .B(
        Red_SignaltoCheck[22]), .Z(Check1_CheckInst_0_n68 ) );
  NAND2_X1 Check1_CheckInst_0_U69  ( .A1(Check1_CheckInst_0_n66 ), .A2(
        Check1_CheckInst_0_n65 ), .ZN(Check1_CheckInst_0_n74 ) );
  XNOR2_X1 Check1_CheckInst_0_U68  ( .A(Red_Feedback3[5]), .B(
        Red_SignaltoCheck[21]), .ZN(Check1_CheckInst_0_n65 ) );
  XNOR2_X1 Check1_CheckInst_0_U67  ( .A(Red_Feedback3[4]), .B(
        Red_SignaltoCheck[20]), .ZN(Check1_CheckInst_0_n66 ) );
  NOR2_X1 Check1_CheckInst_0_U66  ( .A1(Check1_CheckInst_0_n64 ), .A2(
        Check1_CheckInst_0_n63 ), .ZN(Check1_CheckInst_0_n76 ) );
  XOR2_X1 Check1_CheckInst_0_U65  ( .A(Red_Feedback3[1]), .B(
        Red_SignaltoCheck[17]), .Z(Check1_CheckInst_0_n63 ) );
  XOR2_X1 Check1_CheckInst_0_U64  ( .A(Red_Feedback3[2]), .B(
        Red_SignaltoCheck[18]), .Z(Check1_CheckInst_0_n64 ) );
  NAND2_X1 Check1_CheckInst_0_U63  ( .A1(Check1_CheckInst_0_n62 ), .A2(
        Check1_CheckInst_0_n61 ), .ZN(Check1_CheckInst_0_n286 ) );
  NOR2_X1 Check1_CheckInst_0_U62  ( .A1(Check1_CheckInst_0_n60 ), .A2(
        Check1_CheckInst_0_n59 ), .ZN(Check1_CheckInst_0_n61 ) );
  NAND2_X1 Check1_CheckInst_0_U61  ( .A1(Check1_CheckInst_0_n58 ), .A2(
        Check1_CheckInst_0_n57 ), .ZN(Check1_CheckInst_0_n59 ) );
  NOR2_X1 Check1_CheckInst_0_U60  ( .A1(Check1_CheckInst_0_n56 ), .A2(
        Check1_CheckInst_0_n55 ), .ZN(Check1_CheckInst_0_n57 ) );
  NAND2_X1 Check1_CheckInst_0_U59  ( .A1(Check1_CheckInst_0_n54 ), .A2(
        Check1_CheckInst_0_n53 ), .ZN(Check1_CheckInst_0_n55 ) );
  NOR2_X1 Check1_CheckInst_0_U58  ( .A1(Check1_CheckInst_0_n52 ), .A2(
        Check1_CheckInst_0_n51 ), .ZN(Check1_CheckInst_0_n53 ) );
  NAND2_X1 Check1_CheckInst_0_U57  ( .A1(Check1_CheckInst_0_n50 ), .A2(
        Check1_CheckInst_0_n49 ), .ZN(Check1_CheckInst_0_n51 ) );
  XNOR2_X1 Check1_CheckInst_0_U56  ( .A(Red_ShiftRowsOutput3[1]), .B(
        Red_SignaltoCheck[33]), .ZN(Check1_CheckInst_0_n49 ) );
  XNOR2_X1 Check1_CheckInst_0_U55  ( .A(Red_Feedback3[3]), .B(
        Red_SignaltoCheck[19]), .ZN(Check1_CheckInst_0_n50 ) );
  NAND2_X1 Check1_CheckInst_0_U54  ( .A1(Check1_CheckInst_0_n48 ), .A2(
        Check1_CheckInst_0_n47 ), .ZN(Check1_CheckInst_0_n52 ) );
  XNOR2_X1 Check1_CheckInst_0_U53  ( .A(Red_Feedback3[15]), .B(
        Red_SignaltoCheck[31]), .ZN(Check1_CheckInst_0_n47 ) );
  XNOR2_X1 Check1_CheckInst_0_U52  ( .A(Red_ShiftRowsOutput3[2]), .B(
        Red_SignaltoCheck[34]), .ZN(Check1_CheckInst_0_n48 ) );
  NOR2_X1 Check1_CheckInst_0_U51  ( .A1(Check1_CheckInst_0_n46 ), .A2(
        Check1_CheckInst_0_n45 ), .ZN(Check1_CheckInst_0_n54 ) );
  XOR2_X1 Check1_CheckInst_0_U50  ( .A(Red_Feedback3[13]), .B(
        Red_SignaltoCheck[29]), .Z(Check1_CheckInst_0_n45 ) );
  XOR2_X1 Check1_CheckInst_0_U49  ( .A(Red_ShiftRowsOutput3[0]), .B(
        Red_SignaltoCheck[32]), .Z(Check1_CheckInst_0_n46 ) );
  NAND2_X1 Check1_CheckInst_0_U48  ( .A1(Check1_CheckInst_0_n44 ), .A2(
        Check1_CheckInst_0_n43 ), .ZN(Check1_CheckInst_0_n56 ) );
  XNOR2_X1 Check1_CheckInst_0_U47  ( .A(Red_Feedback3[11]), .B(
        Red_SignaltoCheck[27]), .ZN(Check1_CheckInst_0_n43 ) );
  XNOR2_X1 Check1_CheckInst_0_U46  ( .A(Red_Feedback3[14]), .B(
        Red_SignaltoCheck[30]), .ZN(Check1_CheckInst_0_n44 ) );
  NOR2_X1 Check1_CheckInst_0_U45  ( .A1(Check1_CheckInst_0_n42 ), .A2(
        Check1_CheckInst_0_n41 ), .ZN(Check1_CheckInst_0_n58 ) );
  NAND2_X1 Check1_CheckInst_0_U44  ( .A1(Check1_CheckInst_0_n40 ), .A2(
        Check1_CheckInst_0_n39 ), .ZN(Check1_CheckInst_0_n41 ) );
  NOR2_X1 Check1_CheckInst_0_U43  ( .A1(Check1_CheckInst_0_n38 ), .A2(
        Check1_CheckInst_0_n37 ), .ZN(Check1_CheckInst_0_n39 ) );
  NAND2_X1 Check1_CheckInst_0_U42  ( .A1(Check1_CheckInst_0_n36 ), .A2(
        Check1_CheckInst_0_n35 ), .ZN(Check1_CheckInst_0_n37 ) );
  XNOR2_X1 Check1_CheckInst_0_U41  ( .A(Red_Feedback3[12]), .B(
        Red_SignaltoCheck[28]), .ZN(Check1_CheckInst_0_n35 ) );
  XNOR2_X1 Check1_CheckInst_0_U40  ( .A(Red_Feedback3[10]), .B(
        Red_SignaltoCheck[26]), .ZN(Check1_CheckInst_0_n36 ) );
  NAND2_X1 Check1_CheckInst_0_U39  ( .A1(Check1_CheckInst_0_n34 ), .A2(
        Check1_CheckInst_0_n33 ), .ZN(Check1_CheckInst_0_n38 ) );
  XNOR2_X1 Check1_CheckInst_0_U38  ( .A(Red_AddRoundKeyOutput[7]), .B(
        Red_SignaltoCheck[7]), .ZN(Check1_CheckInst_0_n33 ) );
  XNOR2_X1 Check1_CheckInst_0_U37  ( .A(Red_AddRoundKeyOutput[6]), .B(
        Red_SignaltoCheck[6]), .ZN(Check1_CheckInst_0_n34 ) );
  NOR2_X1 Check1_CheckInst_0_U36  ( .A1(Check1_CheckInst_0_n32 ), .A2(
        Check1_CheckInst_0_n31 ), .ZN(Check1_CheckInst_0_n40 ) );
  XOR2_X1 Check1_CheckInst_0_U35  ( .A(Red_AddRoundKeyOutput[5]), .B(
        Red_SignaltoCheck[5]), .Z(Check1_CheckInst_0_n31 ) );
  XOR2_X1 Check1_CheckInst_0_U34  ( .A(Red_AddRoundKeyOutput[4]), .B(
        Red_SignaltoCheck[4]), .Z(Check1_CheckInst_0_n32 ) );
  NAND2_X1 Check1_CheckInst_0_U33  ( .A1(Check1_CheckInst_0_n30 ), .A2(
        Check1_CheckInst_0_n29 ), .ZN(Check1_CheckInst_0_n42 ) );
  XNOR2_X1 Check1_CheckInst_0_U32  ( .A(Red_AddRoundKeyOutput[3]), .B(
        Red_SignaltoCheck[3]), .ZN(Check1_CheckInst_0_n29 ) );
  XNOR2_X1 Check1_CheckInst_0_U31  ( .A(Red_AddRoundKeyOutput[2]), .B(
        Red_SignaltoCheck[2]), .ZN(Check1_CheckInst_0_n30 ) );
  NAND2_X1 Check1_CheckInst_0_U30  ( .A1(Check1_CheckInst_0_n28 ), .A2(
        Check1_CheckInst_0_n27 ), .ZN(Check1_CheckInst_0_n60 ) );
  NOR2_X1 Check1_CheckInst_0_U29  ( .A1(Check1_CheckInst_0_n26 ), .A2(
        Check1_CheckInst_0_n25 ), .ZN(Check1_CheckInst_0_n27 ) );
  NAND2_X1 Check1_CheckInst_0_U28  ( .A1(Check1_CheckInst_0_n24 ), .A2(
        Check1_CheckInst_0_n23 ), .ZN(Check1_CheckInst_0_n25 ) );
  NOR2_X1 Check1_CheckInst_0_U27  ( .A1(Check1_CheckInst_0_n22 ), .A2(
        Check1_CheckInst_0_n21 ), .ZN(Check1_CheckInst_0_n23 ) );
  XOR2_X1 Check1_CheckInst_0_U26  ( .A(Red_SignaltoCheck[1]), .B(
        Red_AddRoundKeyOutput[1]), .Z(Check1_CheckInst_0_n21 ) );
  XOR2_X1 Check1_CheckInst_0_U25  ( .A(Red_AddRoundKeyOutput[0]), .B(
        Red_SignaltoCheck[0]), .Z(Check1_CheckInst_0_n22 ) );
  NOR2_X1 Check1_CheckInst_0_U24  ( .A1(Check1_CheckInst_0_n20 ), .A2(
        Check1_CheckInst_0_n19 ), .ZN(Check1_CheckInst_0_n24 ) );
  XOR2_X1 Check1_CheckInst_0_U23  ( .A(Red_AddRoundKeyOutput[15]), .B(
        Red_SignaltoCheck[15]), .Z(Check1_CheckInst_0_n19 ) );
  XOR2_X1 Check1_CheckInst_0_U22  ( .A(Red_ShiftRowsOutput[15]), .B(
        Red_SignaltoCheck[143]), .Z(Check1_CheckInst_0_n20 ) );
  NAND2_X1 Check1_CheckInst_0_U21  ( .A1(Check1_CheckInst_0_n18 ), .A2(
        Check1_CheckInst_0_n17 ), .ZN(Check1_CheckInst_0_n26 ) );
  XNOR2_X1 Check1_CheckInst_0_U20  ( .A(Red_AddRoundKeyOutput[13]), .B(
        Red_SignaltoCheck[13]), .ZN(Check1_CheckInst_0_n17 ) );
  XNOR2_X1 Check1_CheckInst_0_U19  ( .A(Red_Feedback3[0]), .B(
        Red_SignaltoCheck[16]), .ZN(Check1_CheckInst_0_n18 ) );
  NOR2_X1 Check1_CheckInst_0_U18  ( .A1(Check1_CheckInst_0_n16 ), .A2(
        Check1_CheckInst_0_n15 ), .ZN(Check1_CheckInst_0_n28 ) );
  XOR2_X1 Check1_CheckInst_0_U17  ( .A(Red_AddRoundKeyOutput[11]), .B(
        Red_SignaltoCheck[11]), .Z(Check1_CheckInst_0_n15 ) );
  XOR2_X1 Check1_CheckInst_0_U16  ( .A(Red_AddRoundKeyOutput[14]), .B(
        Red_SignaltoCheck[14]), .Z(Check1_CheckInst_0_n16 ) );
  NOR2_X1 Check1_CheckInst_0_U15  ( .A1(Check1_CheckInst_0_n14 ), .A2(
        Check1_CheckInst_0_n13 ), .ZN(Check1_CheckInst_0_n62 ) );
  NAND2_X1 Check1_CheckInst_0_U14  ( .A1(Check1_CheckInst_0_n12 ), .A2(
        Check1_CheckInst_0_n11 ), .ZN(Check1_CheckInst_0_n13 ) );
  NOR2_X1 Check1_CheckInst_0_U13  ( .A1(Check1_CheckInst_0_n10 ), .A2(
        Check1_CheckInst_0_n9 ), .ZN(Check1_CheckInst_0_n11 ) );
  NAND2_X1 Check1_CheckInst_0_U12  ( .A1(Check1_CheckInst_0_n8 ), .A2(
        Check1_CheckInst_0_n7 ), .ZN(Check1_CheckInst_0_n9 ) );
  XNOR2_X1 Check1_CheckInst_0_U11  ( .A(Red_AddRoundKeyOutput[9]), .B(
        Red_SignaltoCheck[9]), .ZN(Check1_CheckInst_0_n7 ) );
  XNOR2_X1 Check1_CheckInst_0_U10  ( .A(Red_AddRoundKeyOutput[12]), .B(
        Red_SignaltoCheck[12]), .ZN(Check1_CheckInst_0_n8 ) );
  NAND2_X1 Check1_CheckInst_0_U9  ( .A1(Check1_CheckInst_0_n6 ), .A2(
        Check1_CheckInst_0_n5 ), .ZN(Check1_CheckInst_0_n10 ) );
  XNOR2_X1 Check1_CheckInst_0_U8  ( .A(Red_AddRoundKeyOutput[10]), .B(
        Red_SignaltoCheck[10]), .ZN(Check1_CheckInst_0_n5 ) );
  XNOR2_X1 Check1_CheckInst_0_U7  ( .A(Red_AddRoundKeyOutput[8]), .B(
        Red_SignaltoCheck[8]), .ZN(Check1_CheckInst_0_n6 ) );
  NOR2_X1 Check1_CheckInst_0_U6  ( .A1(Check1_CheckInst_0_n4 ), .A2(
        Check1_CheckInst_0_n3 ), .ZN(Check1_CheckInst_0_n12 ) );
  XOR2_X1 Check1_CheckInst_0_U5  ( .A(Red_SubCellInput2[13]), .B(
        Red_SignaltoCheck[61]), .Z(Check1_CheckInst_0_n3 ) );
  XOR2_X1 Check1_CheckInst_0_U4  ( .A(Red_SubCellInput2[12]), .B(
        Red_SignaltoCheck[60]), .Z(Check1_CheckInst_0_n4 ) );
  NAND2_X1 Check1_CheckInst_0_U3  ( .A1(Check1_CheckInst_0_n2 ), .A2(
        Check1_CheckInst_0_n1 ), .ZN(Check1_CheckInst_0_n14 ) );
  XNOR2_X1 Check1_CheckInst_0_U2  ( .A(Red_SubCellInput2[11]), .B(
        Red_SignaltoCheck[59]), .ZN(Check1_CheckInst_0_n1 ) );
  XNOR2_X1 Check1_CheckInst_0_U1  ( .A(Red_SubCellInput2[10]), .B(
        Red_SignaltoCheck[58]), .ZN(Check1_CheckInst_0_n2 ) );
endmodule

