module Cipher ( clk, rst, EncDec, Input, Key, Tweak, Output );
  input [63:0] Input;
  input [127:0] Key;
  output [63:0] Output;
  (* FIRMER="clock" *)input clk;
  (* FIRMER="control" *)input rst;
  wire   MCInst_XOR_r0_Inst_0_n3 , MCInst_XOR_r0_Inst_1_n3 ,
         MCInst_XOR_r0_Inst_2_n3 , MCInst_XOR_r0_Inst_3_n3 ,
         MCInst_XOR_r0_Inst_4_n3 , MCInst_XOR_r0_Inst_5_n3 ,
         MCInst_XOR_r0_Inst_6_n3 , MCInst_XOR_r0_Inst_7_n3 ,
         MCInst_XOR_r0_Inst_8_n3 , MCInst_XOR_r0_Inst_9_n3 ,
         MCInst_XOR_r0_Inst_10_n3 , MCInst_XOR_r0_Inst_11_n3 ,
         MCInst_XOR_r0_Inst_12_n3 , MCInst_XOR_r0_Inst_13_n3 ,
         MCInst_XOR_r0_Inst_14_n3 , MCInst_XOR_r0_Inst_15_n3 ,
         SubCellInst_LFInst_0_n36 , SubCellInst_LFInst_0_n35 ,
         SubCellInst_LFInst_0_n34 , SubCellInst_LFInst_0_n33 ,
         SubCellInst_LFInst_0_n32 , SubCellInst_LFInst_0_n31 ,
         SubCellInst_LFInst_0_n30 , SubCellInst_LFInst_0_n29 ,
         SubCellInst_LFInst_0_n28 , SubCellInst_LFInst_0_n27 ,
         SubCellInst_LFInst_0_n26 , SubCellInst_LFInst_0_n25 ,
         SubCellInst_LFInst_0_n24 , SubCellInst_LFInst_0_n23 ,
         SubCellInst_LFInst_0_n22 , SubCellInst_LFInst_1_n36 ,
         SubCellInst_LFInst_1_n35 , SubCellInst_LFInst_1_n34 ,
         SubCellInst_LFInst_1_n33 , SubCellInst_LFInst_1_n32 ,
         SubCellInst_LFInst_1_n31 , SubCellInst_LFInst_1_n30 ,
         SubCellInst_LFInst_1_n29 , SubCellInst_LFInst_1_n28 ,
         SubCellInst_LFInst_1_n27 , SubCellInst_LFInst_1_n26 ,
         SubCellInst_LFInst_1_n25 , SubCellInst_LFInst_1_n24 ,
         SubCellInst_LFInst_1_n23 , SubCellInst_LFInst_1_n22 ,
         SubCellInst_LFInst_2_n36 , SubCellInst_LFInst_2_n35 ,
         SubCellInst_LFInst_2_n34 , SubCellInst_LFInst_2_n33 ,
         SubCellInst_LFInst_2_n32 , SubCellInst_LFInst_2_n31 ,
         SubCellInst_LFInst_2_n30 , SubCellInst_LFInst_2_n29 ,
         SubCellInst_LFInst_2_n28 , SubCellInst_LFInst_2_n27 ,
         SubCellInst_LFInst_2_n26 , SubCellInst_LFInst_2_n25 ,
         SubCellInst_LFInst_2_n24 , SubCellInst_LFInst_2_n23 ,
         SubCellInst_LFInst_2_n22 , SubCellInst_LFInst_3_n36 ,
         SubCellInst_LFInst_3_n35 , SubCellInst_LFInst_3_n34 ,
         SubCellInst_LFInst_3_n33 , SubCellInst_LFInst_3_n32 ,
         SubCellInst_LFInst_3_n31 , SubCellInst_LFInst_3_n30 ,
         SubCellInst_LFInst_3_n29 , SubCellInst_LFInst_3_n28 ,
         SubCellInst_LFInst_3_n27 , SubCellInst_LFInst_3_n26 ,
         SubCellInst_LFInst_3_n25 , SubCellInst_LFInst_3_n24 ,
         SubCellInst_LFInst_3_n23 , SubCellInst_LFInst_3_n22 ,
         SubCellInst_LFInst_4_n36 , SubCellInst_LFInst_4_n35 ,
         SubCellInst_LFInst_4_n34 , SubCellInst_LFInst_4_n33 ,
         SubCellInst_LFInst_4_n32 , SubCellInst_LFInst_4_n31 ,
         SubCellInst_LFInst_4_n30 , SubCellInst_LFInst_4_n29 ,
         SubCellInst_LFInst_4_n28 , SubCellInst_LFInst_4_n27 ,
         SubCellInst_LFInst_4_n26 , SubCellInst_LFInst_4_n25 ,
         SubCellInst_LFInst_4_n24 , SubCellInst_LFInst_4_n23 ,
         SubCellInst_LFInst_4_n22 , SubCellInst_LFInst_5_n36 ,
         SubCellInst_LFInst_5_n35 , SubCellInst_LFInst_5_n34 ,
         SubCellInst_LFInst_5_n33 , SubCellInst_LFInst_5_n32 ,
         SubCellInst_LFInst_5_n31 , SubCellInst_LFInst_5_n30 ,
         SubCellInst_LFInst_5_n29 , SubCellInst_LFInst_5_n28 ,
         SubCellInst_LFInst_5_n27 , SubCellInst_LFInst_5_n26 ,
         SubCellInst_LFInst_5_n25 , SubCellInst_LFInst_5_n24 ,
         SubCellInst_LFInst_5_n23 , SubCellInst_LFInst_5_n22 ,
         SubCellInst_LFInst_6_n36 , SubCellInst_LFInst_6_n35 ,
         SubCellInst_LFInst_6_n34 , SubCellInst_LFInst_6_n33 ,
         SubCellInst_LFInst_6_n32 , SubCellInst_LFInst_6_n31 ,
         SubCellInst_LFInst_6_n30 , SubCellInst_LFInst_6_n29 ,
         SubCellInst_LFInst_6_n28 , SubCellInst_LFInst_6_n27 ,
         SubCellInst_LFInst_6_n26 , SubCellInst_LFInst_6_n25 ,
         SubCellInst_LFInst_6_n24 , SubCellInst_LFInst_6_n23 ,
         SubCellInst_LFInst_6_n22 , SubCellInst_LFInst_7_n36 ,
         SubCellInst_LFInst_7_n35 , SubCellInst_LFInst_7_n34 ,
         SubCellInst_LFInst_7_n33 , SubCellInst_LFInst_7_n32 ,
         SubCellInst_LFInst_7_n31 , SubCellInst_LFInst_7_n30 ,
         SubCellInst_LFInst_7_n29 , SubCellInst_LFInst_7_n28 ,
         SubCellInst_LFInst_7_n27 , SubCellInst_LFInst_7_n26 ,
         SubCellInst_LFInst_7_n25 , SubCellInst_LFInst_7_n24 ,
         SubCellInst_LFInst_7_n23 , SubCellInst_LFInst_7_n22 ,
         SubCellInst_LFInst_8_n36 , SubCellInst_LFInst_8_n35 ,
         SubCellInst_LFInst_8_n34 , SubCellInst_LFInst_8_n33 ,
         SubCellInst_LFInst_8_n32 , SubCellInst_LFInst_8_n31 ,
         SubCellInst_LFInst_8_n30 , SubCellInst_LFInst_8_n29 ,
         SubCellInst_LFInst_8_n28 , SubCellInst_LFInst_8_n27 ,
         SubCellInst_LFInst_8_n26 , SubCellInst_LFInst_8_n25 ,
         SubCellInst_LFInst_8_n24 , SubCellInst_LFInst_8_n23 ,
         SubCellInst_LFInst_8_n22 , SubCellInst_LFInst_9_n36 ,
         SubCellInst_LFInst_9_n35 , SubCellInst_LFInst_9_n34 ,
         SubCellInst_LFInst_9_n33 , SubCellInst_LFInst_9_n32 ,
         SubCellInst_LFInst_9_n31 , SubCellInst_LFInst_9_n30 ,
         SubCellInst_LFInst_9_n29 , SubCellInst_LFInst_9_n28 ,
         SubCellInst_LFInst_9_n27 , SubCellInst_LFInst_9_n26 ,
         SubCellInst_LFInst_9_n25 , SubCellInst_LFInst_9_n24 ,
         SubCellInst_LFInst_9_n23 , SubCellInst_LFInst_9_n22 ,
         SubCellInst_LFInst_10_n36 , SubCellInst_LFInst_10_n35 ,
         SubCellInst_LFInst_10_n34 , SubCellInst_LFInst_10_n33 ,
         SubCellInst_LFInst_10_n32 , SubCellInst_LFInst_10_n31 ,
         SubCellInst_LFInst_10_n30 , SubCellInst_LFInst_10_n29 ,
         SubCellInst_LFInst_10_n28 , SubCellInst_LFInst_10_n27 ,
         SubCellInst_LFInst_10_n26 , SubCellInst_LFInst_10_n25 ,
         SubCellInst_LFInst_10_n24 , SubCellInst_LFInst_10_n23 ,
         SubCellInst_LFInst_10_n22 , SubCellInst_LFInst_11_n36 ,
         SubCellInst_LFInst_11_n35 , SubCellInst_LFInst_11_n34 ,
         SubCellInst_LFInst_11_n33 , SubCellInst_LFInst_11_n32 ,
         SubCellInst_LFInst_11_n31 , SubCellInst_LFInst_11_n30 ,
         SubCellInst_LFInst_11_n29 , SubCellInst_LFInst_11_n28 ,
         SubCellInst_LFInst_11_n27 , SubCellInst_LFInst_11_n26 ,
         SubCellInst_LFInst_11_n25 , SubCellInst_LFInst_11_n24 ,
         SubCellInst_LFInst_11_n23 , SubCellInst_LFInst_11_n22 ,
         SubCellInst_LFInst_12_n36 , SubCellInst_LFInst_12_n35 ,
         SubCellInst_LFInst_12_n34 , SubCellInst_LFInst_12_n33 ,
         SubCellInst_LFInst_12_n32 , SubCellInst_LFInst_12_n31 ,
         SubCellInst_LFInst_12_n30 , SubCellInst_LFInst_12_n29 ,
         SubCellInst_LFInst_12_n28 , SubCellInst_LFInst_12_n27 ,
         SubCellInst_LFInst_12_n26 , SubCellInst_LFInst_12_n25 ,
         SubCellInst_LFInst_12_n24 , SubCellInst_LFInst_12_n23 ,
         SubCellInst_LFInst_12_n22 , SubCellInst_LFInst_13_n36 ,
         SubCellInst_LFInst_13_n35 , SubCellInst_LFInst_13_n34 ,
         SubCellInst_LFInst_13_n33 , SubCellInst_LFInst_13_n32 ,
         SubCellInst_LFInst_13_n31 , SubCellInst_LFInst_13_n30 ,
         SubCellInst_LFInst_13_n29 , SubCellInst_LFInst_13_n28 ,
         SubCellInst_LFInst_13_n27 , SubCellInst_LFInst_13_n26 ,
         SubCellInst_LFInst_13_n25 , SubCellInst_LFInst_13_n24 ,
         SubCellInst_LFInst_13_n23 , SubCellInst_LFInst_13_n22 ,
         SubCellInst_LFInst_14_n36 , SubCellInst_LFInst_14_n35 ,
         SubCellInst_LFInst_14_n34 , SubCellInst_LFInst_14_n33 ,
         SubCellInst_LFInst_14_n32 , SubCellInst_LFInst_14_n31 ,
         SubCellInst_LFInst_14_n30 , SubCellInst_LFInst_14_n29 ,
         SubCellInst_LFInst_14_n28 , SubCellInst_LFInst_14_n27 ,
         SubCellInst_LFInst_14_n26 , SubCellInst_LFInst_14_n25 ,
         SubCellInst_LFInst_14_n24 , SubCellInst_LFInst_14_n23 ,
         SubCellInst_LFInst_14_n22 , SubCellInst_LFInst_15_n36 ,
         SubCellInst_LFInst_15_n35 , SubCellInst_LFInst_15_n34 ,
         SubCellInst_LFInst_15_n33 , SubCellInst_LFInst_15_n32 ,
         SubCellInst_LFInst_15_n31 , SubCellInst_LFInst_15_n30 ,
         SubCellInst_LFInst_15_n29 , SubCellInst_LFInst_15_n28 ,
         SubCellInst_LFInst_15_n27 , SubCellInst_LFInst_15_n26 ,
         SubCellInst_LFInst_15_n25 , SubCellInst_LFInst_15_n24 ,
         SubCellInst_LFInst_15_n23 , SubCellInst_LFInst_15_n22 ,
         MCInst2_XOR_r0_Inst_0_n3 , MCInst2_XOR_r0_Inst_1_n3 ,
         MCInst2_XOR_r0_Inst_2_n3 , MCInst2_XOR_r0_Inst_3_n3 ,
         MCInst2_XOR_r0_Inst_4_n3 , MCInst2_XOR_r0_Inst_5_n3 ,
         MCInst2_XOR_r0_Inst_6_n3 , MCInst2_XOR_r0_Inst_7_n3 ,
         MCInst2_XOR_r0_Inst_8_n3 , MCInst2_XOR_r0_Inst_9_n3 ,
         MCInst2_XOR_r0_Inst_10_n3 , MCInst2_XOR_r0_Inst_11_n3 ,
         MCInst2_XOR_r0_Inst_12_n3 , MCInst2_XOR_r0_Inst_13_n3 ,
         MCInst2_XOR_r0_Inst_14_n3 , MCInst2_XOR_r0_Inst_15_n3 ,
         SubCellInst2_LFInst_0_n36 , SubCellInst2_LFInst_0_n35 ,
         SubCellInst2_LFInst_0_n34 , SubCellInst2_LFInst_0_n33 ,
         SubCellInst2_LFInst_0_n32 , SubCellInst2_LFInst_0_n31 ,
         SubCellInst2_LFInst_0_n30 , SubCellInst2_LFInst_0_n29 ,
         SubCellInst2_LFInst_0_n28 , SubCellInst2_LFInst_0_n27 ,
         SubCellInst2_LFInst_0_n26 , SubCellInst2_LFInst_0_n25 ,
         SubCellInst2_LFInst_0_n24 , SubCellInst2_LFInst_0_n23 ,
         SubCellInst2_LFInst_0_n22 , SubCellInst2_LFInst_1_n36 ,
         SubCellInst2_LFInst_1_n35 , SubCellInst2_LFInst_1_n34 ,
         SubCellInst2_LFInst_1_n33 , SubCellInst2_LFInst_1_n32 ,
         SubCellInst2_LFInst_1_n31 , SubCellInst2_LFInst_1_n30 ,
         SubCellInst2_LFInst_1_n29 , SubCellInst2_LFInst_1_n28 ,
         SubCellInst2_LFInst_1_n27 , SubCellInst2_LFInst_1_n26 ,
         SubCellInst2_LFInst_1_n25 , SubCellInst2_LFInst_1_n24 ,
         SubCellInst2_LFInst_1_n23 , SubCellInst2_LFInst_1_n22 ,
         SubCellInst2_LFInst_2_n36 , SubCellInst2_LFInst_2_n35 ,
         SubCellInst2_LFInst_2_n34 , SubCellInst2_LFInst_2_n33 ,
         SubCellInst2_LFInst_2_n32 , SubCellInst2_LFInst_2_n31 ,
         SubCellInst2_LFInst_2_n30 , SubCellInst2_LFInst_2_n29 ,
         SubCellInst2_LFInst_2_n28 , SubCellInst2_LFInst_2_n27 ,
         SubCellInst2_LFInst_2_n26 , SubCellInst2_LFInst_2_n25 ,
         SubCellInst2_LFInst_2_n24 , SubCellInst2_LFInst_2_n23 ,
         SubCellInst2_LFInst_2_n22 , SubCellInst2_LFInst_3_n36 ,
         SubCellInst2_LFInst_3_n35 , SubCellInst2_LFInst_3_n34 ,
         SubCellInst2_LFInst_3_n33 , SubCellInst2_LFInst_3_n32 ,
         SubCellInst2_LFInst_3_n31 , SubCellInst2_LFInst_3_n30 ,
         SubCellInst2_LFInst_3_n29 , SubCellInst2_LFInst_3_n28 ,
         SubCellInst2_LFInst_3_n27 , SubCellInst2_LFInst_3_n26 ,
         SubCellInst2_LFInst_3_n25 , SubCellInst2_LFInst_3_n24 ,
         SubCellInst2_LFInst_3_n23 , SubCellInst2_LFInst_3_n22 ,
         SubCellInst2_LFInst_4_n36 , SubCellInst2_LFInst_4_n35 ,
         SubCellInst2_LFInst_4_n34 , SubCellInst2_LFInst_4_n33 ,
         SubCellInst2_LFInst_4_n32 , SubCellInst2_LFInst_4_n31 ,
         SubCellInst2_LFInst_4_n30 , SubCellInst2_LFInst_4_n29 ,
         SubCellInst2_LFInst_4_n28 , SubCellInst2_LFInst_4_n27 ,
         SubCellInst2_LFInst_4_n26 , SubCellInst2_LFInst_4_n25 ,
         SubCellInst2_LFInst_4_n24 , SubCellInst2_LFInst_4_n23 ,
         SubCellInst2_LFInst_4_n22 , SubCellInst2_LFInst_5_n36 ,
         SubCellInst2_LFInst_5_n35 , SubCellInst2_LFInst_5_n34 ,
         SubCellInst2_LFInst_5_n33 , SubCellInst2_LFInst_5_n32 ,
         SubCellInst2_LFInst_5_n31 , SubCellInst2_LFInst_5_n30 ,
         SubCellInst2_LFInst_5_n29 , SubCellInst2_LFInst_5_n28 ,
         SubCellInst2_LFInst_5_n27 , SubCellInst2_LFInst_5_n26 ,
         SubCellInst2_LFInst_5_n25 , SubCellInst2_LFInst_5_n24 ,
         SubCellInst2_LFInst_5_n23 , SubCellInst2_LFInst_5_n22 ,
         SubCellInst2_LFInst_6_n36 , SubCellInst2_LFInst_6_n35 ,
         SubCellInst2_LFInst_6_n34 , SubCellInst2_LFInst_6_n33 ,
         SubCellInst2_LFInst_6_n32 , SubCellInst2_LFInst_6_n31 ,
         SubCellInst2_LFInst_6_n30 , SubCellInst2_LFInst_6_n29 ,
         SubCellInst2_LFInst_6_n28 , SubCellInst2_LFInst_6_n27 ,
         SubCellInst2_LFInst_6_n26 , SubCellInst2_LFInst_6_n25 ,
         SubCellInst2_LFInst_6_n24 , SubCellInst2_LFInst_6_n23 ,
         SubCellInst2_LFInst_6_n22 , SubCellInst2_LFInst_7_n36 ,
         SubCellInst2_LFInst_7_n35 , SubCellInst2_LFInst_7_n34 ,
         SubCellInst2_LFInst_7_n33 , SubCellInst2_LFInst_7_n32 ,
         SubCellInst2_LFInst_7_n31 , SubCellInst2_LFInst_7_n30 ,
         SubCellInst2_LFInst_7_n29 , SubCellInst2_LFInst_7_n28 ,
         SubCellInst2_LFInst_7_n27 , SubCellInst2_LFInst_7_n26 ,
         SubCellInst2_LFInst_7_n25 , SubCellInst2_LFInst_7_n24 ,
         SubCellInst2_LFInst_7_n23 , SubCellInst2_LFInst_7_n22 ,
         SubCellInst2_LFInst_8_n36 , SubCellInst2_LFInst_8_n35 ,
         SubCellInst2_LFInst_8_n34 , SubCellInst2_LFInst_8_n33 ,
         SubCellInst2_LFInst_8_n32 , SubCellInst2_LFInst_8_n31 ,
         SubCellInst2_LFInst_8_n30 , SubCellInst2_LFInst_8_n29 ,
         SubCellInst2_LFInst_8_n28 , SubCellInst2_LFInst_8_n27 ,
         SubCellInst2_LFInst_8_n26 , SubCellInst2_LFInst_8_n25 ,
         SubCellInst2_LFInst_8_n24 , SubCellInst2_LFInst_8_n23 ,
         SubCellInst2_LFInst_8_n22 , SubCellInst2_LFInst_9_n36 ,
         SubCellInst2_LFInst_9_n35 , SubCellInst2_LFInst_9_n34 ,
         SubCellInst2_LFInst_9_n33 , SubCellInst2_LFInst_9_n32 ,
         SubCellInst2_LFInst_9_n31 , SubCellInst2_LFInst_9_n30 ,
         SubCellInst2_LFInst_9_n29 , SubCellInst2_LFInst_9_n28 ,
         SubCellInst2_LFInst_9_n27 , SubCellInst2_LFInst_9_n26 ,
         SubCellInst2_LFInst_9_n25 , SubCellInst2_LFInst_9_n24 ,
         SubCellInst2_LFInst_9_n23 , SubCellInst2_LFInst_9_n22 ,
         SubCellInst2_LFInst_10_n36 , SubCellInst2_LFInst_10_n35 ,
         SubCellInst2_LFInst_10_n34 , SubCellInst2_LFInst_10_n33 ,
         SubCellInst2_LFInst_10_n32 , SubCellInst2_LFInst_10_n31 ,
         SubCellInst2_LFInst_10_n30 , SubCellInst2_LFInst_10_n29 ,
         SubCellInst2_LFInst_10_n28 , SubCellInst2_LFInst_10_n27 ,
         SubCellInst2_LFInst_10_n26 , SubCellInst2_LFInst_10_n25 ,
         SubCellInst2_LFInst_10_n24 , SubCellInst2_LFInst_10_n23 ,
         SubCellInst2_LFInst_10_n22 , SubCellInst2_LFInst_11_n36 ,
         SubCellInst2_LFInst_11_n35 , SubCellInst2_LFInst_11_n34 ,
         SubCellInst2_LFInst_11_n33 , SubCellInst2_LFInst_11_n32 ,
         SubCellInst2_LFInst_11_n31 , SubCellInst2_LFInst_11_n30 ,
         SubCellInst2_LFInst_11_n29 , SubCellInst2_LFInst_11_n28 ,
         SubCellInst2_LFInst_11_n27 , SubCellInst2_LFInst_11_n26 ,
         SubCellInst2_LFInst_11_n25 , SubCellInst2_LFInst_11_n24 ,
         SubCellInst2_LFInst_11_n23 , SubCellInst2_LFInst_11_n22 ,
         SubCellInst2_LFInst_12_n36 , SubCellInst2_LFInst_12_n35 ,
         SubCellInst2_LFInst_12_n34 , SubCellInst2_LFInst_12_n33 ,
         SubCellInst2_LFInst_12_n32 , SubCellInst2_LFInst_12_n31 ,
         SubCellInst2_LFInst_12_n30 , SubCellInst2_LFInst_12_n29 ,
         SubCellInst2_LFInst_12_n28 , SubCellInst2_LFInst_12_n27 ,
         SubCellInst2_LFInst_12_n26 , SubCellInst2_LFInst_12_n25 ,
         SubCellInst2_LFInst_12_n24 , SubCellInst2_LFInst_12_n23 ,
         SubCellInst2_LFInst_12_n22 , SubCellInst2_LFInst_13_n36 ,
         SubCellInst2_LFInst_13_n35 , SubCellInst2_LFInst_13_n34 ,
         SubCellInst2_LFInst_13_n33 , SubCellInst2_LFInst_13_n32 ,
         SubCellInst2_LFInst_13_n31 , SubCellInst2_LFInst_13_n30 ,
         SubCellInst2_LFInst_13_n29 , SubCellInst2_LFInst_13_n28 ,
         SubCellInst2_LFInst_13_n27 , SubCellInst2_LFInst_13_n26 ,
         SubCellInst2_LFInst_13_n25 , SubCellInst2_LFInst_13_n24 ,
         SubCellInst2_LFInst_13_n23 , SubCellInst2_LFInst_13_n22 ,
         SubCellInst2_LFInst_14_n36 , SubCellInst2_LFInst_14_n35 ,
         SubCellInst2_LFInst_14_n34 , SubCellInst2_LFInst_14_n33 ,
         SubCellInst2_LFInst_14_n32 , SubCellInst2_LFInst_14_n31 ,
         SubCellInst2_LFInst_14_n30 , SubCellInst2_LFInst_14_n29 ,
         SubCellInst2_LFInst_14_n28 , SubCellInst2_LFInst_14_n27 ,
         SubCellInst2_LFInst_14_n26 , SubCellInst2_LFInst_14_n25 ,
         SubCellInst2_LFInst_14_n24 , SubCellInst2_LFInst_14_n23 ,
         SubCellInst2_LFInst_14_n22 , SubCellInst2_LFInst_15_n36 ,
         SubCellInst2_LFInst_15_n35 , SubCellInst2_LFInst_15_n34 ,
         SubCellInst2_LFInst_15_n33 , SubCellInst2_LFInst_15_n32 ,
         SubCellInst2_LFInst_15_n31 , SubCellInst2_LFInst_15_n30 ,
         SubCellInst2_LFInst_15_n29 , SubCellInst2_LFInst_15_n28 ,
         SubCellInst2_LFInst_15_n27 , SubCellInst2_LFInst_15_n26 ,
         SubCellInst2_LFInst_15_n25 , SubCellInst2_LFInst_15_n24 ,
         SubCellInst2_LFInst_15_n23 , SubCellInst2_LFInst_15_n22 ;
  wire   [63:0] MCOutput;
  wire   [63:0] AddRoundKeyOutput;
  wire   [63:0] PermutationOutput;
  wire   [63:0] Feedback;
  wire   [63:0] MCOutput2;
  wire   [63:0] AddRoundKeyOutput2;
  wire   [63:0] PermutationOutput2;

  XNOR2_X1 MCInst_XOR_r0_Inst_0_U2  ( .A(MCInst_XOR_r0_Inst_0_n3 ), .B(
        Input[0]), .ZN(MCOutput[48]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_0_U1  ( .A(Input[48]), .B(Input[16]), .ZN(
        MCInst_XOR_r0_Inst_0_n3 ) );
  XOR2_X1 MCInst_XOR_r1_Inst_0_U1  ( .A(Input[32]), .B(Input[0]), .Z(
        MCOutput[32]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_1_U2  ( .A(MCInst_XOR_r0_Inst_1_n3 ), .B(
        Input[1]), .ZN(MCOutput[49]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_1_U1  ( .A(Input[49]), .B(Input[17]), .ZN(
        MCInst_XOR_r0_Inst_1_n3 ) );
  XOR2_X1 MCInst_XOR_r1_Inst_1_U1  ( .A(Input[33]), .B(Input[1]), .Z(
        MCOutput[33]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_2_U2  ( .A(MCInst_XOR_r0_Inst_2_n3 ), .B(
        Input[2]), .ZN(MCOutput[50]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_2_U1  ( .A(Input[50]), .B(Input[18]), .ZN(
        MCInst_XOR_r0_Inst_2_n3 ) );
  XOR2_X1 MCInst_XOR_r1_Inst_2_U1  ( .A(Input[34]), .B(Input[2]), .Z(
        MCOutput[34]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_3_U2  ( .A(MCInst_XOR_r0_Inst_3_n3 ), .B(
        Input[3]), .ZN(MCOutput[51]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_3_U1  ( .A(Input[51]), .B(Input[19]), .ZN(
        MCInst_XOR_r0_Inst_3_n3 ) );
  XOR2_X1 MCInst_XOR_r1_Inst_3_U1  ( .A(Input[35]), .B(Input[3]), .Z(
        MCOutput[35]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_4_U2  ( .A(MCInst_XOR_r0_Inst_4_n3 ), .B(
        Input[4]), .ZN(MCOutput[52]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_4_U1  ( .A(Input[52]), .B(Input[20]), .ZN(
        MCInst_XOR_r0_Inst_4_n3 ) );
  XOR2_X1 MCInst_XOR_r1_Inst_4_U1  ( .A(Input[36]), .B(Input[4]), .Z(
        MCOutput[36]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_5_U2  ( .A(MCInst_XOR_r0_Inst_5_n3 ), .B(
        Input[5]), .ZN(MCOutput[53]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_5_U1  ( .A(Input[53]), .B(Input[21]), .ZN(
        MCInst_XOR_r0_Inst_5_n3 ) );
  XOR2_X1 MCInst_XOR_r1_Inst_5_U1  ( .A(Input[37]), .B(Input[5]), .Z(
        MCOutput[37]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_6_U2  ( .A(MCInst_XOR_r0_Inst_6_n3 ), .B(
        Input[6]), .ZN(MCOutput[54]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_6_U1  ( .A(Input[54]), .B(Input[22]), .ZN(
        MCInst_XOR_r0_Inst_6_n3 ) );
  XOR2_X1 MCInst_XOR_r1_Inst_6_U1  ( .A(Input[38]), .B(Input[6]), .Z(
        MCOutput[38]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_7_U2  ( .A(MCInst_XOR_r0_Inst_7_n3 ), .B(
        Input[7]), .ZN(MCOutput[55]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_7_U1  ( .A(Input[55]), .B(Input[23]), .ZN(
        MCInst_XOR_r0_Inst_7_n3 ) );
  XOR2_X1 MCInst_XOR_r1_Inst_7_U1  ( .A(Input[39]), .B(Input[7]), .Z(
        MCOutput[39]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_8_U2  ( .A(MCInst_XOR_r0_Inst_8_n3 ), .B(
        Input[8]), .ZN(MCOutput[56]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_8_U1  ( .A(Input[56]), .B(Input[24]), .ZN(
        MCInst_XOR_r0_Inst_8_n3 ) );
  XOR2_X1 MCInst_XOR_r1_Inst_8_U1  ( .A(Input[40]), .B(Input[8]), .Z(
        MCOutput[40]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_9_U2  ( .A(MCInst_XOR_r0_Inst_9_n3 ), .B(
        Input[9]), .ZN(MCOutput[57]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_9_U1  ( .A(Input[57]), .B(Input[25]), .ZN(
        MCInst_XOR_r0_Inst_9_n3 ) );
  XOR2_X1 MCInst_XOR_r1_Inst_9_U1  ( .A(Input[41]), .B(Input[9]), .Z(
        MCOutput[41]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_10_U2  ( .A(MCInst_XOR_r0_Inst_10_n3 ), .B(
        Input[10]), .ZN(MCOutput[58]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_10_U1  ( .A(Input[58]), .B(Input[26]), .ZN(
        MCInst_XOR_r0_Inst_10_n3 ) );
  XOR2_X1 MCInst_XOR_r1_Inst_10_U1  ( .A(Input[42]), .B(Input[10]), .Z(
        MCOutput[42]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_11_U2  ( .A(MCInst_XOR_r0_Inst_11_n3 ), .B(
        Input[11]), .ZN(MCOutput[59]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_11_U1  ( .A(Input[59]), .B(Input[27]), .ZN(
        MCInst_XOR_r0_Inst_11_n3 ) );
  XOR2_X1 MCInst_XOR_r1_Inst_11_U1  ( .A(Input[43]), .B(Input[11]), .Z(
        MCOutput[43]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_12_U2  ( .A(MCInst_XOR_r0_Inst_12_n3 ), .B(
        Input[12]), .ZN(MCOutput[60]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_12_U1  ( .A(Input[60]), .B(Input[28]), .ZN(
        MCInst_XOR_r0_Inst_12_n3 ) );
  XOR2_X1 MCInst_XOR_r1_Inst_12_U1  ( .A(Input[44]), .B(Input[12]), .Z(
        MCOutput[44]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_13_U2  ( .A(MCInst_XOR_r0_Inst_13_n3 ), .B(
        Input[13]), .ZN(MCOutput[61]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_13_U1  ( .A(Input[61]), .B(Input[29]), .ZN(
        MCInst_XOR_r0_Inst_13_n3 ) );
  XOR2_X1 MCInst_XOR_r1_Inst_13_U1  ( .A(Input[45]), .B(Input[13]), .Z(
        MCOutput[45]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_14_U2  ( .A(MCInst_XOR_r0_Inst_14_n3 ), .B(
        Input[14]), .ZN(MCOutput[62]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_14_U1  ( .A(Input[62]), .B(Input[30]), .ZN(
        MCInst_XOR_r0_Inst_14_n3 ) );
  XOR2_X1 MCInst_XOR_r1_Inst_14_U1  ( .A(Input[46]), .B(Input[14]), .Z(
        MCOutput[46]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_15_U2  ( .A(MCInst_XOR_r0_Inst_15_n3 ), .B(
        Input[15]), .ZN(MCOutput[63]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_15_U1  ( .A(Input[63]), .B(Input[31]), .ZN(
        MCInst_XOR_r0_Inst_15_n3 ) );
  XOR2_X1 MCInst_XOR_r1_Inst_15_U1  ( .A(Input[47]), .B(Input[15]), .Z(
        MCOutput[47]) );
  XOR2_X1 AddKeyXOR1_XORInst_0_0_U1  ( .A(MCOutput[48]), .B(Key[112]), .Z(
        AddRoundKeyOutput[48]) );
  XOR2_X1 AddKeyXOR1_XORInst_0_1_U1  ( .A(MCOutput[49]), .B(Key[113]), .Z(
        AddRoundKeyOutput[49]) );
  XOR2_X1 AddKeyXOR1_XORInst_0_2_U1  ( .A(MCOutput[50]), .B(Key[114]), .Z(
        AddRoundKeyOutput[50]) );
  XOR2_X1 AddKeyXOR1_XORInst_0_3_U1  ( .A(MCOutput[51]), .B(Key[115]), .Z(
        AddRoundKeyOutput[51]) );
  XOR2_X1 AddKeyXOR1_XORInst_1_0_U1  ( .A(MCOutput[52]), .B(Key[116]), .Z(
        AddRoundKeyOutput[52]) );
  XOR2_X1 AddKeyXOR1_XORInst_1_1_U1  ( .A(MCOutput[53]), .B(Key[117]), .Z(
        AddRoundKeyOutput[53]) );
  XOR2_X1 AddKeyXOR1_XORInst_1_2_U1  ( .A(MCOutput[54]), .B(Key[118]), .Z(
        AddRoundKeyOutput[54]) );
  XOR2_X1 AddKeyXOR1_XORInst_1_3_U1  ( .A(MCOutput[55]), .B(Key[119]), .Z(
        AddRoundKeyOutput[55]) );
  XOR2_X1 AddKeyXOR1_XORInst_2_0_U1  ( .A(MCOutput[56]), .B(Key[120]), .Z(
        AddRoundKeyOutput[56]) );
  XOR2_X1 AddKeyXOR1_XORInst_2_1_U1  ( .A(MCOutput[57]), .B(Key[121]), .Z(
        AddRoundKeyOutput[57]) );
  XOR2_X1 AddKeyXOR1_XORInst_2_2_U1  ( .A(MCOutput[58]), .B(Key[122]), .Z(
        AddRoundKeyOutput[58]) );
  XOR2_X1 AddKeyXOR1_XORInst_2_3_U1  ( .A(MCOutput[59]), .B(Key[123]), .Z(
        AddRoundKeyOutput[59]) );
  XOR2_X1 AddKeyXOR1_XORInst_3_0_U1  ( .A(MCOutput[60]), .B(Key[124]), .Z(
        AddRoundKeyOutput[60]) );
  XOR2_X1 AddKeyXOR1_XORInst_3_1_U1  ( .A(MCOutput[61]), .B(Key[125]), .Z(
        AddRoundKeyOutput[61]) );
  XOR2_X1 AddKeyXOR1_XORInst_3_2_U1  ( .A(MCOutput[62]), .B(Key[126]), .Z(
        AddRoundKeyOutput[62]) );
  XOR2_X1 AddKeyXOR1_XORInst_3_3_U1  ( .A(MCOutput[63]), .B(Key[127]), .Z(
        AddRoundKeyOutput[63]) );
  XOR2_X1 AddKeyConstXOR_XORInst_0_0_U1  ( .A(Key[104]), .B(MCOutput[40]), 
        .Z(AddRoundKeyOutput[40]) );
  XOR2_X1 AddKeyConstXOR_XORInst_0_1_U1  ( .A(Key[105]), .B(MCOutput[41]), 
        .Z(AddRoundKeyOutput[41]) );
  XOR2_X1 AddKeyConstXOR_XORInst_0_2_U1  ( .A(Key[106]), .B(MCOutput[42]), 
        .Z(AddRoundKeyOutput[42]) );
  XOR2_X1 AddKeyConstXOR_XORInst_0_3_U1  ( .A(Key[107]), .B(MCOutput[43]), 
        .Z(AddRoundKeyOutput[43]) );
  XOR2_X1 AddKeyConstXOR_XORInst_1_0_U1  ( .A(Key[108]), .B(MCOutput[44]), 
        .Z(AddRoundKeyOutput[44]) );
  XOR2_X1 AddKeyConstXOR_XORInst_1_1_U1  ( .A(Key[109]), .B(MCOutput[45]), 
        .Z(AddRoundKeyOutput[45]) );
  XOR2_X1 AddKeyConstXOR_XORInst_1_2_U1  ( .A(Key[110]), .B(MCOutput[46]), 
        .Z(AddRoundKeyOutput[46]) );
  XOR2_X1 AddKeyConstXOR_XORInst_1_3_U1  ( .A(Key[111]), .B(MCOutput[47]), 
        .Z(AddRoundKeyOutput[47]) );
  XOR2_X1 AddKeyXOR2_XORInst_0_0_U1  ( .A(Input[0]), .B(Key[64]), .Z(
        AddRoundKeyOutput[0]) );
  XOR2_X1 AddKeyXOR2_XORInst_0_1_U1  ( .A(Input[1]), .B(Key[65]), .Z(
        AddRoundKeyOutput[1]) );
  XOR2_X1 AddKeyXOR2_XORInst_0_2_U1  ( .A(Input[2]), .B(Key[66]), .Z(
        AddRoundKeyOutput[2]) );
  XOR2_X1 AddKeyXOR2_XORInst_0_3_U1  ( .A(Input[3]), .B(Key[67]), .Z(
        AddRoundKeyOutput[3]) );
  XOR2_X1 AddKeyXOR2_XORInst_1_0_U1  ( .A(Input[4]), .B(Key[68]), .Z(
        AddRoundKeyOutput[4]) );
  XOR2_X1 AddKeyXOR2_XORInst_1_1_U1  ( .A(Input[5]), .B(Key[69]), .Z(
        AddRoundKeyOutput[5]) );
  XOR2_X1 AddKeyXOR2_XORInst_1_2_U1  ( .A(Input[6]), .B(Key[70]), .Z(
        AddRoundKeyOutput[6]) );
  XOR2_X1 AddKeyXOR2_XORInst_1_3_U1  ( .A(Input[7]), .B(Key[71]), .Z(
        AddRoundKeyOutput[7]) );
  XOR2_X1 AddKeyXOR2_XORInst_2_0_U1  ( .A(Input[8]), .B(Key[72]), .Z(
        AddRoundKeyOutput[8]) );
  XOR2_X1 AddKeyXOR2_XORInst_2_1_U1  ( .A(Input[9]), .B(Key[73]), .Z(
        AddRoundKeyOutput[9]) );
  XOR2_X1 AddKeyXOR2_XORInst_2_2_U1  ( .A(Input[10]), .B(Key[74]), .Z(
        AddRoundKeyOutput[10]) );
  XOR2_X1 AddKeyXOR2_XORInst_2_3_U1  ( .A(Input[11]), .B(Key[75]), .Z(
        AddRoundKeyOutput[11]) );
  XOR2_X1 AddKeyXOR2_XORInst_3_0_U1  ( .A(Input[12]), .B(Key[76]), .Z(
        AddRoundKeyOutput[12]) );
  XOR2_X1 AddKeyXOR2_XORInst_3_1_U1  ( .A(Input[13]), .B(Key[77]), .Z(
        AddRoundKeyOutput[13]) );
  XOR2_X1 AddKeyXOR2_XORInst_3_2_U1  ( .A(Input[14]), .B(Key[78]), .Z(
        AddRoundKeyOutput[14]) );
  XOR2_X1 AddKeyXOR2_XORInst_3_3_U1  ( .A(Input[15]), .B(Key[79]), .Z(
        AddRoundKeyOutput[15]) );
  XOR2_X1 AddKeyXOR2_XORInst_4_0_U1  ( .A(Input[16]), .B(Key[80]), .Z(
        AddRoundKeyOutput[16]) );
  XOR2_X1 AddKeyXOR2_XORInst_4_1_U1  ( .A(Input[17]), .B(Key[81]), .Z(
        AddRoundKeyOutput[17]) );
  XOR2_X1 AddKeyXOR2_XORInst_4_2_U1  ( .A(Input[18]), .B(Key[82]), .Z(
        AddRoundKeyOutput[18]) );
  XOR2_X1 AddKeyXOR2_XORInst_4_3_U1  ( .A(Input[19]), .B(Key[83]), .Z(
        AddRoundKeyOutput[19]) );
  XOR2_X1 AddKeyXOR2_XORInst_5_0_U1  ( .A(Input[20]), .B(Key[84]), .Z(
        AddRoundKeyOutput[20]) );
  XOR2_X1 AddKeyXOR2_XORInst_5_1_U1  ( .A(Input[21]), .B(Key[85]), .Z(
        AddRoundKeyOutput[21]) );
  XOR2_X1 AddKeyXOR2_XORInst_5_2_U1  ( .A(Input[22]), .B(Key[86]), .Z(
        AddRoundKeyOutput[22]) );
  XOR2_X1 AddKeyXOR2_XORInst_5_3_U1  ( .A(Input[23]), .B(Key[87]), .Z(
        AddRoundKeyOutput[23]) );
  XOR2_X1 AddKeyXOR2_XORInst_6_0_U1  ( .A(Input[24]), .B(Key[88]), .Z(
        AddRoundKeyOutput[24]) );
  XOR2_X1 AddKeyXOR2_XORInst_6_1_U1  ( .A(Input[25]), .B(Key[89]), .Z(
        AddRoundKeyOutput[25]) );
  XOR2_X1 AddKeyXOR2_XORInst_6_2_U1  ( .A(Input[26]), .B(Key[90]), .Z(
        AddRoundKeyOutput[26]) );
  XOR2_X1 AddKeyXOR2_XORInst_6_3_U1  ( .A(Input[27]), .B(Key[91]), .Z(
        AddRoundKeyOutput[27]) );
  XOR2_X1 AddKeyXOR2_XORInst_7_0_U1  ( .A(Input[28]), .B(Key[92]), .Z(
        AddRoundKeyOutput[28]) );
  XOR2_X1 AddKeyXOR2_XORInst_7_1_U1  ( .A(Input[29]), .B(Key[93]), .Z(
        AddRoundKeyOutput[29]) );
  XOR2_X1 AddKeyXOR2_XORInst_7_2_U1  ( .A(Input[30]), .B(Key[94]), .Z(
        AddRoundKeyOutput[30]) );
  XOR2_X1 AddKeyXOR2_XORInst_7_3_U1  ( .A(Input[31]), .B(Key[95]), .Z(
        AddRoundKeyOutput[31]) );
  XOR2_X1 AddKeyXOR2_XORInst_8_0_U1  ( .A(MCOutput[32]), .B(Key[96]), .Z(
        AddRoundKeyOutput[32]) );
  XOR2_X1 AddKeyXOR2_XORInst_8_1_U1  ( .A(MCOutput[33]), .B(Key[97]), .Z(
        AddRoundKeyOutput[33]) );
  XOR2_X1 AddKeyXOR2_XORInst_8_2_U1  ( .A(MCOutput[34]), .B(Key[98]), .Z(
        AddRoundKeyOutput[34]) );
  XOR2_X1 AddKeyXOR2_XORInst_8_3_U1  ( .A(MCOutput[35]), .B(Key[99]), .Z(
        AddRoundKeyOutput[35]) );
  XOR2_X1 AddKeyXOR2_XORInst_9_0_U1  ( .A(MCOutput[36]), .B(Key[100]), .Z(
        AddRoundKeyOutput[36]) );
  XOR2_X1 AddKeyXOR2_XORInst_9_1_U1  ( .A(MCOutput[37]), .B(Key[101]), .Z(
        AddRoundKeyOutput[37]) );
  XOR2_X1 AddKeyXOR2_XORInst_9_2_U1  ( .A(MCOutput[38]), .B(Key[102]), .Z(
        AddRoundKeyOutput[38]) );
  XOR2_X1 AddKeyXOR2_XORInst_9_3_U1  ( .A(MCOutput[39]), .B(Key[103]), .Z(
        AddRoundKeyOutput[39]) );
  DFF_X1 StateReg_s_current_state_reg[0]  ( .D(AddRoundKeyOutput[0]), .CK(clk), .Q(PermutationOutput[60]) );
  DFF_X1 StateReg_s_current_state_reg[1]  ( .D(AddRoundKeyOutput[1]), .CK(clk), .Q(PermutationOutput[61]) );
  DFF_X1 StateReg_s_current_state_reg[2]  ( .D(AddRoundKeyOutput[2]), .CK(clk), .Q(PermutationOutput[62]) );
  DFF_X1 StateReg_s_current_state_reg[3]  ( .D(AddRoundKeyOutput[3]), .CK(clk), .Q(PermutationOutput[63]) );
  DFF_X1 StateReg_s_current_state_reg[4]  ( .D(AddRoundKeyOutput[4]), .CK(clk), .Q(PermutationOutput[48]) );
  DFF_X1 StateReg_s_current_state_reg[5]  ( .D(AddRoundKeyOutput[5]), .CK(clk), .Q(PermutationOutput[49]) );
  DFF_X1 StateReg_s_current_state_reg[6]  ( .D(AddRoundKeyOutput[6]), .CK(clk), .Q(PermutationOutput[50]) );
  DFF_X1 StateReg_s_current_state_reg[7]  ( .D(AddRoundKeyOutput[7]), .CK(clk), .Q(PermutationOutput[51]) );
  DFF_X1 StateReg_s_current_state_reg[8]  ( .D(AddRoundKeyOutput[8]), .CK(clk), .Q(PermutationOutput[52]) );
  DFF_X1 StateReg_s_current_state_reg[9]  ( .D(AddRoundKeyOutput[9]), .CK(clk), .Q(PermutationOutput[53]) );
  DFF_X1 StateReg_s_current_state_reg[10]  ( .D(AddRoundKeyOutput[10]), .CK(
        clk), .Q(PermutationOutput[54]) );
  DFF_X1 StateReg_s_current_state_reg[11]  ( .D(AddRoundKeyOutput[11]), .CK(
        clk), .Q(PermutationOutput[55]) );
  DFF_X1 StateReg_s_current_state_reg[12]  ( .D(AddRoundKeyOutput[12]), .CK(
        clk), .Q(PermutationOutput[56]) );
  DFF_X1 StateReg_s_current_state_reg[13]  ( .D(AddRoundKeyOutput[13]), .CK(
        clk), .Q(PermutationOutput[57]) );
  DFF_X1 StateReg_s_current_state_reg[14]  ( .D(AddRoundKeyOutput[14]), .CK(
        clk), .Q(PermutationOutput[58]) );
  DFF_X1 StateReg_s_current_state_reg[15]  ( .D(AddRoundKeyOutput[15]), .CK(
        clk), .Q(PermutationOutput[59]) );
  DFF_X1 StateReg_s_current_state_reg[16]  ( .D(AddRoundKeyOutput[16]), .CK(
        clk), .Q(PermutationOutput[32]) );
  DFF_X1 StateReg_s_current_state_reg[17]  ( .D(AddRoundKeyOutput[17]), .CK(
        clk), .Q(PermutationOutput[33]) );
  DFF_X1 StateReg_s_current_state_reg[18]  ( .D(AddRoundKeyOutput[18]), .CK(
        clk), .Q(PermutationOutput[34]) );
  DFF_X1 StateReg_s_current_state_reg[19]  ( .D(AddRoundKeyOutput[19]), .CK(
        clk), .Q(PermutationOutput[35]) );
  DFF_X1 StateReg_s_current_state_reg[20]  ( .D(AddRoundKeyOutput[20]), .CK(
        clk), .Q(PermutationOutput[44]) );
  DFF_X1 StateReg_s_current_state_reg[21]  ( .D(AddRoundKeyOutput[21]), .CK(
        clk), .Q(PermutationOutput[45]) );
  DFF_X1 StateReg_s_current_state_reg[22]  ( .D(AddRoundKeyOutput[22]), .CK(
        clk), .Q(PermutationOutput[46]) );
  DFF_X1 StateReg_s_current_state_reg[23]  ( .D(AddRoundKeyOutput[23]), .CK(
        clk), .Q(PermutationOutput[47]) );
  DFF_X1 StateReg_s_current_state_reg[24]  ( .D(AddRoundKeyOutput[24]), .CK(
        clk), .Q(PermutationOutput[40]) );
  DFF_X1 StateReg_s_current_state_reg[25]  ( .D(AddRoundKeyOutput[25]), .CK(
        clk), .Q(PermutationOutput[41]) );
  DFF_X1 StateReg_s_current_state_reg[26]  ( .D(AddRoundKeyOutput[26]), .CK(
        clk), .Q(PermutationOutput[42]) );
  DFF_X1 StateReg_s_current_state_reg[27]  ( .D(AddRoundKeyOutput[27]), .CK(
        clk), .Q(PermutationOutput[43]) );
  DFF_X1 StateReg_s_current_state_reg[28]  ( .D(AddRoundKeyOutput[28]), .CK(
        clk), .Q(PermutationOutput[36]) );
  DFF_X1 StateReg_s_current_state_reg[29]  ( .D(AddRoundKeyOutput[29]), .CK(
        clk), .Q(PermutationOutput[37]) );
  DFF_X1 StateReg_s_current_state_reg[30]  ( .D(AddRoundKeyOutput[30]), .CK(
        clk), .Q(PermutationOutput[38]) );
  DFF_X1 StateReg_s_current_state_reg[31]  ( .D(AddRoundKeyOutput[31]), .CK(
        clk), .Q(PermutationOutput[39]) );
  DFF_X1 StateReg_s_current_state_reg[32]  ( .D(AddRoundKeyOutput[32]), .CK(
        clk), .Q(PermutationOutput[16]) );
  DFF_X1 StateReg_s_current_state_reg[33]  ( .D(AddRoundKeyOutput[33]), .CK(
        clk), .Q(PermutationOutput[17]) );
  DFF_X1 StateReg_s_current_state_reg[34]  ( .D(AddRoundKeyOutput[34]), .CK(
        clk), .Q(PermutationOutput[18]) );
  DFF_X1 StateReg_s_current_state_reg[35]  ( .D(AddRoundKeyOutput[35]), .CK(
        clk), .Q(PermutationOutput[19]) );
  DFF_X1 StateReg_s_current_state_reg[36]  ( .D(AddRoundKeyOutput[36]), .CK(
        clk), .Q(PermutationOutput[28]) );
  DFF_X1 StateReg_s_current_state_reg[37]  ( .D(AddRoundKeyOutput[37]), .CK(
        clk), .Q(PermutationOutput[29]) );
  DFF_X1 StateReg_s_current_state_reg[38]  ( .D(AddRoundKeyOutput[38]), .CK(
        clk), .Q(PermutationOutput[30]) );
  DFF_X1 StateReg_s_current_state_reg[39]  ( .D(AddRoundKeyOutput[39]), .CK(
        clk), .Q(PermutationOutput[31]) );
  DFF_X1 StateReg_s_current_state_reg[40]  ( .D(AddRoundKeyOutput[40]), .CK(
        clk), .Q(PermutationOutput[24]) );
  DFF_X1 StateReg_s_current_state_reg[41]  ( .D(AddRoundKeyOutput[41]), .CK(
        clk), .Q(PermutationOutput[25]) );
  DFF_X1 StateReg_s_current_state_reg[42]  ( .D(AddRoundKeyOutput[42]), .CK(
        clk), .Q(PermutationOutput[26]) );
  DFF_X1 StateReg_s_current_state_reg[43]  ( .D(AddRoundKeyOutput[43]), .CK(
        clk), .Q(PermutationOutput[27]) );
  DFF_X1 StateReg_s_current_state_reg[44]  ( .D(AddRoundKeyOutput[44]), .CK(
        clk), .Q(PermutationOutput[20]) );
  DFF_X1 StateReg_s_current_state_reg[45]  ( .D(AddRoundKeyOutput[45]), .CK(
        clk), .Q(PermutationOutput[21]) );
  DFF_X1 StateReg_s_current_state_reg[46]  ( .D(AddRoundKeyOutput[46]), .CK(
        clk), .Q(PermutationOutput[22]) );
  DFF_X1 StateReg_s_current_state_reg[47]  ( .D(AddRoundKeyOutput[47]), .CK(
        clk), .Q(PermutationOutput[23]) );
  DFF_X1 StateReg_s_current_state_reg[48]  ( .D(AddRoundKeyOutput[48]), .CK(
        clk), .Q(PermutationOutput[4]) );
  DFF_X1 StateReg_s_current_state_reg[49]  ( .D(AddRoundKeyOutput[49]), .CK(
        clk), .Q(PermutationOutput[5]) );
  DFF_X1 StateReg_s_current_state_reg[50]  ( .D(AddRoundKeyOutput[50]), .CK(
        clk), .Q(PermutationOutput[6]) );
  DFF_X1 StateReg_s_current_state_reg[51]  ( .D(AddRoundKeyOutput[51]), .CK(
        clk), .Q(PermutationOutput[7]) );
  DFF_X1 StateReg_s_current_state_reg[52]  ( .D(AddRoundKeyOutput[52]), .CK(
        clk), .Q(PermutationOutput[8]) );
  DFF_X1 StateReg_s_current_state_reg[53]  ( .D(AddRoundKeyOutput[53]), .CK(
        clk), .Q(PermutationOutput[9]) );
  DFF_X1 StateReg_s_current_state_reg[54]  ( .D(AddRoundKeyOutput[54]), .CK(
        clk), .Q(PermutationOutput[10]) );
  DFF_X1 StateReg_s_current_state_reg[55]  ( .D(AddRoundKeyOutput[55]), .CK(
        clk), .Q(PermutationOutput[11]) );
  DFF_X1 StateReg_s_current_state_reg[56]  ( .D(AddRoundKeyOutput[56]), .CK(
        clk), .Q(PermutationOutput[12]) );
  DFF_X1 StateReg_s_current_state_reg[57]  ( .D(AddRoundKeyOutput[57]), .CK(
        clk), .Q(PermutationOutput[13]) );
  DFF_X1 StateReg_s_current_state_reg[58]  ( .D(AddRoundKeyOutput[58]), .CK(
        clk), .Q(PermutationOutput[14]) );
  DFF_X1 StateReg_s_current_state_reg[59]  ( .D(AddRoundKeyOutput[59]), .CK(
        clk), .Q(PermutationOutput[15]) );
  DFF_X1 StateReg_s_current_state_reg[60]  ( .D(AddRoundKeyOutput[60]), .CK(
        clk), .Q(PermutationOutput[0]) );
  DFF_X1 StateReg_s_current_state_reg[61]  ( .D(AddRoundKeyOutput[61]), .CK(
        clk), .Q(PermutationOutput[1]) );
  DFF_X1 StateReg_s_current_state_reg[62]  ( .D(AddRoundKeyOutput[62]), .CK(
        clk), .Q(PermutationOutput[2]) );
  DFF_X1 StateReg_s_current_state_reg[63]  ( .D(AddRoundKeyOutput[63]), .CK(
        clk), .Q(PermutationOutput[3]) );
  NOR2_X1 SubCellInst_LFInst_0_U21  ( .A1(SubCellInst_LFInst_0_n36 ), .A2(
        SubCellInst_LFInst_0_n35 ), .ZN(MCOutput2[0]) );
  NOR2_X1 SubCellInst_LFInst_0_U20  ( .A1(PermutationOutput[1]), .A2(
        SubCellInst_LFInst_0_n34 ), .ZN(SubCellInst_LFInst_0_n36 ) );
  NOR2_X1 SubCellInst_LFInst_0_U19  ( .A1(SubCellInst_LFInst_0_n33 ), .A2(
        SubCellInst_LFInst_0_n32 ), .ZN(SubCellInst_LFInst_0_n34 ) );
  NOR2_X1 SubCellInst_LFInst_0_U18  ( .A1(PermutationOutput[2]), .A2(
        PermutationOutput[3]), .ZN(SubCellInst_LFInst_0_n32 ) );
  NAND2_X1 SubCellInst_LFInst_0_U17  ( .A1(SubCellInst_LFInst_0_n31 ), .A2(
        SubCellInst_LFInst_0_n30 ), .ZN(MCOutput2[1]) );
  NAND2_X1 SubCellInst_LFInst_0_U16  ( .A1(PermutationOutput[0]), .A2(
        SubCellInst_LFInst_0_n29 ), .ZN(SubCellInst_LFInst_0_n30 ) );
  NAND2_X1 SubCellInst_LFInst_0_U15  ( .A1(PermutationOutput[2]), .A2(
        SubCellInst_LFInst_0_n28 ), .ZN(SubCellInst_LFInst_0_n31 ) );
  NAND2_X1 SubCellInst_LFInst_0_U14  ( .A1(PermutationOutput[3]), .A2(
        SubCellInst_LFInst_0_n33 ), .ZN(SubCellInst_LFInst_0_n28 ) );
  NAND2_X1 SubCellInst_LFInst_0_U13  ( .A1(SubCellInst_LFInst_0_n27 ), .A2(
        SubCellInst_LFInst_0_n26 ), .ZN(MCOutput2[2]) );
  NAND2_X1 SubCellInst_LFInst_0_U12  ( .A1(SubCellInst_LFInst_0_n25 ), .A2(
        PermutationOutput[1]), .ZN(SubCellInst_LFInst_0_n27 ) );
  NAND2_X1 SubCellInst_LFInst_0_U11  ( .A1(SubCellInst_LFInst_0_n24 ), .A2(
        SubCellInst_LFInst_0_n23 ), .ZN(SubCellInst_LFInst_0_n25 ) );
  NAND2_X1 SubCellInst_LFInst_0_U10  ( .A1(PermutationOutput[0]), .A2(
        PermutationOutput[3]), .ZN(SubCellInst_LFInst_0_n24 ) );
  NAND2_X1 SubCellInst_LFInst_0_U9  ( .A1(SubCellInst_LFInst_0_n26 ), .A2(
        SubCellInst_LFInst_0_n22 ), .ZN(MCOutput2[3]) );
  OR2_X1 SubCellInst_LFInst_0_U8  ( .A1(PermutationOutput[1]), .A2(
        SubCellInst_LFInst_0_n35 ), .ZN(SubCellInst_LFInst_0_n22 ) );
  NOR2_X1 SubCellInst_LFInst_0_U7  ( .A1(SubCellInst_LFInst_0_n23 ), .A2(
        SubCellInst_LFInst_0_n29 ), .ZN(SubCellInst_LFInst_0_n35 ) );
  INV_X1 SubCellInst_LFInst_0_U6  ( .A(PermutationOutput[2]), .ZN(
        SubCellInst_LFInst_0_n23 ) );
  NAND2_X1 SubCellInst_LFInst_0_U5  ( .A1(SubCellInst_LFInst_0_n29 ), .A2(
        SubCellInst_LFInst_0_n33 ), .ZN(SubCellInst_LFInst_0_n26 ) );
  INV_X1 SubCellInst_LFInst_0_U4  ( .A(PermutationOutput[0]), .ZN(
        SubCellInst_LFInst_0_n33 ) );
  INV_X1 SubCellInst_LFInst_0_U3  ( .A(PermutationOutput[3]), .ZN(
        SubCellInst_LFInst_0_n29 ) );
  NOR2_X1 SubCellInst_LFInst_1_U21  ( .A1(SubCellInst_LFInst_1_n36 ), .A2(
        SubCellInst_LFInst_1_n35 ), .ZN(MCOutput2[4]) );
  NOR2_X1 SubCellInst_LFInst_1_U20  ( .A1(PermutationOutput[5]), .A2(
        SubCellInst_LFInst_1_n34 ), .ZN(SubCellInst_LFInst_1_n36 ) );
  NOR2_X1 SubCellInst_LFInst_1_U19  ( .A1(SubCellInst_LFInst_1_n33 ), .A2(
        SubCellInst_LFInst_1_n32 ), .ZN(SubCellInst_LFInst_1_n34 ) );
  NOR2_X1 SubCellInst_LFInst_1_U18  ( .A1(PermutationOutput[6]), .A2(
        PermutationOutput[7]), .ZN(SubCellInst_LFInst_1_n32 ) );
  NAND2_X1 SubCellInst_LFInst_1_U17  ( .A1(SubCellInst_LFInst_1_n31 ), .A2(
        SubCellInst_LFInst_1_n30 ), .ZN(MCOutput2[5]) );
  NAND2_X1 SubCellInst_LFInst_1_U16  ( .A1(PermutationOutput[4]), .A2(
        SubCellInst_LFInst_1_n29 ), .ZN(SubCellInst_LFInst_1_n30 ) );
  NAND2_X1 SubCellInst_LFInst_1_U15  ( .A1(PermutationOutput[6]), .A2(
        SubCellInst_LFInst_1_n28 ), .ZN(SubCellInst_LFInst_1_n31 ) );
  NAND2_X1 SubCellInst_LFInst_1_U14  ( .A1(PermutationOutput[7]), .A2(
        SubCellInst_LFInst_1_n33 ), .ZN(SubCellInst_LFInst_1_n28 ) );
  NAND2_X1 SubCellInst_LFInst_1_U13  ( .A1(SubCellInst_LFInst_1_n27 ), .A2(
        SubCellInst_LFInst_1_n26 ), .ZN(MCOutput2[6]) );
  NAND2_X1 SubCellInst_LFInst_1_U12  ( .A1(SubCellInst_LFInst_1_n25 ), .A2(
        PermutationOutput[5]), .ZN(SubCellInst_LFInst_1_n27 ) );
  NAND2_X1 SubCellInst_LFInst_1_U11  ( .A1(SubCellInst_LFInst_1_n24 ), .A2(
        SubCellInst_LFInst_1_n23 ), .ZN(SubCellInst_LFInst_1_n25 ) );
  NAND2_X1 SubCellInst_LFInst_1_U10  ( .A1(PermutationOutput[4]), .A2(
        PermutationOutput[7]), .ZN(SubCellInst_LFInst_1_n24 ) );
  NAND2_X1 SubCellInst_LFInst_1_U9  ( .A1(SubCellInst_LFInst_1_n26 ), .A2(
        SubCellInst_LFInst_1_n22 ), .ZN(MCOutput2[7]) );
  OR2_X1 SubCellInst_LFInst_1_U8  ( .A1(PermutationOutput[5]), .A2(
        SubCellInst_LFInst_1_n35 ), .ZN(SubCellInst_LFInst_1_n22 ) );
  NOR2_X1 SubCellInst_LFInst_1_U7  ( .A1(SubCellInst_LFInst_1_n23 ), .A2(
        SubCellInst_LFInst_1_n29 ), .ZN(SubCellInst_LFInst_1_n35 ) );
  INV_X1 SubCellInst_LFInst_1_U6  ( .A(PermutationOutput[6]), .ZN(
        SubCellInst_LFInst_1_n23 ) );
  NAND2_X1 SubCellInst_LFInst_1_U5  ( .A1(SubCellInst_LFInst_1_n29 ), .A2(
        SubCellInst_LFInst_1_n33 ), .ZN(SubCellInst_LFInst_1_n26 ) );
  INV_X1 SubCellInst_LFInst_1_U4  ( .A(PermutationOutput[4]), .ZN(
        SubCellInst_LFInst_1_n33 ) );
  INV_X1 SubCellInst_LFInst_1_U3  ( .A(PermutationOutput[7]), .ZN(
        SubCellInst_LFInst_1_n29 ) );
  NOR2_X1 SubCellInst_LFInst_2_U21  ( .A1(SubCellInst_LFInst_2_n36 ), .A2(
        SubCellInst_LFInst_2_n35 ), .ZN(MCOutput2[8]) );
  NOR2_X1 SubCellInst_LFInst_2_U20  ( .A1(PermutationOutput[9]), .A2(
        SubCellInst_LFInst_2_n34 ), .ZN(SubCellInst_LFInst_2_n36 ) );
  NOR2_X1 SubCellInst_LFInst_2_U19  ( .A1(SubCellInst_LFInst_2_n33 ), .A2(
        SubCellInst_LFInst_2_n32 ), .ZN(SubCellInst_LFInst_2_n34 ) );
  NOR2_X1 SubCellInst_LFInst_2_U18  ( .A1(PermutationOutput[10]), .A2(
        PermutationOutput[11]), .ZN(SubCellInst_LFInst_2_n32 ) );
  NAND2_X1 SubCellInst_LFInst_2_U17  ( .A1(SubCellInst_LFInst_2_n31 ), .A2(
        SubCellInst_LFInst_2_n30 ), .ZN(MCOutput2[9]) );
  NAND2_X1 SubCellInst_LFInst_2_U16  ( .A1(PermutationOutput[8]), .A2(
        SubCellInst_LFInst_2_n29 ), .ZN(SubCellInst_LFInst_2_n30 ) );
  NAND2_X1 SubCellInst_LFInst_2_U15  ( .A1(PermutationOutput[10]), .A2(
        SubCellInst_LFInst_2_n28 ), .ZN(SubCellInst_LFInst_2_n31 ) );
  NAND2_X1 SubCellInst_LFInst_2_U14  ( .A1(PermutationOutput[11]), .A2(
        SubCellInst_LFInst_2_n33 ), .ZN(SubCellInst_LFInst_2_n28 ) );
  NAND2_X1 SubCellInst_LFInst_2_U13  ( .A1(SubCellInst_LFInst_2_n27 ), .A2(
        SubCellInst_LFInst_2_n26 ), .ZN(MCOutput2[10]) );
  NAND2_X1 SubCellInst_LFInst_2_U12  ( .A1(SubCellInst_LFInst_2_n25 ), .A2(
        PermutationOutput[9]), .ZN(SubCellInst_LFInst_2_n27 ) );
  NAND2_X1 SubCellInst_LFInst_2_U11  ( .A1(SubCellInst_LFInst_2_n24 ), .A2(
        SubCellInst_LFInst_2_n23 ), .ZN(SubCellInst_LFInst_2_n25 ) );
  NAND2_X1 SubCellInst_LFInst_2_U10  ( .A1(PermutationOutput[8]), .A2(
        PermutationOutput[11]), .ZN(SubCellInst_LFInst_2_n24 ) );
  NAND2_X1 SubCellInst_LFInst_2_U9  ( .A1(SubCellInst_LFInst_2_n26 ), .A2(
        SubCellInst_LFInst_2_n22 ), .ZN(MCOutput2[11]) );
  OR2_X1 SubCellInst_LFInst_2_U8  ( .A1(PermutationOutput[9]), .A2(
        SubCellInst_LFInst_2_n35 ), .ZN(SubCellInst_LFInst_2_n22 ) );
  NOR2_X1 SubCellInst_LFInst_2_U7  ( .A1(SubCellInst_LFInst_2_n23 ), .A2(
        SubCellInst_LFInst_2_n29 ), .ZN(SubCellInst_LFInst_2_n35 ) );
  INV_X1 SubCellInst_LFInst_2_U6  ( .A(PermutationOutput[10]), .ZN(
        SubCellInst_LFInst_2_n23 ) );
  NAND2_X1 SubCellInst_LFInst_2_U5  ( .A1(SubCellInst_LFInst_2_n29 ), .A2(
        SubCellInst_LFInst_2_n33 ), .ZN(SubCellInst_LFInst_2_n26 ) );
  INV_X1 SubCellInst_LFInst_2_U4  ( .A(PermutationOutput[8]), .ZN(
        SubCellInst_LFInst_2_n33 ) );
  INV_X1 SubCellInst_LFInst_2_U3  ( .A(PermutationOutput[11]), .ZN(
        SubCellInst_LFInst_2_n29 ) );
  NOR2_X1 SubCellInst_LFInst_3_U21  ( .A1(SubCellInst_LFInst_3_n36 ), .A2(
        SubCellInst_LFInst_3_n35 ), .ZN(MCOutput2[12]) );
  NOR2_X1 SubCellInst_LFInst_3_U20  ( .A1(PermutationOutput[13]), .A2(
        SubCellInst_LFInst_3_n34 ), .ZN(SubCellInst_LFInst_3_n36 ) );
  NOR2_X1 SubCellInst_LFInst_3_U19  ( .A1(SubCellInst_LFInst_3_n33 ), .A2(
        SubCellInst_LFInst_3_n32 ), .ZN(SubCellInst_LFInst_3_n34 ) );
  NOR2_X1 SubCellInst_LFInst_3_U18  ( .A1(PermutationOutput[14]), .A2(
        PermutationOutput[15]), .ZN(SubCellInst_LFInst_3_n32 ) );
  NAND2_X1 SubCellInst_LFInst_3_U17  ( .A1(SubCellInst_LFInst_3_n31 ), .A2(
        SubCellInst_LFInst_3_n30 ), .ZN(MCOutput2[13]) );
  NAND2_X1 SubCellInst_LFInst_3_U16  ( .A1(PermutationOutput[12]), .A2(
        SubCellInst_LFInst_3_n29 ), .ZN(SubCellInst_LFInst_3_n30 ) );
  NAND2_X1 SubCellInst_LFInst_3_U15  ( .A1(PermutationOutput[14]), .A2(
        SubCellInst_LFInst_3_n28 ), .ZN(SubCellInst_LFInst_3_n31 ) );
  NAND2_X1 SubCellInst_LFInst_3_U14  ( .A1(PermutationOutput[15]), .A2(
        SubCellInst_LFInst_3_n33 ), .ZN(SubCellInst_LFInst_3_n28 ) );
  NAND2_X1 SubCellInst_LFInst_3_U13  ( .A1(SubCellInst_LFInst_3_n27 ), .A2(
        SubCellInst_LFInst_3_n26 ), .ZN(MCOutput2[14]) );
  NAND2_X1 SubCellInst_LFInst_3_U12  ( .A1(SubCellInst_LFInst_3_n25 ), .A2(
        PermutationOutput[13]), .ZN(SubCellInst_LFInst_3_n27 ) );
  NAND2_X1 SubCellInst_LFInst_3_U11  ( .A1(SubCellInst_LFInst_3_n24 ), .A2(
        SubCellInst_LFInst_3_n23 ), .ZN(SubCellInst_LFInst_3_n25 ) );
  NAND2_X1 SubCellInst_LFInst_3_U10  ( .A1(PermutationOutput[12]), .A2(
        PermutationOutput[15]), .ZN(SubCellInst_LFInst_3_n24 ) );
  NAND2_X1 SubCellInst_LFInst_3_U9  ( .A1(SubCellInst_LFInst_3_n26 ), .A2(
        SubCellInst_LFInst_3_n22 ), .ZN(MCOutput2[15]) );
  OR2_X1 SubCellInst_LFInst_3_U8  ( .A1(PermutationOutput[13]), .A2(
        SubCellInst_LFInst_3_n35 ), .ZN(SubCellInst_LFInst_3_n22 ) );
  NOR2_X1 SubCellInst_LFInst_3_U7  ( .A1(SubCellInst_LFInst_3_n23 ), .A2(
        SubCellInst_LFInst_3_n29 ), .ZN(SubCellInst_LFInst_3_n35 ) );
  INV_X1 SubCellInst_LFInst_3_U6  ( .A(PermutationOutput[14]), .ZN(
        SubCellInst_LFInst_3_n23 ) );
  NAND2_X1 SubCellInst_LFInst_3_U5  ( .A1(SubCellInst_LFInst_3_n29 ), .A2(
        SubCellInst_LFInst_3_n33 ), .ZN(SubCellInst_LFInst_3_n26 ) );
  INV_X1 SubCellInst_LFInst_3_U4  ( .A(PermutationOutput[12]), .ZN(
        SubCellInst_LFInst_3_n33 ) );
  INV_X1 SubCellInst_LFInst_3_U3  ( .A(PermutationOutput[15]), .ZN(
        SubCellInst_LFInst_3_n29 ) );
  NOR2_X1 SubCellInst_LFInst_4_U21  ( .A1(SubCellInst_LFInst_4_n36 ), .A2(
        SubCellInst_LFInst_4_n35 ), .ZN(MCOutput2[16]) );
  NOR2_X1 SubCellInst_LFInst_4_U20  ( .A1(PermutationOutput[17]), .A2(
        SubCellInst_LFInst_4_n34 ), .ZN(SubCellInst_LFInst_4_n36 ) );
  NOR2_X1 SubCellInst_LFInst_4_U19  ( .A1(SubCellInst_LFInst_4_n33 ), .A2(
        SubCellInst_LFInst_4_n32 ), .ZN(SubCellInst_LFInst_4_n34 ) );
  NOR2_X1 SubCellInst_LFInst_4_U18  ( .A1(PermutationOutput[18]), .A2(
        PermutationOutput[19]), .ZN(SubCellInst_LFInst_4_n32 ) );
  NAND2_X1 SubCellInst_LFInst_4_U17  ( .A1(SubCellInst_LFInst_4_n31 ), .A2(
        SubCellInst_LFInst_4_n30 ), .ZN(MCOutput2[17]) );
  NAND2_X1 SubCellInst_LFInst_4_U16  ( .A1(PermutationOutput[16]), .A2(
        SubCellInst_LFInst_4_n29 ), .ZN(SubCellInst_LFInst_4_n30 ) );
  NAND2_X1 SubCellInst_LFInst_4_U15  ( .A1(PermutationOutput[18]), .A2(
        SubCellInst_LFInst_4_n28 ), .ZN(SubCellInst_LFInst_4_n31 ) );
  NAND2_X1 SubCellInst_LFInst_4_U14  ( .A1(PermutationOutput[19]), .A2(
        SubCellInst_LFInst_4_n33 ), .ZN(SubCellInst_LFInst_4_n28 ) );
  NAND2_X1 SubCellInst_LFInst_4_U13  ( .A1(SubCellInst_LFInst_4_n27 ), .A2(
        SubCellInst_LFInst_4_n26 ), .ZN(MCOutput2[18]) );
  NAND2_X1 SubCellInst_LFInst_4_U12  ( .A1(SubCellInst_LFInst_4_n25 ), .A2(
        PermutationOutput[17]), .ZN(SubCellInst_LFInst_4_n27 ) );
  NAND2_X1 SubCellInst_LFInst_4_U11  ( .A1(SubCellInst_LFInst_4_n24 ), .A2(
        SubCellInst_LFInst_4_n23 ), .ZN(SubCellInst_LFInst_4_n25 ) );
  NAND2_X1 SubCellInst_LFInst_4_U10  ( .A1(PermutationOutput[16]), .A2(
        PermutationOutput[19]), .ZN(SubCellInst_LFInst_4_n24 ) );
  NAND2_X1 SubCellInst_LFInst_4_U9  ( .A1(SubCellInst_LFInst_4_n26 ), .A2(
        SubCellInst_LFInst_4_n22 ), .ZN(MCOutput2[19]) );
  OR2_X1 SubCellInst_LFInst_4_U8  ( .A1(PermutationOutput[17]), .A2(
        SubCellInst_LFInst_4_n35 ), .ZN(SubCellInst_LFInst_4_n22 ) );
  NOR2_X1 SubCellInst_LFInst_4_U7  ( .A1(SubCellInst_LFInst_4_n23 ), .A2(
        SubCellInst_LFInst_4_n29 ), .ZN(SubCellInst_LFInst_4_n35 ) );
  INV_X1 SubCellInst_LFInst_4_U6  ( .A(PermutationOutput[18]), .ZN(
        SubCellInst_LFInst_4_n23 ) );
  NAND2_X1 SubCellInst_LFInst_4_U5  ( .A1(SubCellInst_LFInst_4_n29 ), .A2(
        SubCellInst_LFInst_4_n33 ), .ZN(SubCellInst_LFInst_4_n26 ) );
  INV_X1 SubCellInst_LFInst_4_U4  ( .A(PermutationOutput[16]), .ZN(
        SubCellInst_LFInst_4_n33 ) );
  INV_X1 SubCellInst_LFInst_4_U3  ( .A(PermutationOutput[19]), .ZN(
        SubCellInst_LFInst_4_n29 ) );
  NOR2_X1 SubCellInst_LFInst_5_U21  ( .A1(SubCellInst_LFInst_5_n36 ), .A2(
        SubCellInst_LFInst_5_n35 ), .ZN(MCOutput2[20]) );
  NOR2_X1 SubCellInst_LFInst_5_U20  ( .A1(PermutationOutput[21]), .A2(
        SubCellInst_LFInst_5_n34 ), .ZN(SubCellInst_LFInst_5_n36 ) );
  NOR2_X1 SubCellInst_LFInst_5_U19  ( .A1(SubCellInst_LFInst_5_n33 ), .A2(
        SubCellInst_LFInst_5_n32 ), .ZN(SubCellInst_LFInst_5_n34 ) );
  NOR2_X1 SubCellInst_LFInst_5_U18  ( .A1(PermutationOutput[22]), .A2(
        PermutationOutput[23]), .ZN(SubCellInst_LFInst_5_n32 ) );
  NAND2_X1 SubCellInst_LFInst_5_U17  ( .A1(SubCellInst_LFInst_5_n31 ), .A2(
        SubCellInst_LFInst_5_n30 ), .ZN(MCOutput2[21]) );
  NAND2_X1 SubCellInst_LFInst_5_U16  ( .A1(PermutationOutput[20]), .A2(
        SubCellInst_LFInst_5_n29 ), .ZN(SubCellInst_LFInst_5_n30 ) );
  NAND2_X1 SubCellInst_LFInst_5_U15  ( .A1(PermutationOutput[22]), .A2(
        SubCellInst_LFInst_5_n28 ), .ZN(SubCellInst_LFInst_5_n31 ) );
  NAND2_X1 SubCellInst_LFInst_5_U14  ( .A1(PermutationOutput[23]), .A2(
        SubCellInst_LFInst_5_n33 ), .ZN(SubCellInst_LFInst_5_n28 ) );
  NAND2_X1 SubCellInst_LFInst_5_U13  ( .A1(SubCellInst_LFInst_5_n27 ), .A2(
        SubCellInst_LFInst_5_n26 ), .ZN(MCOutput2[22]) );
  NAND2_X1 SubCellInst_LFInst_5_U12  ( .A1(SubCellInst_LFInst_5_n25 ), .A2(
        PermutationOutput[21]), .ZN(SubCellInst_LFInst_5_n27 ) );
  NAND2_X1 SubCellInst_LFInst_5_U11  ( .A1(SubCellInst_LFInst_5_n24 ), .A2(
        SubCellInst_LFInst_5_n23 ), .ZN(SubCellInst_LFInst_5_n25 ) );
  NAND2_X1 SubCellInst_LFInst_5_U10  ( .A1(PermutationOutput[20]), .A2(
        PermutationOutput[23]), .ZN(SubCellInst_LFInst_5_n24 ) );
  NAND2_X1 SubCellInst_LFInst_5_U9  ( .A1(SubCellInst_LFInst_5_n26 ), .A2(
        SubCellInst_LFInst_5_n22 ), .ZN(MCOutput2[23]) );
  OR2_X1 SubCellInst_LFInst_5_U8  ( .A1(PermutationOutput[21]), .A2(
        SubCellInst_LFInst_5_n35 ), .ZN(SubCellInst_LFInst_5_n22 ) );
  NOR2_X1 SubCellInst_LFInst_5_U7  ( .A1(SubCellInst_LFInst_5_n23 ), .A2(
        SubCellInst_LFInst_5_n29 ), .ZN(SubCellInst_LFInst_5_n35 ) );
  INV_X1 SubCellInst_LFInst_5_U6  ( .A(PermutationOutput[22]), .ZN(
        SubCellInst_LFInst_5_n23 ) );
  NAND2_X1 SubCellInst_LFInst_5_U5  ( .A1(SubCellInst_LFInst_5_n29 ), .A2(
        SubCellInst_LFInst_5_n33 ), .ZN(SubCellInst_LFInst_5_n26 ) );
  INV_X1 SubCellInst_LFInst_5_U4  ( .A(PermutationOutput[20]), .ZN(
        SubCellInst_LFInst_5_n33 ) );
  INV_X1 SubCellInst_LFInst_5_U3  ( .A(PermutationOutput[23]), .ZN(
        SubCellInst_LFInst_5_n29 ) );
  NOR2_X1 SubCellInst_LFInst_6_U21  ( .A1(SubCellInst_LFInst_6_n36 ), .A2(
        SubCellInst_LFInst_6_n35 ), .ZN(MCOutput2[24]) );
  NOR2_X1 SubCellInst_LFInst_6_U20  ( .A1(PermutationOutput[25]), .A2(
        SubCellInst_LFInst_6_n34 ), .ZN(SubCellInst_LFInst_6_n36 ) );
  NOR2_X1 SubCellInst_LFInst_6_U19  ( .A1(SubCellInst_LFInst_6_n33 ), .A2(
        SubCellInst_LFInst_6_n32 ), .ZN(SubCellInst_LFInst_6_n34 ) );
  NOR2_X1 SubCellInst_LFInst_6_U18  ( .A1(PermutationOutput[26]), .A2(
        PermutationOutput[27]), .ZN(SubCellInst_LFInst_6_n32 ) );
  NAND2_X1 SubCellInst_LFInst_6_U17  ( .A1(SubCellInst_LFInst_6_n31 ), .A2(
        SubCellInst_LFInst_6_n30 ), .ZN(MCOutput2[25]) );
  NAND2_X1 SubCellInst_LFInst_6_U16  ( .A1(PermutationOutput[24]), .A2(
        SubCellInst_LFInst_6_n29 ), .ZN(SubCellInst_LFInst_6_n30 ) );
  NAND2_X1 SubCellInst_LFInst_6_U15  ( .A1(PermutationOutput[26]), .A2(
        SubCellInst_LFInst_6_n28 ), .ZN(SubCellInst_LFInst_6_n31 ) );
  NAND2_X1 SubCellInst_LFInst_6_U14  ( .A1(PermutationOutput[27]), .A2(
        SubCellInst_LFInst_6_n33 ), .ZN(SubCellInst_LFInst_6_n28 ) );
  NAND2_X1 SubCellInst_LFInst_6_U13  ( .A1(SubCellInst_LFInst_6_n27 ), .A2(
        SubCellInst_LFInst_6_n26 ), .ZN(MCOutput2[26]) );
  NAND2_X1 SubCellInst_LFInst_6_U12  ( .A1(SubCellInst_LFInst_6_n25 ), .A2(
        PermutationOutput[25]), .ZN(SubCellInst_LFInst_6_n27 ) );
  NAND2_X1 SubCellInst_LFInst_6_U11  ( .A1(SubCellInst_LFInst_6_n24 ), .A2(
        SubCellInst_LFInst_6_n23 ), .ZN(SubCellInst_LFInst_6_n25 ) );
  NAND2_X1 SubCellInst_LFInst_6_U10  ( .A1(PermutationOutput[24]), .A2(
        PermutationOutput[27]), .ZN(SubCellInst_LFInst_6_n24 ) );
  NAND2_X1 SubCellInst_LFInst_6_U9  ( .A1(SubCellInst_LFInst_6_n26 ), .A2(
        SubCellInst_LFInst_6_n22 ), .ZN(MCOutput2[27]) );
  OR2_X1 SubCellInst_LFInst_6_U8  ( .A1(PermutationOutput[25]), .A2(
        SubCellInst_LFInst_6_n35 ), .ZN(SubCellInst_LFInst_6_n22 ) );
  NOR2_X1 SubCellInst_LFInst_6_U7  ( .A1(SubCellInst_LFInst_6_n23 ), .A2(
        SubCellInst_LFInst_6_n29 ), .ZN(SubCellInst_LFInst_6_n35 ) );
  INV_X1 SubCellInst_LFInst_6_U6  ( .A(PermutationOutput[26]), .ZN(
        SubCellInst_LFInst_6_n23 ) );
  NAND2_X1 SubCellInst_LFInst_6_U5  ( .A1(SubCellInst_LFInst_6_n29 ), .A2(
        SubCellInst_LFInst_6_n33 ), .ZN(SubCellInst_LFInst_6_n26 ) );
  INV_X1 SubCellInst_LFInst_6_U4  ( .A(PermutationOutput[24]), .ZN(
        SubCellInst_LFInst_6_n33 ) );
  INV_X1 SubCellInst_LFInst_6_U3  ( .A(PermutationOutput[27]), .ZN(
        SubCellInst_LFInst_6_n29 ) );
  NOR2_X1 SubCellInst_LFInst_7_U21  ( .A1(SubCellInst_LFInst_7_n36 ), .A2(
        SubCellInst_LFInst_7_n35 ), .ZN(MCOutput2[28]) );
  NOR2_X1 SubCellInst_LFInst_7_U20  ( .A1(PermutationOutput[29]), .A2(
        SubCellInst_LFInst_7_n34 ), .ZN(SubCellInst_LFInst_7_n36 ) );
  NOR2_X1 SubCellInst_LFInst_7_U19  ( .A1(SubCellInst_LFInst_7_n33 ), .A2(
        SubCellInst_LFInst_7_n32 ), .ZN(SubCellInst_LFInst_7_n34 ) );
  NOR2_X1 SubCellInst_LFInst_7_U18  ( .A1(PermutationOutput[30]), .A2(
        PermutationOutput[31]), .ZN(SubCellInst_LFInst_7_n32 ) );
  NAND2_X1 SubCellInst_LFInst_7_U17  ( .A1(SubCellInst_LFInst_7_n31 ), .A2(
        SubCellInst_LFInst_7_n30 ), .ZN(MCOutput2[29]) );
  NAND2_X1 SubCellInst_LFInst_7_U16  ( .A1(PermutationOutput[28]), .A2(
        SubCellInst_LFInst_7_n29 ), .ZN(SubCellInst_LFInst_7_n30 ) );
  NAND2_X1 SubCellInst_LFInst_7_U15  ( .A1(PermutationOutput[30]), .A2(
        SubCellInst_LFInst_7_n28 ), .ZN(SubCellInst_LFInst_7_n31 ) );
  NAND2_X1 SubCellInst_LFInst_7_U14  ( .A1(PermutationOutput[31]), .A2(
        SubCellInst_LFInst_7_n33 ), .ZN(SubCellInst_LFInst_7_n28 ) );
  NAND2_X1 SubCellInst_LFInst_7_U13  ( .A1(SubCellInst_LFInst_7_n27 ), .A2(
        SubCellInst_LFInst_7_n26 ), .ZN(MCOutput2[30]) );
  NAND2_X1 SubCellInst_LFInst_7_U12  ( .A1(SubCellInst_LFInst_7_n25 ), .A2(
        PermutationOutput[29]), .ZN(SubCellInst_LFInst_7_n27 ) );
  NAND2_X1 SubCellInst_LFInst_7_U11  ( .A1(SubCellInst_LFInst_7_n24 ), .A2(
        SubCellInst_LFInst_7_n23 ), .ZN(SubCellInst_LFInst_7_n25 ) );
  NAND2_X1 SubCellInst_LFInst_7_U10  ( .A1(PermutationOutput[28]), .A2(
        PermutationOutput[31]), .ZN(SubCellInst_LFInst_7_n24 ) );
  NAND2_X1 SubCellInst_LFInst_7_U9  ( .A1(SubCellInst_LFInst_7_n26 ), .A2(
        SubCellInst_LFInst_7_n22 ), .ZN(MCOutput2[31]) );
  OR2_X1 SubCellInst_LFInst_7_U8  ( .A1(PermutationOutput[29]), .A2(
        SubCellInst_LFInst_7_n35 ), .ZN(SubCellInst_LFInst_7_n22 ) );
  NOR2_X1 SubCellInst_LFInst_7_U7  ( .A1(SubCellInst_LFInst_7_n23 ), .A2(
        SubCellInst_LFInst_7_n29 ), .ZN(SubCellInst_LFInst_7_n35 ) );
  INV_X1 SubCellInst_LFInst_7_U6  ( .A(PermutationOutput[30]), .ZN(
        SubCellInst_LFInst_7_n23 ) );
  NAND2_X1 SubCellInst_LFInst_7_U5  ( .A1(SubCellInst_LFInst_7_n29 ), .A2(
        SubCellInst_LFInst_7_n33 ), .ZN(SubCellInst_LFInst_7_n26 ) );
  INV_X1 SubCellInst_LFInst_7_U4  ( .A(PermutationOutput[28]), .ZN(
        SubCellInst_LFInst_7_n33 ) );
  INV_X1 SubCellInst_LFInst_7_U3  ( .A(PermutationOutput[31]), .ZN(
        SubCellInst_LFInst_7_n29 ) );
  NOR2_X1 SubCellInst_LFInst_8_U21  ( .A1(SubCellInst_LFInst_8_n36 ), .A2(
        SubCellInst_LFInst_8_n35 ), .ZN(Feedback[32]) );
  NOR2_X1 SubCellInst_LFInst_8_U20  ( .A1(PermutationOutput[33]), .A2(
        SubCellInst_LFInst_8_n34 ), .ZN(SubCellInst_LFInst_8_n36 ) );
  NOR2_X1 SubCellInst_LFInst_8_U19  ( .A1(SubCellInst_LFInst_8_n33 ), .A2(
        SubCellInst_LFInst_8_n32 ), .ZN(SubCellInst_LFInst_8_n34 ) );
  NOR2_X1 SubCellInst_LFInst_8_U18  ( .A1(PermutationOutput[34]), .A2(
        PermutationOutput[35]), .ZN(SubCellInst_LFInst_8_n32 ) );
  NAND2_X1 SubCellInst_LFInst_8_U17  ( .A1(SubCellInst_LFInst_8_n31 ), .A2(
        SubCellInst_LFInst_8_n30 ), .ZN(Feedback[33]) );
  NAND2_X1 SubCellInst_LFInst_8_U16  ( .A1(PermutationOutput[32]), .A2(
        SubCellInst_LFInst_8_n29 ), .ZN(SubCellInst_LFInst_8_n30 ) );
  NAND2_X1 SubCellInst_LFInst_8_U15  ( .A1(PermutationOutput[34]), .A2(
        SubCellInst_LFInst_8_n28 ), .ZN(SubCellInst_LFInst_8_n31 ) );
  NAND2_X1 SubCellInst_LFInst_8_U14  ( .A1(PermutationOutput[35]), .A2(
        SubCellInst_LFInst_8_n33 ), .ZN(SubCellInst_LFInst_8_n28 ) );
  NAND2_X1 SubCellInst_LFInst_8_U13  ( .A1(SubCellInst_LFInst_8_n27 ), .A2(
        SubCellInst_LFInst_8_n26 ), .ZN(Feedback[34]) );
  NAND2_X1 SubCellInst_LFInst_8_U12  ( .A1(SubCellInst_LFInst_8_n25 ), .A2(
        PermutationOutput[33]), .ZN(SubCellInst_LFInst_8_n27 ) );
  NAND2_X1 SubCellInst_LFInst_8_U11  ( .A1(SubCellInst_LFInst_8_n24 ), .A2(
        SubCellInst_LFInst_8_n23 ), .ZN(SubCellInst_LFInst_8_n25 ) );
  NAND2_X1 SubCellInst_LFInst_8_U10  ( .A1(PermutationOutput[32]), .A2(
        PermutationOutput[35]), .ZN(SubCellInst_LFInst_8_n24 ) );
  NAND2_X1 SubCellInst_LFInst_8_U9  ( .A1(SubCellInst_LFInst_8_n26 ), .A2(
        SubCellInst_LFInst_8_n22 ), .ZN(Feedback[35]) );
  OR2_X1 SubCellInst_LFInst_8_U8  ( .A1(PermutationOutput[33]), .A2(
        SubCellInst_LFInst_8_n35 ), .ZN(SubCellInst_LFInst_8_n22 ) );
  NOR2_X1 SubCellInst_LFInst_8_U7  ( .A1(SubCellInst_LFInst_8_n23 ), .A2(
        SubCellInst_LFInst_8_n29 ), .ZN(SubCellInst_LFInst_8_n35 ) );
  INV_X1 SubCellInst_LFInst_8_U6  ( .A(PermutationOutput[34]), .ZN(
        SubCellInst_LFInst_8_n23 ) );
  NAND2_X1 SubCellInst_LFInst_8_U5  ( .A1(SubCellInst_LFInst_8_n29 ), .A2(
        SubCellInst_LFInst_8_n33 ), .ZN(SubCellInst_LFInst_8_n26 ) );
  INV_X1 SubCellInst_LFInst_8_U4  ( .A(PermutationOutput[32]), .ZN(
        SubCellInst_LFInst_8_n33 ) );
  INV_X1 SubCellInst_LFInst_8_U3  ( .A(PermutationOutput[35]), .ZN(
        SubCellInst_LFInst_8_n29 ) );
  NOR2_X1 SubCellInst_LFInst_9_U21  ( .A1(SubCellInst_LFInst_9_n36 ), .A2(
        SubCellInst_LFInst_9_n35 ), .ZN(Feedback[36]) );
  NOR2_X1 SubCellInst_LFInst_9_U20  ( .A1(PermutationOutput[37]), .A2(
        SubCellInst_LFInst_9_n34 ), .ZN(SubCellInst_LFInst_9_n36 ) );
  NOR2_X1 SubCellInst_LFInst_9_U19  ( .A1(SubCellInst_LFInst_9_n33 ), .A2(
        SubCellInst_LFInst_9_n32 ), .ZN(SubCellInst_LFInst_9_n34 ) );
  NOR2_X1 SubCellInst_LFInst_9_U18  ( .A1(PermutationOutput[38]), .A2(
        PermutationOutput[39]), .ZN(SubCellInst_LFInst_9_n32 ) );
  NAND2_X1 SubCellInst_LFInst_9_U17  ( .A1(SubCellInst_LFInst_9_n31 ), .A2(
        SubCellInst_LFInst_9_n30 ), .ZN(Feedback[37]) );
  NAND2_X1 SubCellInst_LFInst_9_U16  ( .A1(PermutationOutput[36]), .A2(
        SubCellInst_LFInst_9_n29 ), .ZN(SubCellInst_LFInst_9_n30 ) );
  NAND2_X1 SubCellInst_LFInst_9_U15  ( .A1(PermutationOutput[38]), .A2(
        SubCellInst_LFInst_9_n28 ), .ZN(SubCellInst_LFInst_9_n31 ) );
  NAND2_X1 SubCellInst_LFInst_9_U14  ( .A1(PermutationOutput[39]), .A2(
        SubCellInst_LFInst_9_n33 ), .ZN(SubCellInst_LFInst_9_n28 ) );
  NAND2_X1 SubCellInst_LFInst_9_U13  ( .A1(SubCellInst_LFInst_9_n27 ), .A2(
        SubCellInst_LFInst_9_n26 ), .ZN(Feedback[38]) );
  NAND2_X1 SubCellInst_LFInst_9_U12  ( .A1(SubCellInst_LFInst_9_n25 ), .A2(
        PermutationOutput[37]), .ZN(SubCellInst_LFInst_9_n27 ) );
  NAND2_X1 SubCellInst_LFInst_9_U11  ( .A1(SubCellInst_LFInst_9_n24 ), .A2(
        SubCellInst_LFInst_9_n23 ), .ZN(SubCellInst_LFInst_9_n25 ) );
  NAND2_X1 SubCellInst_LFInst_9_U10  ( .A1(PermutationOutput[36]), .A2(
        PermutationOutput[39]), .ZN(SubCellInst_LFInst_9_n24 ) );
  NAND2_X1 SubCellInst_LFInst_9_U9  ( .A1(SubCellInst_LFInst_9_n26 ), .A2(
        SubCellInst_LFInst_9_n22 ), .ZN(Feedback[39]) );
  OR2_X1 SubCellInst_LFInst_9_U8  ( .A1(PermutationOutput[37]), .A2(
        SubCellInst_LFInst_9_n35 ), .ZN(SubCellInst_LFInst_9_n22 ) );
  NOR2_X1 SubCellInst_LFInst_9_U7  ( .A1(SubCellInst_LFInst_9_n23 ), .A2(
        SubCellInst_LFInst_9_n29 ), .ZN(SubCellInst_LFInst_9_n35 ) );
  INV_X1 SubCellInst_LFInst_9_U6  ( .A(PermutationOutput[38]), .ZN(
        SubCellInst_LFInst_9_n23 ) );
  NAND2_X1 SubCellInst_LFInst_9_U5  ( .A1(SubCellInst_LFInst_9_n29 ), .A2(
        SubCellInst_LFInst_9_n33 ), .ZN(SubCellInst_LFInst_9_n26 ) );
  INV_X1 SubCellInst_LFInst_9_U4  ( .A(PermutationOutput[36]), .ZN(
        SubCellInst_LFInst_9_n33 ) );
  INV_X1 SubCellInst_LFInst_9_U3  ( .A(PermutationOutput[39]), .ZN(
        SubCellInst_LFInst_9_n29 ) );
  NOR2_X1 SubCellInst_LFInst_10_U21  ( .A1(SubCellInst_LFInst_10_n36 ), .A2(
        SubCellInst_LFInst_10_n35 ), .ZN(Feedback[40]) );
  NOR2_X1 SubCellInst_LFInst_10_U20  ( .A1(PermutationOutput[41]), .A2(
        SubCellInst_LFInst_10_n34 ), .ZN(SubCellInst_LFInst_10_n36 ) );
  NOR2_X1 SubCellInst_LFInst_10_U19  ( .A1(SubCellInst_LFInst_10_n33 ), .A2(
        SubCellInst_LFInst_10_n32 ), .ZN(SubCellInst_LFInst_10_n34 ) );
  NOR2_X1 SubCellInst_LFInst_10_U18  ( .A1(PermutationOutput[42]), .A2(
        PermutationOutput[43]), .ZN(SubCellInst_LFInst_10_n32 ) );
  NAND2_X1 SubCellInst_LFInst_10_U17  ( .A1(SubCellInst_LFInst_10_n31 ), 
        .A2(SubCellInst_LFInst_10_n30 ), .ZN(Feedback[41]) );
  NAND2_X1 SubCellInst_LFInst_10_U16  ( .A1(PermutationOutput[40]), .A2(
        SubCellInst_LFInst_10_n29 ), .ZN(SubCellInst_LFInst_10_n30 ) );
  NAND2_X1 SubCellInst_LFInst_10_U15  ( .A1(PermutationOutput[42]), .A2(
        SubCellInst_LFInst_10_n28 ), .ZN(SubCellInst_LFInst_10_n31 ) );
  NAND2_X1 SubCellInst_LFInst_10_U14  ( .A1(PermutationOutput[43]), .A2(
        SubCellInst_LFInst_10_n33 ), .ZN(SubCellInst_LFInst_10_n28 ) );
  NAND2_X1 SubCellInst_LFInst_10_U13  ( .A1(SubCellInst_LFInst_10_n27 ), 
        .A2(SubCellInst_LFInst_10_n26 ), .ZN(Feedback[42]) );
  NAND2_X1 SubCellInst_LFInst_10_U12  ( .A1(SubCellInst_LFInst_10_n25 ), 
        .A2(PermutationOutput[41]), .ZN(SubCellInst_LFInst_10_n27 ) );
  NAND2_X1 SubCellInst_LFInst_10_U11  ( .A1(SubCellInst_LFInst_10_n24 ), 
        .A2(SubCellInst_LFInst_10_n23 ), .ZN(SubCellInst_LFInst_10_n25 ) );
  NAND2_X1 SubCellInst_LFInst_10_U10  ( .A1(PermutationOutput[40]), .A2(
        PermutationOutput[43]), .ZN(SubCellInst_LFInst_10_n24 ) );
  NAND2_X1 SubCellInst_LFInst_10_U9  ( .A1(SubCellInst_LFInst_10_n26 ), .A2(
        SubCellInst_LFInst_10_n22 ), .ZN(Feedback[43]) );
  OR2_X1 SubCellInst_LFInst_10_U8  ( .A1(PermutationOutput[41]), .A2(
        SubCellInst_LFInst_10_n35 ), .ZN(SubCellInst_LFInst_10_n22 ) );
  NOR2_X1 SubCellInst_LFInst_10_U7  ( .A1(SubCellInst_LFInst_10_n23 ), .A2(
        SubCellInst_LFInst_10_n29 ), .ZN(SubCellInst_LFInst_10_n35 ) );
  INV_X1 SubCellInst_LFInst_10_U6  ( .A(PermutationOutput[42]), .ZN(
        SubCellInst_LFInst_10_n23 ) );
  NAND2_X1 SubCellInst_LFInst_10_U5  ( .A1(SubCellInst_LFInst_10_n29 ), .A2(
        SubCellInst_LFInst_10_n33 ), .ZN(SubCellInst_LFInst_10_n26 ) );
  INV_X1 SubCellInst_LFInst_10_U4  ( .A(PermutationOutput[40]), .ZN(
        SubCellInst_LFInst_10_n33 ) );
  INV_X1 SubCellInst_LFInst_10_U3  ( .A(PermutationOutput[43]), .ZN(
        SubCellInst_LFInst_10_n29 ) );
  NOR2_X1 SubCellInst_LFInst_11_U21  ( .A1(SubCellInst_LFInst_11_n36 ), .A2(
        SubCellInst_LFInst_11_n35 ), .ZN(Feedback[44]) );
  NOR2_X1 SubCellInst_LFInst_11_U20  ( .A1(PermutationOutput[45]), .A2(
        SubCellInst_LFInst_11_n34 ), .ZN(SubCellInst_LFInst_11_n36 ) );
  NOR2_X1 SubCellInst_LFInst_11_U19  ( .A1(SubCellInst_LFInst_11_n33 ), .A2(
        SubCellInst_LFInst_11_n32 ), .ZN(SubCellInst_LFInst_11_n34 ) );
  NOR2_X1 SubCellInst_LFInst_11_U18  ( .A1(PermutationOutput[46]), .A2(
        PermutationOutput[47]), .ZN(SubCellInst_LFInst_11_n32 ) );
  NAND2_X1 SubCellInst_LFInst_11_U17  ( .A1(SubCellInst_LFInst_11_n31 ), 
        .A2(SubCellInst_LFInst_11_n30 ), .ZN(Feedback[45]) );
  NAND2_X1 SubCellInst_LFInst_11_U16  ( .A1(PermutationOutput[44]), .A2(
        SubCellInst_LFInst_11_n29 ), .ZN(SubCellInst_LFInst_11_n30 ) );
  NAND2_X1 SubCellInst_LFInst_11_U15  ( .A1(PermutationOutput[46]), .A2(
        SubCellInst_LFInst_11_n28 ), .ZN(SubCellInst_LFInst_11_n31 ) );
  NAND2_X1 SubCellInst_LFInst_11_U14  ( .A1(PermutationOutput[47]), .A2(
        SubCellInst_LFInst_11_n33 ), .ZN(SubCellInst_LFInst_11_n28 ) );
  NAND2_X1 SubCellInst_LFInst_11_U13  ( .A1(SubCellInst_LFInst_11_n27 ), 
        .A2(SubCellInst_LFInst_11_n26 ), .ZN(Feedback[46]) );
  NAND2_X1 SubCellInst_LFInst_11_U12  ( .A1(SubCellInst_LFInst_11_n25 ), 
        .A2(PermutationOutput[45]), .ZN(SubCellInst_LFInst_11_n27 ) );
  NAND2_X1 SubCellInst_LFInst_11_U11  ( .A1(SubCellInst_LFInst_11_n24 ), 
        .A2(SubCellInst_LFInst_11_n23 ), .ZN(SubCellInst_LFInst_11_n25 ) );
  NAND2_X1 SubCellInst_LFInst_11_U10  ( .A1(PermutationOutput[44]), .A2(
        PermutationOutput[47]), .ZN(SubCellInst_LFInst_11_n24 ) );
  NAND2_X1 SubCellInst_LFInst_11_U9  ( .A1(SubCellInst_LFInst_11_n26 ), .A2(
        SubCellInst_LFInst_11_n22 ), .ZN(Feedback[47]) );
  OR2_X1 SubCellInst_LFInst_11_U8  ( .A1(PermutationOutput[45]), .A2(
        SubCellInst_LFInst_11_n35 ), .ZN(SubCellInst_LFInst_11_n22 ) );
  NOR2_X1 SubCellInst_LFInst_11_U7  ( .A1(SubCellInst_LFInst_11_n23 ), .A2(
        SubCellInst_LFInst_11_n29 ), .ZN(SubCellInst_LFInst_11_n35 ) );
  INV_X1 SubCellInst_LFInst_11_U6  ( .A(PermutationOutput[46]), .ZN(
        SubCellInst_LFInst_11_n23 ) );
  NAND2_X1 SubCellInst_LFInst_11_U5  ( .A1(SubCellInst_LFInst_11_n29 ), .A2(
        SubCellInst_LFInst_11_n33 ), .ZN(SubCellInst_LFInst_11_n26 ) );
  INV_X1 SubCellInst_LFInst_11_U4  ( .A(PermutationOutput[44]), .ZN(
        SubCellInst_LFInst_11_n33 ) );
  INV_X1 SubCellInst_LFInst_11_U3  ( .A(PermutationOutput[47]), .ZN(
        SubCellInst_LFInst_11_n29 ) );
  NOR2_X1 SubCellInst_LFInst_12_U21  ( .A1(SubCellInst_LFInst_12_n36 ), .A2(
        SubCellInst_LFInst_12_n35 ), .ZN(Feedback[48]) );
  NOR2_X1 SubCellInst_LFInst_12_U20  ( .A1(PermutationOutput[49]), .A2(
        SubCellInst_LFInst_12_n34 ), .ZN(SubCellInst_LFInst_12_n36 ) );
  NOR2_X1 SubCellInst_LFInst_12_U19  ( .A1(SubCellInst_LFInst_12_n33 ), .A2(
        SubCellInst_LFInst_12_n32 ), .ZN(SubCellInst_LFInst_12_n34 ) );
  NOR2_X1 SubCellInst_LFInst_12_U18  ( .A1(PermutationOutput[50]), .A2(
        PermutationOutput[51]), .ZN(SubCellInst_LFInst_12_n32 ) );
  NAND2_X1 SubCellInst_LFInst_12_U17  ( .A1(SubCellInst_LFInst_12_n31 ), 
        .A2(SubCellInst_LFInst_12_n30 ), .ZN(Feedback[49]) );
  NAND2_X1 SubCellInst_LFInst_12_U16  ( .A1(PermutationOutput[48]), .A2(
        SubCellInst_LFInst_12_n29 ), .ZN(SubCellInst_LFInst_12_n30 ) );
  NAND2_X1 SubCellInst_LFInst_12_U15  ( .A1(PermutationOutput[50]), .A2(
        SubCellInst_LFInst_12_n28 ), .ZN(SubCellInst_LFInst_12_n31 ) );
  NAND2_X1 SubCellInst_LFInst_12_U14  ( .A1(PermutationOutput[51]), .A2(
        SubCellInst_LFInst_12_n33 ), .ZN(SubCellInst_LFInst_12_n28 ) );
  NAND2_X1 SubCellInst_LFInst_12_U13  ( .A1(SubCellInst_LFInst_12_n27 ), 
        .A2(SubCellInst_LFInst_12_n26 ), .ZN(Feedback[50]) );
  NAND2_X1 SubCellInst_LFInst_12_U12  ( .A1(SubCellInst_LFInst_12_n25 ), 
        .A2(PermutationOutput[49]), .ZN(SubCellInst_LFInst_12_n27 ) );
  NAND2_X1 SubCellInst_LFInst_12_U11  ( .A1(SubCellInst_LFInst_12_n24 ), 
        .A2(SubCellInst_LFInst_12_n23 ), .ZN(SubCellInst_LFInst_12_n25 ) );
  NAND2_X1 SubCellInst_LFInst_12_U10  ( .A1(PermutationOutput[48]), .A2(
        PermutationOutput[51]), .ZN(SubCellInst_LFInst_12_n24 ) );
  NAND2_X1 SubCellInst_LFInst_12_U9  ( .A1(SubCellInst_LFInst_12_n26 ), .A2(
        SubCellInst_LFInst_12_n22 ), .ZN(Feedback[51]) );
  OR2_X1 SubCellInst_LFInst_12_U8  ( .A1(PermutationOutput[49]), .A2(
        SubCellInst_LFInst_12_n35 ), .ZN(SubCellInst_LFInst_12_n22 ) );
  NOR2_X1 SubCellInst_LFInst_12_U7  ( .A1(SubCellInst_LFInst_12_n23 ), .A2(
        SubCellInst_LFInst_12_n29 ), .ZN(SubCellInst_LFInst_12_n35 ) );
  INV_X1 SubCellInst_LFInst_12_U6  ( .A(PermutationOutput[50]), .ZN(
        SubCellInst_LFInst_12_n23 ) );
  NAND2_X1 SubCellInst_LFInst_12_U5  ( .A1(SubCellInst_LFInst_12_n29 ), .A2(
        SubCellInst_LFInst_12_n33 ), .ZN(SubCellInst_LFInst_12_n26 ) );
  INV_X1 SubCellInst_LFInst_12_U4  ( .A(PermutationOutput[48]), .ZN(
        SubCellInst_LFInst_12_n33 ) );
  INV_X1 SubCellInst_LFInst_12_U3  ( .A(PermutationOutput[51]), .ZN(
        SubCellInst_LFInst_12_n29 ) );
  NOR2_X1 SubCellInst_LFInst_13_U21  ( .A1(SubCellInst_LFInst_13_n36 ), .A2(
        SubCellInst_LFInst_13_n35 ), .ZN(Feedback[52]) );
  NOR2_X1 SubCellInst_LFInst_13_U20  ( .A1(PermutationOutput[53]), .A2(
        SubCellInst_LFInst_13_n34 ), .ZN(SubCellInst_LFInst_13_n36 ) );
  NOR2_X1 SubCellInst_LFInst_13_U19  ( .A1(SubCellInst_LFInst_13_n33 ), .A2(
        SubCellInst_LFInst_13_n32 ), .ZN(SubCellInst_LFInst_13_n34 ) );
  NOR2_X1 SubCellInst_LFInst_13_U18  ( .A1(PermutationOutput[54]), .A2(
        PermutationOutput[55]), .ZN(SubCellInst_LFInst_13_n32 ) );
  NAND2_X1 SubCellInst_LFInst_13_U17  ( .A1(SubCellInst_LFInst_13_n31 ), 
        .A2(SubCellInst_LFInst_13_n30 ), .ZN(Feedback[53]) );
  NAND2_X1 SubCellInst_LFInst_13_U16  ( .A1(PermutationOutput[52]), .A2(
        SubCellInst_LFInst_13_n29 ), .ZN(SubCellInst_LFInst_13_n30 ) );
  NAND2_X1 SubCellInst_LFInst_13_U15  ( .A1(PermutationOutput[54]), .A2(
        SubCellInst_LFInst_13_n28 ), .ZN(SubCellInst_LFInst_13_n31 ) );
  NAND2_X1 SubCellInst_LFInst_13_U14  ( .A1(PermutationOutput[55]), .A2(
        SubCellInst_LFInst_13_n33 ), .ZN(SubCellInst_LFInst_13_n28 ) );
  NAND2_X1 SubCellInst_LFInst_13_U13  ( .A1(SubCellInst_LFInst_13_n27 ), 
        .A2(SubCellInst_LFInst_13_n26 ), .ZN(Feedback[54]) );
  NAND2_X1 SubCellInst_LFInst_13_U12  ( .A1(SubCellInst_LFInst_13_n25 ), 
        .A2(PermutationOutput[53]), .ZN(SubCellInst_LFInst_13_n27 ) );
  NAND2_X1 SubCellInst_LFInst_13_U11  ( .A1(SubCellInst_LFInst_13_n24 ), 
        .A2(SubCellInst_LFInst_13_n23 ), .ZN(SubCellInst_LFInst_13_n25 ) );
  NAND2_X1 SubCellInst_LFInst_13_U10  ( .A1(PermutationOutput[52]), .A2(
        PermutationOutput[55]), .ZN(SubCellInst_LFInst_13_n24 ) );
  NAND2_X1 SubCellInst_LFInst_13_U9  ( .A1(SubCellInst_LFInst_13_n26 ), .A2(
        SubCellInst_LFInst_13_n22 ), .ZN(Feedback[55]) );
  OR2_X1 SubCellInst_LFInst_13_U8  ( .A1(PermutationOutput[53]), .A2(
        SubCellInst_LFInst_13_n35 ), .ZN(SubCellInst_LFInst_13_n22 ) );
  NOR2_X1 SubCellInst_LFInst_13_U7  ( .A1(SubCellInst_LFInst_13_n23 ), .A2(
        SubCellInst_LFInst_13_n29 ), .ZN(SubCellInst_LFInst_13_n35 ) );
  INV_X1 SubCellInst_LFInst_13_U6  ( .A(PermutationOutput[54]), .ZN(
        SubCellInst_LFInst_13_n23 ) );
  NAND2_X1 SubCellInst_LFInst_13_U5  ( .A1(SubCellInst_LFInst_13_n29 ), .A2(
        SubCellInst_LFInst_13_n33 ), .ZN(SubCellInst_LFInst_13_n26 ) );
  INV_X1 SubCellInst_LFInst_13_U4  ( .A(PermutationOutput[52]), .ZN(
        SubCellInst_LFInst_13_n33 ) );
  INV_X1 SubCellInst_LFInst_13_U3  ( .A(PermutationOutput[55]), .ZN(
        SubCellInst_LFInst_13_n29 ) );
  NOR2_X1 SubCellInst_LFInst_14_U21  ( .A1(SubCellInst_LFInst_14_n36 ), .A2(
        SubCellInst_LFInst_14_n35 ), .ZN(Feedback[56]) );
  NOR2_X1 SubCellInst_LFInst_14_U20  ( .A1(PermutationOutput[57]), .A2(
        SubCellInst_LFInst_14_n34 ), .ZN(SubCellInst_LFInst_14_n36 ) );
  NOR2_X1 SubCellInst_LFInst_14_U19  ( .A1(SubCellInst_LFInst_14_n33 ), .A2(
        SubCellInst_LFInst_14_n32 ), .ZN(SubCellInst_LFInst_14_n34 ) );
  NOR2_X1 SubCellInst_LFInst_14_U18  ( .A1(PermutationOutput[58]), .A2(
        PermutationOutput[59]), .ZN(SubCellInst_LFInst_14_n32 ) );
  NAND2_X1 SubCellInst_LFInst_14_U17  ( .A1(SubCellInst_LFInst_14_n31 ), 
        .A2(SubCellInst_LFInst_14_n30 ), .ZN(Feedback[57]) );
  NAND2_X1 SubCellInst_LFInst_14_U16  ( .A1(PermutationOutput[56]), .A2(
        SubCellInst_LFInst_14_n29 ), .ZN(SubCellInst_LFInst_14_n30 ) );
  NAND2_X1 SubCellInst_LFInst_14_U15  ( .A1(PermutationOutput[58]), .A2(
        SubCellInst_LFInst_14_n28 ), .ZN(SubCellInst_LFInst_14_n31 ) );
  NAND2_X1 SubCellInst_LFInst_14_U14  ( .A1(PermutationOutput[59]), .A2(
        SubCellInst_LFInst_14_n33 ), .ZN(SubCellInst_LFInst_14_n28 ) );
  NAND2_X1 SubCellInst_LFInst_14_U13  ( .A1(SubCellInst_LFInst_14_n27 ), 
        .A2(SubCellInst_LFInst_14_n26 ), .ZN(Feedback[58]) );
  NAND2_X1 SubCellInst_LFInst_14_U12  ( .A1(SubCellInst_LFInst_14_n25 ), 
        .A2(PermutationOutput[57]), .ZN(SubCellInst_LFInst_14_n27 ) );
  NAND2_X1 SubCellInst_LFInst_14_U11  ( .A1(SubCellInst_LFInst_14_n24 ), 
        .A2(SubCellInst_LFInst_14_n23 ), .ZN(SubCellInst_LFInst_14_n25 ) );
  NAND2_X1 SubCellInst_LFInst_14_U10  ( .A1(PermutationOutput[56]), .A2(
        PermutationOutput[59]), .ZN(SubCellInst_LFInst_14_n24 ) );
  NAND2_X1 SubCellInst_LFInst_14_U9  ( .A1(SubCellInst_LFInst_14_n26 ), .A2(
        SubCellInst_LFInst_14_n22 ), .ZN(Feedback[59]) );
  OR2_X1 SubCellInst_LFInst_14_U8  ( .A1(PermutationOutput[57]), .A2(
        SubCellInst_LFInst_14_n35 ), .ZN(SubCellInst_LFInst_14_n22 ) );
  NOR2_X1 SubCellInst_LFInst_14_U7  ( .A1(SubCellInst_LFInst_14_n23 ), .A2(
        SubCellInst_LFInst_14_n29 ), .ZN(SubCellInst_LFInst_14_n35 ) );
  INV_X1 SubCellInst_LFInst_14_U6  ( .A(PermutationOutput[58]), .ZN(
        SubCellInst_LFInst_14_n23 ) );
  NAND2_X1 SubCellInst_LFInst_14_U5  ( .A1(SubCellInst_LFInst_14_n29 ), .A2(
        SubCellInst_LFInst_14_n33 ), .ZN(SubCellInst_LFInst_14_n26 ) );
  INV_X1 SubCellInst_LFInst_14_U4  ( .A(PermutationOutput[56]), .ZN(
        SubCellInst_LFInst_14_n33 ) );
  INV_X1 SubCellInst_LFInst_14_U3  ( .A(PermutationOutput[59]), .ZN(
        SubCellInst_LFInst_14_n29 ) );
  NOR2_X1 SubCellInst_LFInst_15_U21  ( .A1(SubCellInst_LFInst_15_n36 ), .A2(
        SubCellInst_LFInst_15_n35 ), .ZN(Feedback[60]) );
  NOR2_X1 SubCellInst_LFInst_15_U20  ( .A1(PermutationOutput[61]), .A2(
        SubCellInst_LFInst_15_n34 ), .ZN(SubCellInst_LFInst_15_n36 ) );
  NOR2_X1 SubCellInst_LFInst_15_U19  ( .A1(SubCellInst_LFInst_15_n33 ), .A2(
        SubCellInst_LFInst_15_n32 ), .ZN(SubCellInst_LFInst_15_n34 ) );
  NOR2_X1 SubCellInst_LFInst_15_U18  ( .A1(PermutationOutput[62]), .A2(
        PermutationOutput[63]), .ZN(SubCellInst_LFInst_15_n32 ) );
  NAND2_X1 SubCellInst_LFInst_15_U17  ( .A1(SubCellInst_LFInst_15_n31 ), 
        .A2(SubCellInst_LFInst_15_n30 ), .ZN(Feedback[61]) );
  NAND2_X1 SubCellInst_LFInst_15_U16  ( .A1(PermutationOutput[60]), .A2(
        SubCellInst_LFInst_15_n29 ), .ZN(SubCellInst_LFInst_15_n30 ) );
  NAND2_X1 SubCellInst_LFInst_15_U15  ( .A1(PermutationOutput[62]), .A2(
        SubCellInst_LFInst_15_n28 ), .ZN(SubCellInst_LFInst_15_n31 ) );
  NAND2_X1 SubCellInst_LFInst_15_U14  ( .A1(PermutationOutput[63]), .A2(
        SubCellInst_LFInst_15_n33 ), .ZN(SubCellInst_LFInst_15_n28 ) );
  NAND2_X1 SubCellInst_LFInst_15_U13  ( .A1(SubCellInst_LFInst_15_n27 ), 
        .A2(SubCellInst_LFInst_15_n26 ), .ZN(Feedback[62]) );
  NAND2_X1 SubCellInst_LFInst_15_U12  ( .A1(SubCellInst_LFInst_15_n25 ), 
        .A2(PermutationOutput[61]), .ZN(SubCellInst_LFInst_15_n27 ) );
  NAND2_X1 SubCellInst_LFInst_15_U11  ( .A1(SubCellInst_LFInst_15_n24 ), 
        .A2(SubCellInst_LFInst_15_n23 ), .ZN(SubCellInst_LFInst_15_n25 ) );
  NAND2_X1 SubCellInst_LFInst_15_U10  ( .A1(PermutationOutput[60]), .A2(
        PermutationOutput[63]), .ZN(SubCellInst_LFInst_15_n24 ) );
  NAND2_X1 SubCellInst_LFInst_15_U9  ( .A1(SubCellInst_LFInst_15_n26 ), .A2(
        SubCellInst_LFInst_15_n22 ), .ZN(Feedback[63]) );
  OR2_X1 SubCellInst_LFInst_15_U8  ( .A1(PermutationOutput[61]), .A2(
        SubCellInst_LFInst_15_n35 ), .ZN(SubCellInst_LFInst_15_n22 ) );
  NOR2_X1 SubCellInst_LFInst_15_U7  ( .A1(SubCellInst_LFInst_15_n23 ), .A2(
        SubCellInst_LFInst_15_n29 ), .ZN(SubCellInst_LFInst_15_n35 ) );
  INV_X1 SubCellInst_LFInst_15_U6  ( .A(PermutationOutput[62]), .ZN(
        SubCellInst_LFInst_15_n23 ) );
  NAND2_X1 SubCellInst_LFInst_15_U5  ( .A1(SubCellInst_LFInst_15_n29 ), .A2(
        SubCellInst_LFInst_15_n33 ), .ZN(SubCellInst_LFInst_15_n26 ) );
  INV_X1 SubCellInst_LFInst_15_U4  ( .A(PermutationOutput[60]), .ZN(
        SubCellInst_LFInst_15_n33 ) );
  INV_X1 SubCellInst_LFInst_15_U3  ( .A(PermutationOutput[63]), .ZN(
        SubCellInst_LFInst_15_n29 ) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_0_U2  ( .A(MCInst2_XOR_r0_Inst_0_n3 ), .B(
        MCOutput2[0]), .ZN(MCOutput2[48]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_0_U1  ( .A(Feedback[48]), .B(MCOutput2[16]), 
        .ZN(MCInst2_XOR_r0_Inst_0_n3 ) );
  XOR2_X1 MCInst2_XOR_r1_Inst_0_U1  ( .A(Feedback[32]), .B(MCOutput2[0]), .Z(
        MCOutput2[32]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_1_U2  ( .A(MCInst2_XOR_r0_Inst_1_n3 ), .B(
        MCOutput2[1]), .ZN(MCOutput2[49]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_1_U1  ( .A(Feedback[49]), .B(MCOutput2[17]), 
        .ZN(MCInst2_XOR_r0_Inst_1_n3 ) );
  XOR2_X1 MCInst2_XOR_r1_Inst_1_U1  ( .A(Feedback[33]), .B(MCOutput2[1]), .Z(
        MCOutput2[33]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_2_U2  ( .A(MCInst2_XOR_r0_Inst_2_n3 ), .B(
        MCOutput2[2]), .ZN(MCOutput2[50]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_2_U1  ( .A(Feedback[50]), .B(MCOutput2[18]), 
        .ZN(MCInst2_XOR_r0_Inst_2_n3 ) );
  XOR2_X1 MCInst2_XOR_r1_Inst_2_U1  ( .A(Feedback[34]), .B(MCOutput2[2]), .Z(
        MCOutput2[34]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_3_U2  ( .A(MCInst2_XOR_r0_Inst_3_n3 ), .B(
        MCOutput2[3]), .ZN(MCOutput2[51]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_3_U1  ( .A(Feedback[51]), .B(MCOutput2[19]), 
        .ZN(MCInst2_XOR_r0_Inst_3_n3 ) );
  XOR2_X1 MCInst2_XOR_r1_Inst_3_U1  ( .A(Feedback[35]), .B(MCOutput2[3]), .Z(
        MCOutput2[35]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_4_U2  ( .A(MCInst2_XOR_r0_Inst_4_n3 ), .B(
        MCOutput2[4]), .ZN(MCOutput2[52]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_4_U1  ( .A(Feedback[52]), .B(MCOutput2[20]), 
        .ZN(MCInst2_XOR_r0_Inst_4_n3 ) );
  XOR2_X1 MCInst2_XOR_r1_Inst_4_U1  ( .A(Feedback[36]), .B(MCOutput2[4]), .Z(
        MCOutput2[36]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_5_U2  ( .A(MCInst2_XOR_r0_Inst_5_n3 ), .B(
        MCOutput2[5]), .ZN(MCOutput2[53]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_5_U1  ( .A(Feedback[53]), .B(MCOutput2[21]), 
        .ZN(MCInst2_XOR_r0_Inst_5_n3 ) );
  XOR2_X1 MCInst2_XOR_r1_Inst_5_U1  ( .A(Feedback[37]), .B(MCOutput2[5]), .Z(
        MCOutput2[37]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_6_U2  ( .A(MCInst2_XOR_r0_Inst_6_n3 ), .B(
        MCOutput2[6]), .ZN(MCOutput2[54]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_6_U1  ( .A(Feedback[54]), .B(MCOutput2[22]), 
        .ZN(MCInst2_XOR_r0_Inst_6_n3 ) );
  XOR2_X1 MCInst2_XOR_r1_Inst_6_U1  ( .A(Feedback[38]), .B(MCOutput2[6]), .Z(
        MCOutput2[38]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_7_U2  ( .A(MCInst2_XOR_r0_Inst_7_n3 ), .B(
        MCOutput2[7]), .ZN(MCOutput2[55]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_7_U1  ( .A(Feedback[55]), .B(MCOutput2[23]), 
        .ZN(MCInst2_XOR_r0_Inst_7_n3 ) );
  XOR2_X1 MCInst2_XOR_r1_Inst_7_U1  ( .A(Feedback[39]), .B(MCOutput2[7]), .Z(
        MCOutput2[39]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_8_U2  ( .A(MCInst2_XOR_r0_Inst_8_n3 ), .B(
        MCOutput2[8]), .ZN(MCOutput2[56]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_8_U1  ( .A(Feedback[56]), .B(MCOutput2[24]), 
        .ZN(MCInst2_XOR_r0_Inst_8_n3 ) );
  XOR2_X1 MCInst2_XOR_r1_Inst_8_U1  ( .A(Feedback[40]), .B(MCOutput2[8]), .Z(
        MCOutput2[40]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_9_U2  ( .A(MCInst2_XOR_r0_Inst_9_n3 ), .B(
        MCOutput2[9]), .ZN(MCOutput2[57]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_9_U1  ( .A(Feedback[57]), .B(MCOutput2[25]), 
        .ZN(MCInst2_XOR_r0_Inst_9_n3 ) );
  XOR2_X1 MCInst2_XOR_r1_Inst_9_U1  ( .A(Feedback[41]), .B(MCOutput2[9]), .Z(
        MCOutput2[41]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_10_U2  ( .A(MCInst2_XOR_r0_Inst_10_n3 ), .B(
        MCOutput2[10]), .ZN(MCOutput2[58]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_10_U1  ( .A(Feedback[58]), .B(MCOutput2[26]), 
        .ZN(MCInst2_XOR_r0_Inst_10_n3 ) );
  XOR2_X1 MCInst2_XOR_r1_Inst_10_U1  ( .A(Feedback[42]), .B(MCOutput2[10]), 
        .Z(MCOutput2[42]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_11_U2  ( .A(MCInst2_XOR_r0_Inst_11_n3 ), .B(
        MCOutput2[11]), .ZN(MCOutput2[59]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_11_U1  ( .A(Feedback[59]), .B(MCOutput2[27]), 
        .ZN(MCInst2_XOR_r0_Inst_11_n3 ) );
  XOR2_X1 MCInst2_XOR_r1_Inst_11_U1  ( .A(Feedback[43]), .B(MCOutput2[11]), 
        .Z(MCOutput2[43]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_12_U2  ( .A(MCInst2_XOR_r0_Inst_12_n3 ), .B(
        MCOutput2[12]), .ZN(MCOutput2[60]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_12_U1  ( .A(Feedback[60]), .B(MCOutput2[28]), 
        .ZN(MCInst2_XOR_r0_Inst_12_n3 ) );
  XOR2_X1 MCInst2_XOR_r1_Inst_12_U1  ( .A(Feedback[44]), .B(MCOutput2[12]), 
        .Z(MCOutput2[44]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_13_U2  ( .A(MCInst2_XOR_r0_Inst_13_n3 ), .B(
        MCOutput2[13]), .ZN(MCOutput2[61]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_13_U1  ( .A(Feedback[61]), .B(MCOutput2[29]), 
        .ZN(MCInst2_XOR_r0_Inst_13_n3 ) );
  XOR2_X1 MCInst2_XOR_r1_Inst_13_U1  ( .A(Feedback[45]), .B(MCOutput2[13]), 
        .Z(MCOutput2[45]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_14_U2  ( .A(MCInst2_XOR_r0_Inst_14_n3 ), .B(
        MCOutput2[14]), .ZN(MCOutput2[62]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_14_U1  ( .A(Feedback[62]), .B(MCOutput2[30]), 
        .ZN(MCInst2_XOR_r0_Inst_14_n3 ) );
  XOR2_X1 MCInst2_XOR_r1_Inst_14_U1  ( .A(Feedback[46]), .B(MCOutput2[14]), 
        .Z(MCOutput2[46]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_15_U2  ( .A(MCInst2_XOR_r0_Inst_15_n3 ), .B(
        MCOutput2[15]), .ZN(MCOutput2[63]) );
  XNOR2_X1 MCInst2_XOR_r0_Inst_15_U1  ( .A(Feedback[63]), .B(MCOutput2[31]), 
        .ZN(MCInst2_XOR_r0_Inst_15_n3 ) );
  XOR2_X1 MCInst2_XOR_r1_Inst_15_U1  ( .A(Feedback[47]), .B(MCOutput2[15]), 
        .Z(MCOutput2[47]) );
  XOR2_X1 AddKeyXOR12_XORInst_0_0_U1  ( .A(MCOutput2[48]), .B(Key[48]), .Z(
        AddRoundKeyOutput2[48]) );
  XOR2_X1 AddKeyXOR12_XORInst_0_1_U1  ( .A(MCOutput2[49]), .B(Key[49]), .Z(
        AddRoundKeyOutput2[49]) );
  XOR2_X1 AddKeyXOR12_XORInst_0_2_U1  ( .A(MCOutput2[50]), .B(Key[50]), .Z(
        AddRoundKeyOutput2[50]) );
  XOR2_X1 AddKeyXOR12_XORInst_0_3_U1  ( .A(MCOutput2[51]), .B(Key[51]), .Z(
        AddRoundKeyOutput2[51]) );
  XOR2_X1 AddKeyXOR12_XORInst_1_0_U1  ( .A(MCOutput2[52]), .B(Key[52]), .Z(
        AddRoundKeyOutput2[52]) );
  XOR2_X1 AddKeyXOR12_XORInst_1_1_U1  ( .A(MCOutput2[53]), .B(Key[53]), .Z(
        AddRoundKeyOutput2[53]) );
  XOR2_X1 AddKeyXOR12_XORInst_1_2_U1  ( .A(MCOutput2[54]), .B(Key[54]), .Z(
        AddRoundKeyOutput2[54]) );
  XOR2_X1 AddKeyXOR12_XORInst_1_3_U1  ( .A(MCOutput2[55]), .B(Key[55]), .Z(
        AddRoundKeyOutput2[55]) );
  XOR2_X1 AddKeyXOR12_XORInst_2_0_U1  ( .A(MCOutput2[56]), .B(Key[56]), .Z(
        AddRoundKeyOutput2[56]) );
  XOR2_X1 AddKeyXOR12_XORInst_2_1_U1  ( .A(MCOutput2[57]), .B(Key[57]), .Z(
        AddRoundKeyOutput2[57]) );
  XOR2_X1 AddKeyXOR12_XORInst_2_2_U1  ( .A(MCOutput2[58]), .B(Key[58]), .Z(
        AddRoundKeyOutput2[58]) );
  XOR2_X1 AddKeyXOR12_XORInst_2_3_U1  ( .A(MCOutput2[59]), .B(Key[59]), .Z(
        AddRoundKeyOutput2[59]) );
  XOR2_X1 AddKeyXOR12_XORInst_3_0_U1  ( .A(MCOutput2[60]), .B(Key[60]), .Z(
        AddRoundKeyOutput2[60]) );
  XOR2_X1 AddKeyXOR12_XORInst_3_1_U1  ( .A(MCOutput2[61]), .B(Key[61]), .Z(
        AddRoundKeyOutput2[61]) );
  XOR2_X1 AddKeyXOR12_XORInst_3_2_U1  ( .A(MCOutput2[62]), .B(Key[62]), .Z(
        AddRoundKeyOutput2[62]) );
  XOR2_X1 AddKeyXOR12_XORInst_3_3_U1  ( .A(MCOutput2[63]), .B(Key[63]), .Z(
        AddRoundKeyOutput2[63]) );
  XOR2_X1 AddKeyConstXOR2_XORInst_0_0_U1  ( .A(Key[40]), .B(MCOutput2[40]), 
        .Z(AddRoundKeyOutput2[40]) );
  XOR2_X1 AddKeyConstXOR2_XORInst_0_1_U1  ( .A(Key[41]), .B(MCOutput2[41]), 
        .Z(AddRoundKeyOutput2[41]) );
  XOR2_X1 AddKeyConstXOR2_XORInst_0_2_U1  ( .A(Key[42]), .B(MCOutput2[42]), 
        .Z(AddRoundKeyOutput2[42]) );
  XOR2_X1 AddKeyConstXOR2_XORInst_0_3_U1  ( .A(Key[43]), .B(MCOutput2[43]), 
        .Z(AddRoundKeyOutput2[43]) );
  XOR2_X1 AddKeyConstXOR2_XORInst_1_0_U1  ( .A(Key[44]), .B(MCOutput2[44]), 
        .Z(AddRoundKeyOutput2[44]) );
  XOR2_X1 AddKeyConstXOR2_XORInst_1_1_U1  ( .A(Key[45]), .B(MCOutput2[45]), 
        .Z(AddRoundKeyOutput2[45]) );
  XOR2_X1 AddKeyConstXOR2_XORInst_1_2_U1  ( .A(Key[46]), .B(MCOutput2[46]), 
        .Z(AddRoundKeyOutput2[46]) );
  XOR2_X1 AddKeyConstXOR2_XORInst_1_3_U1  ( .A(Key[47]), .B(MCOutput2[47]), 
        .Z(AddRoundKeyOutput2[47]) );
  XOR2_X1 AddKeyXOR22_XORInst_0_0_U1  ( .A(MCOutput2[0]), .B(Key[0]), .Z(
        AddRoundKeyOutput2[0]) );
  XOR2_X1 AddKeyXOR22_XORInst_0_1_U1  ( .A(MCOutput2[1]), .B(Key[1]), .Z(
        AddRoundKeyOutput2[1]) );
  XOR2_X1 AddKeyXOR22_XORInst_0_2_U1  ( .A(MCOutput2[2]), .B(Key[2]), .Z(
        AddRoundKeyOutput2[2]) );
  XOR2_X1 AddKeyXOR22_XORInst_0_3_U1  ( .A(MCOutput2[3]), .B(Key[3]), .Z(
        AddRoundKeyOutput2[3]) );
  XOR2_X1 AddKeyXOR22_XORInst_1_0_U1  ( .A(MCOutput2[4]), .B(Key[4]), .Z(
        AddRoundKeyOutput2[4]) );
  XOR2_X1 AddKeyXOR22_XORInst_1_1_U1  ( .A(MCOutput2[5]), .B(Key[5]), .Z(
        AddRoundKeyOutput2[5]) );
  XOR2_X1 AddKeyXOR22_XORInst_1_2_U1  ( .A(MCOutput2[6]), .B(Key[6]), .Z(
        AddRoundKeyOutput2[6]) );
  XOR2_X1 AddKeyXOR22_XORInst_1_3_U1  ( .A(MCOutput2[7]), .B(Key[7]), .Z(
        AddRoundKeyOutput2[7]) );
  XOR2_X1 AddKeyXOR22_XORInst_2_0_U1  ( .A(MCOutput2[8]), .B(Key[8]), .Z(
        AddRoundKeyOutput2[8]) );
  XOR2_X1 AddKeyXOR22_XORInst_2_1_U1  ( .A(MCOutput2[9]), .B(Key[9]), .Z(
        AddRoundKeyOutput2[9]) );
  XOR2_X1 AddKeyXOR22_XORInst_2_2_U1  ( .A(MCOutput2[10]), .B(Key[10]), .Z(
        AddRoundKeyOutput2[10]) );
  XOR2_X1 AddKeyXOR22_XORInst_2_3_U1  ( .A(MCOutput2[11]), .B(Key[11]), .Z(
        AddRoundKeyOutput2[11]) );
  XOR2_X1 AddKeyXOR22_XORInst_3_0_U1  ( .A(MCOutput2[12]), .B(Key[12]), .Z(
        AddRoundKeyOutput2[12]) );
  XOR2_X1 AddKeyXOR22_XORInst_3_1_U1  ( .A(MCOutput2[13]), .B(Key[13]), .Z(
        AddRoundKeyOutput2[13]) );
  XOR2_X1 AddKeyXOR22_XORInst_3_2_U1  ( .A(MCOutput2[14]), .B(Key[14]), .Z(
        AddRoundKeyOutput2[14]) );
  XOR2_X1 AddKeyXOR22_XORInst_3_3_U1  ( .A(MCOutput2[15]), .B(Key[15]), .Z(
        AddRoundKeyOutput2[15]) );
  XOR2_X1 AddKeyXOR22_XORInst_4_0_U1  ( .A(MCOutput2[16]), .B(Key[16]), .Z(
        AddRoundKeyOutput2[16]) );
  XOR2_X1 AddKeyXOR22_XORInst_4_1_U1  ( .A(MCOutput2[17]), .B(Key[17]), .Z(
        AddRoundKeyOutput2[17]) );
  XOR2_X1 AddKeyXOR22_XORInst_4_2_U1  ( .A(MCOutput2[18]), .B(Key[18]), .Z(
        AddRoundKeyOutput2[18]) );
  XOR2_X1 AddKeyXOR22_XORInst_4_3_U1  ( .A(MCOutput2[19]), .B(Key[19]), .Z(
        AddRoundKeyOutput2[19]) );
  XOR2_X1 AddKeyXOR22_XORInst_5_0_U1  ( .A(MCOutput2[20]), .B(Key[20]), .Z(
        AddRoundKeyOutput2[20]) );
  XOR2_X1 AddKeyXOR22_XORInst_5_1_U1  ( .A(MCOutput2[21]), .B(Key[21]), .Z(
        AddRoundKeyOutput2[21]) );
  XOR2_X1 AddKeyXOR22_XORInst_5_2_U1  ( .A(MCOutput2[22]), .B(Key[22]), .Z(
        AddRoundKeyOutput2[22]) );
  XOR2_X1 AddKeyXOR22_XORInst_5_3_U1  ( .A(MCOutput2[23]), .B(Key[23]), .Z(
        AddRoundKeyOutput2[23]) );
  XOR2_X1 AddKeyXOR22_XORInst_6_0_U1  ( .A(MCOutput2[24]), .B(Key[24]), .Z(
        AddRoundKeyOutput2[24]) );
  XOR2_X1 AddKeyXOR22_XORInst_6_1_U1  ( .A(MCOutput2[25]), .B(Key[25]), .Z(
        AddRoundKeyOutput2[25]) );
  XOR2_X1 AddKeyXOR22_XORInst_6_2_U1  ( .A(MCOutput2[26]), .B(Key[26]), .Z(
        AddRoundKeyOutput2[26]) );
  XOR2_X1 AddKeyXOR22_XORInst_6_3_U1  ( .A(MCOutput2[27]), .B(Key[27]), .Z(
        AddRoundKeyOutput2[27]) );
  XOR2_X1 AddKeyXOR22_XORInst_7_0_U1  ( .A(MCOutput2[28]), .B(Key[28]), .Z(
        AddRoundKeyOutput2[28]) );
  XOR2_X1 AddKeyXOR22_XORInst_7_1_U1  ( .A(MCOutput2[29]), .B(Key[29]), .Z(
        AddRoundKeyOutput2[29]) );
  XOR2_X1 AddKeyXOR22_XORInst_7_2_U1  ( .A(MCOutput2[30]), .B(Key[30]), .Z(
        AddRoundKeyOutput2[30]) );
  XOR2_X1 AddKeyXOR22_XORInst_7_3_U1  ( .A(MCOutput2[31]), .B(Key[31]), .Z(
        AddRoundKeyOutput2[31]) );
  XOR2_X1 AddKeyXOR22_XORInst_8_0_U1  ( .A(MCOutput2[32]), .B(Key[32]), .Z(
        AddRoundKeyOutput2[32]) );
  XOR2_X1 AddKeyXOR22_XORInst_8_1_U1  ( .A(MCOutput2[33]), .B(Key[33]), .Z(
        AddRoundKeyOutput2[33]) );
  XOR2_X1 AddKeyXOR22_XORInst_8_2_U1  ( .A(MCOutput2[34]), .B(Key[34]), .Z(
        AddRoundKeyOutput2[34]) );
  XOR2_X1 AddKeyXOR22_XORInst_8_3_U1  ( .A(MCOutput2[35]), .B(Key[35]), .Z(
        AddRoundKeyOutput2[35]) );
  XOR2_X1 AddKeyXOR22_XORInst_9_0_U1  ( .A(MCOutput2[36]), .B(Key[36]), .Z(
        AddRoundKeyOutput2[36]) );
  XOR2_X1 AddKeyXOR22_XORInst_9_1_U1  ( .A(MCOutput2[37]), .B(Key[37]), .Z(
        AddRoundKeyOutput2[37]) );
  XOR2_X1 AddKeyXOR22_XORInst_9_2_U1  ( .A(MCOutput2[38]), .B(Key[38]), .Z(
        AddRoundKeyOutput2[38]) );
  XOR2_X1 AddKeyXOR22_XORInst_9_3_U1  ( .A(MCOutput2[39]), .B(Key[39]), .Z(
        AddRoundKeyOutput2[39]) );
  DFF_X1 StateReg2_s_current_state_reg[0]  ( .D(AddRoundKeyOutput2[0]), .CK(
        clk), .Q(PermutationOutput2[60]) );
  DFF_X1 StateReg2_s_current_state_reg[1]  ( .D(AddRoundKeyOutput2[1]), .CK(
        clk), .Q(PermutationOutput2[61]) );
  DFF_X1 StateReg2_s_current_state_reg[2]  ( .D(AddRoundKeyOutput2[2]), .CK(
        clk), .Q(PermutationOutput2[62]) );
  DFF_X1 StateReg2_s_current_state_reg[3]  ( .D(AddRoundKeyOutput2[3]), .CK(
        clk), .Q(PermutationOutput2[63]) );
  DFF_X1 StateReg2_s_current_state_reg[4]  ( .D(AddRoundKeyOutput2[4]), .CK(
        clk), .Q(PermutationOutput2[48]) );
  DFF_X1 StateReg2_s_current_state_reg[5]  ( .D(AddRoundKeyOutput2[5]), .CK(
        clk), .Q(PermutationOutput2[49]) );
  DFF_X1 StateReg2_s_current_state_reg[6]  ( .D(AddRoundKeyOutput2[6]), .CK(
        clk), .Q(PermutationOutput2[50]) );
  DFF_X1 StateReg2_s_current_state_reg[7]  ( .D(AddRoundKeyOutput2[7]), .CK(
        clk), .Q(PermutationOutput2[51]) );
  DFF_X1 StateReg2_s_current_state_reg[8]  ( .D(AddRoundKeyOutput2[8]), .CK(
        clk), .Q(PermutationOutput2[52]) );
  DFF_X1 StateReg2_s_current_state_reg[9]  ( .D(AddRoundKeyOutput2[9]), .CK(
        clk), .Q(PermutationOutput2[53]) );
  DFF_X1 StateReg2_s_current_state_reg[10]  ( .D(AddRoundKeyOutput2[10]), 
        .CK(clk), .Q(PermutationOutput2[54]) );
  DFF_X1 StateReg2_s_current_state_reg[11]  ( .D(AddRoundKeyOutput2[11]), 
        .CK(clk), .Q(PermutationOutput2[55]) );
  DFF_X1 StateReg2_s_current_state_reg[12]  ( .D(AddRoundKeyOutput2[12]), 
        .CK(clk), .Q(PermutationOutput2[56]) );
  DFF_X1 StateReg2_s_current_state_reg[13]  ( .D(AddRoundKeyOutput2[13]), 
        .CK(clk), .Q(PermutationOutput2[57]) );
  DFF_X1 StateReg2_s_current_state_reg[14]  ( .D(AddRoundKeyOutput2[14]), 
        .CK(clk), .Q(PermutationOutput2[58]) );
  DFF_X1 StateReg2_s_current_state_reg[15]  ( .D(AddRoundKeyOutput2[15]), 
        .CK(clk), .Q(PermutationOutput2[59]) );
  DFF_X1 StateReg2_s_current_state_reg[16]  ( .D(AddRoundKeyOutput2[16]), 
        .CK(clk), .Q(PermutationOutput2[32]) );
  DFF_X1 StateReg2_s_current_state_reg[17]  ( .D(AddRoundKeyOutput2[17]), 
        .CK(clk), .Q(PermutationOutput2[33]) );
  DFF_X1 StateReg2_s_current_state_reg[18]  ( .D(AddRoundKeyOutput2[18]), 
        .CK(clk), .Q(PermutationOutput2[34]) );
  DFF_X1 StateReg2_s_current_state_reg[19]  ( .D(AddRoundKeyOutput2[19]), 
        .CK(clk), .Q(PermutationOutput2[35]) );
  DFF_X1 StateReg2_s_current_state_reg[20]  ( .D(AddRoundKeyOutput2[20]), 
        .CK(clk), .Q(PermutationOutput2[44]) );
  DFF_X1 StateReg2_s_current_state_reg[21]  ( .D(AddRoundKeyOutput2[21]), 
        .CK(clk), .Q(PermutationOutput2[45]) );
  DFF_X1 StateReg2_s_current_state_reg[22]  ( .D(AddRoundKeyOutput2[22]), 
        .CK(clk), .Q(PermutationOutput2[46]) );
  DFF_X1 StateReg2_s_current_state_reg[23]  ( .D(AddRoundKeyOutput2[23]), 
        .CK(clk), .Q(PermutationOutput2[47]) );
  DFF_X1 StateReg2_s_current_state_reg[24]  ( .D(AddRoundKeyOutput2[24]), 
        .CK(clk), .Q(PermutationOutput2[40]) );
  DFF_X1 StateReg2_s_current_state_reg[25]  ( .D(AddRoundKeyOutput2[25]), 
        .CK(clk), .Q(PermutationOutput2[41]) );
  DFF_X1 StateReg2_s_current_state_reg[26]  ( .D(AddRoundKeyOutput2[26]), 
        .CK(clk), .Q(PermutationOutput2[42]) );
  DFF_X1 StateReg2_s_current_state_reg[27]  ( .D(AddRoundKeyOutput2[27]), 
        .CK(clk), .Q(PermutationOutput2[43]) );
  DFF_X1 StateReg2_s_current_state_reg[28]  ( .D(AddRoundKeyOutput2[28]), 
        .CK(clk), .Q(PermutationOutput2[36]) );
  DFF_X1 StateReg2_s_current_state_reg[29]  ( .D(AddRoundKeyOutput2[29]), 
        .CK(clk), .Q(PermutationOutput2[37]) );
  DFF_X1 StateReg2_s_current_state_reg[30]  ( .D(AddRoundKeyOutput2[30]), 
        .CK(clk), .Q(PermutationOutput2[38]) );
  DFF_X1 StateReg2_s_current_state_reg[31]  ( .D(AddRoundKeyOutput2[31]), 
        .CK(clk), .Q(PermutationOutput2[39]) );
  DFF_X1 StateReg2_s_current_state_reg[32]  ( .D(AddRoundKeyOutput2[32]), 
        .CK(clk), .Q(PermutationOutput2[16]) );
  DFF_X1 StateReg2_s_current_state_reg[33]  ( .D(AddRoundKeyOutput2[33]), 
        .CK(clk), .Q(PermutationOutput2[17]) );
  DFF_X1 StateReg2_s_current_state_reg[34]  ( .D(AddRoundKeyOutput2[34]), 
        .CK(clk), .Q(PermutationOutput2[18]) );
  DFF_X1 StateReg2_s_current_state_reg[35]  ( .D(AddRoundKeyOutput2[35]), 
        .CK(clk), .Q(PermutationOutput2[19]) );
  DFF_X1 StateReg2_s_current_state_reg[36]  ( .D(AddRoundKeyOutput2[36]), 
        .CK(clk), .Q(PermutationOutput2[28]) );
  DFF_X1 StateReg2_s_current_state_reg[37]  ( .D(AddRoundKeyOutput2[37]), 
        .CK(clk), .Q(PermutationOutput2[29]) );
  DFF_X1 StateReg2_s_current_state_reg[38]  ( .D(AddRoundKeyOutput2[38]), 
        .CK(clk), .Q(PermutationOutput2[30]) );
  DFF_X1 StateReg2_s_current_state_reg[39]  ( .D(AddRoundKeyOutput2[39]), 
        .CK(clk), .Q(PermutationOutput2[31]) );
  DFF_X1 StateReg2_s_current_state_reg[40]  ( .D(AddRoundKeyOutput2[40]), 
        .CK(clk), .Q(PermutationOutput2[24]) );
  DFF_X1 StateReg2_s_current_state_reg[41]  ( .D(AddRoundKeyOutput2[41]), 
        .CK(clk), .Q(PermutationOutput2[25]) );
  DFF_X1 StateReg2_s_current_state_reg[42]  ( .D(AddRoundKeyOutput2[42]), 
        .CK(clk), .Q(PermutationOutput2[26]) );
  DFF_X1 StateReg2_s_current_state_reg[43]  ( .D(AddRoundKeyOutput2[43]), 
        .CK(clk), .Q(PermutationOutput2[27]) );
  DFF_X1 StateReg2_s_current_state_reg[44]  ( .D(AddRoundKeyOutput2[44]), 
        .CK(clk), .Q(PermutationOutput2[20]) );
  DFF_X1 StateReg2_s_current_state_reg[45]  ( .D(AddRoundKeyOutput2[45]), 
        .CK(clk), .Q(PermutationOutput2[21]) );
  DFF_X1 StateReg2_s_current_state_reg[46]  ( .D(AddRoundKeyOutput2[46]), 
        .CK(clk), .Q(PermutationOutput2[22]) );
  DFF_X1 StateReg2_s_current_state_reg[47]  ( .D(AddRoundKeyOutput2[47]), 
        .CK(clk), .Q(PermutationOutput2[23]) );
  DFF_X1 StateReg2_s_current_state_reg[48]  ( .D(AddRoundKeyOutput2[48]), 
        .CK(clk), .Q(PermutationOutput2[4]) );
  DFF_X1 StateReg2_s_current_state_reg[49]  ( .D(AddRoundKeyOutput2[49]), 
        .CK(clk), .Q(PermutationOutput2[5]) );
  DFF_X1 StateReg2_s_current_state_reg[50]  ( .D(AddRoundKeyOutput2[50]), 
        .CK(clk), .Q(PermutationOutput2[6]) );
  DFF_X1 StateReg2_s_current_state_reg[51]  ( .D(AddRoundKeyOutput2[51]), 
        .CK(clk), .Q(PermutationOutput2[7]) );
  DFF_X1 StateReg2_s_current_state_reg[52]  ( .D(AddRoundKeyOutput2[52]), 
        .CK(clk), .Q(PermutationOutput2[8]) );
  DFF_X1 StateReg2_s_current_state_reg[53]  ( .D(AddRoundKeyOutput2[53]), 
        .CK(clk), .Q(PermutationOutput2[9]) );
  DFF_X1 StateReg2_s_current_state_reg[54]  ( .D(AddRoundKeyOutput2[54]), 
        .CK(clk), .Q(PermutationOutput2[10]) );
  DFF_X1 StateReg2_s_current_state_reg[55]  ( .D(AddRoundKeyOutput2[55]), 
        .CK(clk), .Q(PermutationOutput2[11]) );
  DFF_X1 StateReg2_s_current_state_reg[56]  ( .D(AddRoundKeyOutput2[56]), 
        .CK(clk), .Q(PermutationOutput2[12]) );
  DFF_X1 StateReg2_s_current_state_reg[57]  ( .D(AddRoundKeyOutput2[57]), 
        .CK(clk), .Q(PermutationOutput2[13]) );
  DFF_X1 StateReg2_s_current_state_reg[58]  ( .D(AddRoundKeyOutput2[58]), 
        .CK(clk), .Q(PermutationOutput2[14]) );
  DFF_X1 StateReg2_s_current_state_reg[59]  ( .D(AddRoundKeyOutput2[59]), 
        .CK(clk), .Q(PermutationOutput2[15]) );
  DFF_X1 StateReg2_s_current_state_reg[60]  ( .D(AddRoundKeyOutput2[60]), 
        .CK(clk), .Q(PermutationOutput2[0]) );
  DFF_X1 StateReg2_s_current_state_reg[61]  ( .D(AddRoundKeyOutput2[61]), 
        .CK(clk), .Q(PermutationOutput2[1]) );
  DFF_X1 StateReg2_s_current_state_reg[62]  ( .D(AddRoundKeyOutput2[62]), 
        .CK(clk), .Q(PermutationOutput2[2]) );
  DFF_X1 StateReg2_s_current_state_reg[63]  ( .D(AddRoundKeyOutput2[63]), 
        .CK(clk), .Q(PermutationOutput2[3]) );
  NOR2_X1 SubCellInst2_LFInst_0_U21  ( .A1(SubCellInst2_LFInst_0_n36 ), .A2(
        SubCellInst2_LFInst_0_n35 ), .ZN(Output[0]) );
  NOR2_X1 SubCellInst2_LFInst_0_U20  ( .A1(PermutationOutput2[1]), .A2(
        SubCellInst2_LFInst_0_n34 ), .ZN(SubCellInst2_LFInst_0_n36 ) );
  NOR2_X1 SubCellInst2_LFInst_0_U19  ( .A1(SubCellInst2_LFInst_0_n33 ), .A2(
        SubCellInst2_LFInst_0_n32 ), .ZN(SubCellInst2_LFInst_0_n34 ) );
  NOR2_X1 SubCellInst2_LFInst_0_U18  ( .A1(PermutationOutput2[2]), .A2(
        PermutationOutput2[3]), .ZN(SubCellInst2_LFInst_0_n32 ) );
  NAND2_X1 SubCellInst2_LFInst_0_U17  ( .A1(SubCellInst2_LFInst_0_n31 ), 
        .A2(SubCellInst2_LFInst_0_n30 ), .ZN(Output[1]) );
  NAND2_X1 SubCellInst2_LFInst_0_U16  ( .A1(PermutationOutput2[0]), .A2(
        SubCellInst2_LFInst_0_n29 ), .ZN(SubCellInst2_LFInst_0_n30 ) );
  NAND2_X1 SubCellInst2_LFInst_0_U15  ( .A1(PermutationOutput2[2]), .A2(
        SubCellInst2_LFInst_0_n28 ), .ZN(SubCellInst2_LFInst_0_n31 ) );
  NAND2_X1 SubCellInst2_LFInst_0_U14  ( .A1(PermutationOutput2[3]), .A2(
        SubCellInst2_LFInst_0_n33 ), .ZN(SubCellInst2_LFInst_0_n28 ) );
  NAND2_X1 SubCellInst2_LFInst_0_U13  ( .A1(SubCellInst2_LFInst_0_n27 ), 
        .A2(SubCellInst2_LFInst_0_n26 ), .ZN(Output[2]) );
  NAND2_X1 SubCellInst2_LFInst_0_U12  ( .A1(SubCellInst2_LFInst_0_n25 ), 
        .A2(PermutationOutput2[1]), .ZN(SubCellInst2_LFInst_0_n27 ) );
  NAND2_X1 SubCellInst2_LFInst_0_U11  ( .A1(SubCellInst2_LFInst_0_n24 ), 
        .A2(SubCellInst2_LFInst_0_n23 ), .ZN(SubCellInst2_LFInst_0_n25 ) );
  NAND2_X1 SubCellInst2_LFInst_0_U10  ( .A1(PermutationOutput2[0]), .A2(
        PermutationOutput2[3]), .ZN(SubCellInst2_LFInst_0_n24 ) );
  NAND2_X1 SubCellInst2_LFInst_0_U9  ( .A1(SubCellInst2_LFInst_0_n26 ), .A2(
        SubCellInst2_LFInst_0_n22 ), .ZN(Output[3]) );
  OR2_X1 SubCellInst2_LFInst_0_U8  ( .A1(PermutationOutput2[1]), .A2(
        SubCellInst2_LFInst_0_n35 ), .ZN(SubCellInst2_LFInst_0_n22 ) );
  NOR2_X1 SubCellInst2_LFInst_0_U7  ( .A1(SubCellInst2_LFInst_0_n23 ), .A2(
        SubCellInst2_LFInst_0_n29 ), .ZN(SubCellInst2_LFInst_0_n35 ) );
  INV_X1 SubCellInst2_LFInst_0_U6  ( .A(PermutationOutput2[2]), .ZN(
        SubCellInst2_LFInst_0_n23 ) );
  NAND2_X1 SubCellInst2_LFInst_0_U5  ( .A1(SubCellInst2_LFInst_0_n29 ), .A2(
        SubCellInst2_LFInst_0_n33 ), .ZN(SubCellInst2_LFInst_0_n26 ) );
  INV_X1 SubCellInst2_LFInst_0_U4  ( .A(PermutationOutput2[0]), .ZN(
        SubCellInst2_LFInst_0_n33 ) );
  INV_X1 SubCellInst2_LFInst_0_U3  ( .A(PermutationOutput2[3]), .ZN(
        SubCellInst2_LFInst_0_n29 ) );
  NOR2_X1 SubCellInst2_LFInst_1_U21  ( .A1(SubCellInst2_LFInst_1_n36 ), .A2(
        SubCellInst2_LFInst_1_n35 ), .ZN(Output[4]) );
  NOR2_X1 SubCellInst2_LFInst_1_U20  ( .A1(PermutationOutput2[5]), .A2(
        SubCellInst2_LFInst_1_n34 ), .ZN(SubCellInst2_LFInst_1_n36 ) );
  NOR2_X1 SubCellInst2_LFInst_1_U19  ( .A1(SubCellInst2_LFInst_1_n33 ), .A2(
        SubCellInst2_LFInst_1_n32 ), .ZN(SubCellInst2_LFInst_1_n34 ) );
  NOR2_X1 SubCellInst2_LFInst_1_U18  ( .A1(PermutationOutput2[6]), .A2(
        PermutationOutput2[7]), .ZN(SubCellInst2_LFInst_1_n32 ) );
  NAND2_X1 SubCellInst2_LFInst_1_U17  ( .A1(SubCellInst2_LFInst_1_n31 ), 
        .A2(SubCellInst2_LFInst_1_n30 ), .ZN(Output[5]) );
  NAND2_X1 SubCellInst2_LFInst_1_U16  ( .A1(PermutationOutput2[4]), .A2(
        SubCellInst2_LFInst_1_n29 ), .ZN(SubCellInst2_LFInst_1_n30 ) );
  NAND2_X1 SubCellInst2_LFInst_1_U15  ( .A1(PermutationOutput2[6]), .A2(
        SubCellInst2_LFInst_1_n28 ), .ZN(SubCellInst2_LFInst_1_n31 ) );
  NAND2_X1 SubCellInst2_LFInst_1_U14  ( .A1(PermutationOutput2[7]), .A2(
        SubCellInst2_LFInst_1_n33 ), .ZN(SubCellInst2_LFInst_1_n28 ) );
  NAND2_X1 SubCellInst2_LFInst_1_U13  ( .A1(SubCellInst2_LFInst_1_n27 ), 
        .A2(SubCellInst2_LFInst_1_n26 ), .ZN(Output[6]) );
  NAND2_X1 SubCellInst2_LFInst_1_U12  ( .A1(SubCellInst2_LFInst_1_n25 ), 
        .A2(PermutationOutput2[5]), .ZN(SubCellInst2_LFInst_1_n27 ) );
  NAND2_X1 SubCellInst2_LFInst_1_U11  ( .A1(SubCellInst2_LFInst_1_n24 ), 
        .A2(SubCellInst2_LFInst_1_n23 ), .ZN(SubCellInst2_LFInst_1_n25 ) );
  NAND2_X1 SubCellInst2_LFInst_1_U10  ( .A1(PermutationOutput2[4]), .A2(
        PermutationOutput2[7]), .ZN(SubCellInst2_LFInst_1_n24 ) );
  NAND2_X1 SubCellInst2_LFInst_1_U9  ( .A1(SubCellInst2_LFInst_1_n26 ), .A2(
        SubCellInst2_LFInst_1_n22 ), .ZN(Output[7]) );
  OR2_X1 SubCellInst2_LFInst_1_U8  ( .A1(PermutationOutput2[5]), .A2(
        SubCellInst2_LFInst_1_n35 ), .ZN(SubCellInst2_LFInst_1_n22 ) );
  NOR2_X1 SubCellInst2_LFInst_1_U7  ( .A1(SubCellInst2_LFInst_1_n23 ), .A2(
        SubCellInst2_LFInst_1_n29 ), .ZN(SubCellInst2_LFInst_1_n35 ) );
  INV_X1 SubCellInst2_LFInst_1_U6  ( .A(PermutationOutput2[6]), .ZN(
        SubCellInst2_LFInst_1_n23 ) );
  NAND2_X1 SubCellInst2_LFInst_1_U5  ( .A1(SubCellInst2_LFInst_1_n29 ), .A2(
        SubCellInst2_LFInst_1_n33 ), .ZN(SubCellInst2_LFInst_1_n26 ) );
  INV_X1 SubCellInst2_LFInst_1_U4  ( .A(PermutationOutput2[4]), .ZN(
        SubCellInst2_LFInst_1_n33 ) );
  INV_X1 SubCellInst2_LFInst_1_U3  ( .A(PermutationOutput2[7]), .ZN(
        SubCellInst2_LFInst_1_n29 ) );
  NOR2_X1 SubCellInst2_LFInst_2_U21  ( .A1(SubCellInst2_LFInst_2_n36 ), .A2(
        SubCellInst2_LFInst_2_n35 ), .ZN(Output[8]) );
  NOR2_X1 SubCellInst2_LFInst_2_U20  ( .A1(PermutationOutput2[9]), .A2(
        SubCellInst2_LFInst_2_n34 ), .ZN(SubCellInst2_LFInst_2_n36 ) );
  NOR2_X1 SubCellInst2_LFInst_2_U19  ( .A1(SubCellInst2_LFInst_2_n33 ), .A2(
        SubCellInst2_LFInst_2_n32 ), .ZN(SubCellInst2_LFInst_2_n34 ) );
  NOR2_X1 SubCellInst2_LFInst_2_U18  ( .A1(PermutationOutput2[10]), .A2(
        PermutationOutput2[11]), .ZN(SubCellInst2_LFInst_2_n32 ) );
  NAND2_X1 SubCellInst2_LFInst_2_U17  ( .A1(SubCellInst2_LFInst_2_n31 ), 
        .A2(SubCellInst2_LFInst_2_n30 ), .ZN(Output[9]) );
  NAND2_X1 SubCellInst2_LFInst_2_U16  ( .A1(PermutationOutput2[8]), .A2(
        SubCellInst2_LFInst_2_n29 ), .ZN(SubCellInst2_LFInst_2_n30 ) );
  NAND2_X1 SubCellInst2_LFInst_2_U15  ( .A1(PermutationOutput2[10]), .A2(
        SubCellInst2_LFInst_2_n28 ), .ZN(SubCellInst2_LFInst_2_n31 ) );
  NAND2_X1 SubCellInst2_LFInst_2_U14  ( .A1(PermutationOutput2[11]), .A2(
        SubCellInst2_LFInst_2_n33 ), .ZN(SubCellInst2_LFInst_2_n28 ) );
  NAND2_X1 SubCellInst2_LFInst_2_U13  ( .A1(SubCellInst2_LFInst_2_n27 ), 
        .A2(SubCellInst2_LFInst_2_n26 ), .ZN(Output[10]) );
  NAND2_X1 SubCellInst2_LFInst_2_U12  ( .A1(SubCellInst2_LFInst_2_n25 ), 
        .A2(PermutationOutput2[9]), .ZN(SubCellInst2_LFInst_2_n27 ) );
  NAND2_X1 SubCellInst2_LFInst_2_U11  ( .A1(SubCellInst2_LFInst_2_n24 ), 
        .A2(SubCellInst2_LFInst_2_n23 ), .ZN(SubCellInst2_LFInst_2_n25 ) );
  NAND2_X1 SubCellInst2_LFInst_2_U10  ( .A1(PermutationOutput2[8]), .A2(
        PermutationOutput2[11]), .ZN(SubCellInst2_LFInst_2_n24 ) );
  NAND2_X1 SubCellInst2_LFInst_2_U9  ( .A1(SubCellInst2_LFInst_2_n26 ), .A2(
        SubCellInst2_LFInst_2_n22 ), .ZN(Output[11]) );
  OR2_X1 SubCellInst2_LFInst_2_U8  ( .A1(PermutationOutput2[9]), .A2(
        SubCellInst2_LFInst_2_n35 ), .ZN(SubCellInst2_LFInst_2_n22 ) );
  NOR2_X1 SubCellInst2_LFInst_2_U7  ( .A1(SubCellInst2_LFInst_2_n23 ), .A2(
        SubCellInst2_LFInst_2_n29 ), .ZN(SubCellInst2_LFInst_2_n35 ) );
  INV_X1 SubCellInst2_LFInst_2_U6  ( .A(PermutationOutput2[10]), .ZN(
        SubCellInst2_LFInst_2_n23 ) );
  NAND2_X1 SubCellInst2_LFInst_2_U5  ( .A1(SubCellInst2_LFInst_2_n29 ), .A2(
        SubCellInst2_LFInst_2_n33 ), .ZN(SubCellInst2_LFInst_2_n26 ) );
  INV_X1 SubCellInst2_LFInst_2_U4  ( .A(PermutationOutput2[8]), .ZN(
        SubCellInst2_LFInst_2_n33 ) );
  INV_X1 SubCellInst2_LFInst_2_U3  ( .A(PermutationOutput2[11]), .ZN(
        SubCellInst2_LFInst_2_n29 ) );
  NOR2_X1 SubCellInst2_LFInst_3_U21  ( .A1(SubCellInst2_LFInst_3_n36 ), .A2(
        SubCellInst2_LFInst_3_n35 ), .ZN(Output[12]) );
  NOR2_X1 SubCellInst2_LFInst_3_U20  ( .A1(PermutationOutput2[13]), .A2(
        SubCellInst2_LFInst_3_n34 ), .ZN(SubCellInst2_LFInst_3_n36 ) );
  NOR2_X1 SubCellInst2_LFInst_3_U19  ( .A1(SubCellInst2_LFInst_3_n33 ), .A2(
        SubCellInst2_LFInst_3_n32 ), .ZN(SubCellInst2_LFInst_3_n34 ) );
  NOR2_X1 SubCellInst2_LFInst_3_U18  ( .A1(PermutationOutput2[14]), .A2(
        PermutationOutput2[15]), .ZN(SubCellInst2_LFInst_3_n32 ) );
  NAND2_X1 SubCellInst2_LFInst_3_U17  ( .A1(SubCellInst2_LFInst_3_n31 ), 
        .A2(SubCellInst2_LFInst_3_n30 ), .ZN(Output[13]) );
  NAND2_X1 SubCellInst2_LFInst_3_U16  ( .A1(PermutationOutput2[12]), .A2(
        SubCellInst2_LFInst_3_n29 ), .ZN(SubCellInst2_LFInst_3_n30 ) );
  NAND2_X1 SubCellInst2_LFInst_3_U15  ( .A1(PermutationOutput2[14]), .A2(
        SubCellInst2_LFInst_3_n28 ), .ZN(SubCellInst2_LFInst_3_n31 ) );
  NAND2_X1 SubCellInst2_LFInst_3_U14  ( .A1(PermutationOutput2[15]), .A2(
        SubCellInst2_LFInst_3_n33 ), .ZN(SubCellInst2_LFInst_3_n28 ) );
  NAND2_X1 SubCellInst2_LFInst_3_U13  ( .A1(SubCellInst2_LFInst_3_n27 ), 
        .A2(SubCellInst2_LFInst_3_n26 ), .ZN(Output[14]) );
  NAND2_X1 SubCellInst2_LFInst_3_U12  ( .A1(SubCellInst2_LFInst_3_n25 ), 
        .A2(PermutationOutput2[13]), .ZN(SubCellInst2_LFInst_3_n27 ) );
  NAND2_X1 SubCellInst2_LFInst_3_U11  ( .A1(SubCellInst2_LFInst_3_n24 ), 
        .A2(SubCellInst2_LFInst_3_n23 ), .ZN(SubCellInst2_LFInst_3_n25 ) );
  NAND2_X1 SubCellInst2_LFInst_3_U10  ( .A1(PermutationOutput2[12]), .A2(
        PermutationOutput2[15]), .ZN(SubCellInst2_LFInst_3_n24 ) );
  NAND2_X1 SubCellInst2_LFInst_3_U9  ( .A1(SubCellInst2_LFInst_3_n26 ), .A2(
        SubCellInst2_LFInst_3_n22 ), .ZN(Output[15]) );
  OR2_X1 SubCellInst2_LFInst_3_U8  ( .A1(PermutationOutput2[13]), .A2(
        SubCellInst2_LFInst_3_n35 ), .ZN(SubCellInst2_LFInst_3_n22 ) );
  NOR2_X1 SubCellInst2_LFInst_3_U7  ( .A1(SubCellInst2_LFInst_3_n23 ), .A2(
        SubCellInst2_LFInst_3_n29 ), .ZN(SubCellInst2_LFInst_3_n35 ) );
  INV_X1 SubCellInst2_LFInst_3_U6  ( .A(PermutationOutput2[14]), .ZN(
        SubCellInst2_LFInst_3_n23 ) );
  NAND2_X1 SubCellInst2_LFInst_3_U5  ( .A1(SubCellInst2_LFInst_3_n29 ), .A2(
        SubCellInst2_LFInst_3_n33 ), .ZN(SubCellInst2_LFInst_3_n26 ) );
  INV_X1 SubCellInst2_LFInst_3_U4  ( .A(PermutationOutput2[12]), .ZN(
        SubCellInst2_LFInst_3_n33 ) );
  INV_X1 SubCellInst2_LFInst_3_U3  ( .A(PermutationOutput2[15]), .ZN(
        SubCellInst2_LFInst_3_n29 ) );
  NOR2_X1 SubCellInst2_LFInst_4_U21  ( .A1(SubCellInst2_LFInst_4_n36 ), .A2(
        SubCellInst2_LFInst_4_n35 ), .ZN(Output[16]) );
  NOR2_X1 SubCellInst2_LFInst_4_U20  ( .A1(PermutationOutput2[17]), .A2(
        SubCellInst2_LFInst_4_n34 ), .ZN(SubCellInst2_LFInst_4_n36 ) );
  NOR2_X1 SubCellInst2_LFInst_4_U19  ( .A1(SubCellInst2_LFInst_4_n33 ), .A2(
        SubCellInst2_LFInst_4_n32 ), .ZN(SubCellInst2_LFInst_4_n34 ) );
  NOR2_X1 SubCellInst2_LFInst_4_U18  ( .A1(PermutationOutput2[18]), .A2(
        PermutationOutput2[19]), .ZN(SubCellInst2_LFInst_4_n32 ) );
  NAND2_X1 SubCellInst2_LFInst_4_U17  ( .A1(SubCellInst2_LFInst_4_n31 ), 
        .A2(SubCellInst2_LFInst_4_n30 ), .ZN(Output[17]) );
  NAND2_X1 SubCellInst2_LFInst_4_U16  ( .A1(PermutationOutput2[16]), .A2(
        SubCellInst2_LFInst_4_n29 ), .ZN(SubCellInst2_LFInst_4_n30 ) );
  NAND2_X1 SubCellInst2_LFInst_4_U15  ( .A1(PermutationOutput2[18]), .A2(
        SubCellInst2_LFInst_4_n28 ), .ZN(SubCellInst2_LFInst_4_n31 ) );
  NAND2_X1 SubCellInst2_LFInst_4_U14  ( .A1(PermutationOutput2[19]), .A2(
        SubCellInst2_LFInst_4_n33 ), .ZN(SubCellInst2_LFInst_4_n28 ) );
  NAND2_X1 SubCellInst2_LFInst_4_U13  ( .A1(SubCellInst2_LFInst_4_n27 ), 
        .A2(SubCellInst2_LFInst_4_n26 ), .ZN(Output[18]) );
  NAND2_X1 SubCellInst2_LFInst_4_U12  ( .A1(SubCellInst2_LFInst_4_n25 ), 
        .A2(PermutationOutput2[17]), .ZN(SubCellInst2_LFInst_4_n27 ) );
  NAND2_X1 SubCellInst2_LFInst_4_U11  ( .A1(SubCellInst2_LFInst_4_n24 ), 
        .A2(SubCellInst2_LFInst_4_n23 ), .ZN(SubCellInst2_LFInst_4_n25 ) );
  NAND2_X1 SubCellInst2_LFInst_4_U10  ( .A1(PermutationOutput2[16]), .A2(
        PermutationOutput2[19]), .ZN(SubCellInst2_LFInst_4_n24 ) );
  NAND2_X1 SubCellInst2_LFInst_4_U9  ( .A1(SubCellInst2_LFInst_4_n26 ), .A2(
        SubCellInst2_LFInst_4_n22 ), .ZN(Output[19]) );
  OR2_X1 SubCellInst2_LFInst_4_U8  ( .A1(PermutationOutput2[17]), .A2(
        SubCellInst2_LFInst_4_n35 ), .ZN(SubCellInst2_LFInst_4_n22 ) );
  NOR2_X1 SubCellInst2_LFInst_4_U7  ( .A1(SubCellInst2_LFInst_4_n23 ), .A2(
        SubCellInst2_LFInst_4_n29 ), .ZN(SubCellInst2_LFInst_4_n35 ) );
  INV_X1 SubCellInst2_LFInst_4_U6  ( .A(PermutationOutput2[18]), .ZN(
        SubCellInst2_LFInst_4_n23 ) );
  NAND2_X1 SubCellInst2_LFInst_4_U5  ( .A1(SubCellInst2_LFInst_4_n29 ), .A2(
        SubCellInst2_LFInst_4_n33 ), .ZN(SubCellInst2_LFInst_4_n26 ) );
  INV_X1 SubCellInst2_LFInst_4_U4  ( .A(PermutationOutput2[16]), .ZN(
        SubCellInst2_LFInst_4_n33 ) );
  INV_X1 SubCellInst2_LFInst_4_U3  ( .A(PermutationOutput2[19]), .ZN(
        SubCellInst2_LFInst_4_n29 ) );
  NOR2_X1 SubCellInst2_LFInst_5_U21  ( .A1(SubCellInst2_LFInst_5_n36 ), .A2(
        SubCellInst2_LFInst_5_n35 ), .ZN(Output[20]) );
  NOR2_X1 SubCellInst2_LFInst_5_U20  ( .A1(PermutationOutput2[21]), .A2(
        SubCellInst2_LFInst_5_n34 ), .ZN(SubCellInst2_LFInst_5_n36 ) );
  NOR2_X1 SubCellInst2_LFInst_5_U19  ( .A1(SubCellInst2_LFInst_5_n33 ), .A2(
        SubCellInst2_LFInst_5_n32 ), .ZN(SubCellInst2_LFInst_5_n34 ) );
  NOR2_X1 SubCellInst2_LFInst_5_U18  ( .A1(PermutationOutput2[22]), .A2(
        PermutationOutput2[23]), .ZN(SubCellInst2_LFInst_5_n32 ) );
  NAND2_X1 SubCellInst2_LFInst_5_U17  ( .A1(SubCellInst2_LFInst_5_n31 ), 
        .A2(SubCellInst2_LFInst_5_n30 ), .ZN(Output[21]) );
  NAND2_X1 SubCellInst2_LFInst_5_U16  ( .A1(PermutationOutput2[20]), .A2(
        SubCellInst2_LFInst_5_n29 ), .ZN(SubCellInst2_LFInst_5_n30 ) );
  NAND2_X1 SubCellInst2_LFInst_5_U15  ( .A1(PermutationOutput2[22]), .A2(
        SubCellInst2_LFInst_5_n28 ), .ZN(SubCellInst2_LFInst_5_n31 ) );
  NAND2_X1 SubCellInst2_LFInst_5_U14  ( .A1(PermutationOutput2[23]), .A2(
        SubCellInst2_LFInst_5_n33 ), .ZN(SubCellInst2_LFInst_5_n28 ) );
  NAND2_X1 SubCellInst2_LFInst_5_U13  ( .A1(SubCellInst2_LFInst_5_n27 ), 
        .A2(SubCellInst2_LFInst_5_n26 ), .ZN(Output[22]) );
  NAND2_X1 SubCellInst2_LFInst_5_U12  ( .A1(SubCellInst2_LFInst_5_n25 ), 
        .A2(PermutationOutput2[21]), .ZN(SubCellInst2_LFInst_5_n27 ) );
  NAND2_X1 SubCellInst2_LFInst_5_U11  ( .A1(SubCellInst2_LFInst_5_n24 ), 
        .A2(SubCellInst2_LFInst_5_n23 ), .ZN(SubCellInst2_LFInst_5_n25 ) );
  NAND2_X1 SubCellInst2_LFInst_5_U10  ( .A1(PermutationOutput2[20]), .A2(
        PermutationOutput2[23]), .ZN(SubCellInst2_LFInst_5_n24 ) );
  NAND2_X1 SubCellInst2_LFInst_5_U9  ( .A1(SubCellInst2_LFInst_5_n26 ), .A2(
        SubCellInst2_LFInst_5_n22 ), .ZN(Output[23]) );
  OR2_X1 SubCellInst2_LFInst_5_U8  ( .A1(PermutationOutput2[21]), .A2(
        SubCellInst2_LFInst_5_n35 ), .ZN(SubCellInst2_LFInst_5_n22 ) );
  NOR2_X1 SubCellInst2_LFInst_5_U7  ( .A1(SubCellInst2_LFInst_5_n23 ), .A2(
        SubCellInst2_LFInst_5_n29 ), .ZN(SubCellInst2_LFInst_5_n35 ) );
  INV_X1 SubCellInst2_LFInst_5_U6  ( .A(PermutationOutput2[22]), .ZN(
        SubCellInst2_LFInst_5_n23 ) );
  NAND2_X1 SubCellInst2_LFInst_5_U5  ( .A1(SubCellInst2_LFInst_5_n29 ), .A2(
        SubCellInst2_LFInst_5_n33 ), .ZN(SubCellInst2_LFInst_5_n26 ) );
  INV_X1 SubCellInst2_LFInst_5_U4  ( .A(PermutationOutput2[20]), .ZN(
        SubCellInst2_LFInst_5_n33 ) );
  INV_X1 SubCellInst2_LFInst_5_U3  ( .A(PermutationOutput2[23]), .ZN(
        SubCellInst2_LFInst_5_n29 ) );
  NOR2_X1 SubCellInst2_LFInst_6_U21  ( .A1(SubCellInst2_LFInst_6_n36 ), .A2(
        SubCellInst2_LFInst_6_n35 ), .ZN(Output[24]) );
  NOR2_X1 SubCellInst2_LFInst_6_U20  ( .A1(PermutationOutput2[25]), .A2(
        SubCellInst2_LFInst_6_n34 ), .ZN(SubCellInst2_LFInst_6_n36 ) );
  NOR2_X1 SubCellInst2_LFInst_6_U19  ( .A1(SubCellInst2_LFInst_6_n33 ), .A2(
        SubCellInst2_LFInst_6_n32 ), .ZN(SubCellInst2_LFInst_6_n34 ) );
  NOR2_X1 SubCellInst2_LFInst_6_U18  ( .A1(PermutationOutput2[26]), .A2(
        PermutationOutput2[27]), .ZN(SubCellInst2_LFInst_6_n32 ) );
  NAND2_X1 SubCellInst2_LFInst_6_U17  ( .A1(SubCellInst2_LFInst_6_n31 ), 
        .A2(SubCellInst2_LFInst_6_n30 ), .ZN(Output[25]) );
  NAND2_X1 SubCellInst2_LFInst_6_U16  ( .A1(PermutationOutput2[24]), .A2(
        SubCellInst2_LFInst_6_n29 ), .ZN(SubCellInst2_LFInst_6_n30 ) );
  NAND2_X1 SubCellInst2_LFInst_6_U15  ( .A1(PermutationOutput2[26]), .A2(
        SubCellInst2_LFInst_6_n28 ), .ZN(SubCellInst2_LFInst_6_n31 ) );
  NAND2_X1 SubCellInst2_LFInst_6_U14  ( .A1(PermutationOutput2[27]), .A2(
        SubCellInst2_LFInst_6_n33 ), .ZN(SubCellInst2_LFInst_6_n28 ) );
  NAND2_X1 SubCellInst2_LFInst_6_U13  ( .A1(SubCellInst2_LFInst_6_n27 ), 
        .A2(SubCellInst2_LFInst_6_n26 ), .ZN(Output[26]) );
  NAND2_X1 SubCellInst2_LFInst_6_U12  ( .A1(SubCellInst2_LFInst_6_n25 ), 
        .A2(PermutationOutput2[25]), .ZN(SubCellInst2_LFInst_6_n27 ) );
  NAND2_X1 SubCellInst2_LFInst_6_U11  ( .A1(SubCellInst2_LFInst_6_n24 ), 
        .A2(SubCellInst2_LFInst_6_n23 ), .ZN(SubCellInst2_LFInst_6_n25 ) );
  NAND2_X1 SubCellInst2_LFInst_6_U10  ( .A1(PermutationOutput2[24]), .A2(
        PermutationOutput2[27]), .ZN(SubCellInst2_LFInst_6_n24 ) );
  NAND2_X1 SubCellInst2_LFInst_6_U9  ( .A1(SubCellInst2_LFInst_6_n26 ), .A2(
        SubCellInst2_LFInst_6_n22 ), .ZN(Output[27]) );
  OR2_X1 SubCellInst2_LFInst_6_U8  ( .A1(PermutationOutput2[25]), .A2(
        SubCellInst2_LFInst_6_n35 ), .ZN(SubCellInst2_LFInst_6_n22 ) );
  NOR2_X1 SubCellInst2_LFInst_6_U7  ( .A1(SubCellInst2_LFInst_6_n23 ), .A2(
        SubCellInst2_LFInst_6_n29 ), .ZN(SubCellInst2_LFInst_6_n35 ) );
  INV_X1 SubCellInst2_LFInst_6_U6  ( .A(PermutationOutput2[26]), .ZN(
        SubCellInst2_LFInst_6_n23 ) );
  NAND2_X1 SubCellInst2_LFInst_6_U5  ( .A1(SubCellInst2_LFInst_6_n29 ), .A2(
        SubCellInst2_LFInst_6_n33 ), .ZN(SubCellInst2_LFInst_6_n26 ) );
  INV_X1 SubCellInst2_LFInst_6_U4  ( .A(PermutationOutput2[24]), .ZN(
        SubCellInst2_LFInst_6_n33 ) );
  INV_X1 SubCellInst2_LFInst_6_U3  ( .A(PermutationOutput2[27]), .ZN(
        SubCellInst2_LFInst_6_n29 ) );
  NOR2_X1 SubCellInst2_LFInst_7_U21  ( .A1(SubCellInst2_LFInst_7_n36 ), .A2(
        SubCellInst2_LFInst_7_n35 ), .ZN(Output[28]) );
  NOR2_X1 SubCellInst2_LFInst_7_U20  ( .A1(PermutationOutput2[29]), .A2(
        SubCellInst2_LFInst_7_n34 ), .ZN(SubCellInst2_LFInst_7_n36 ) );
  NOR2_X1 SubCellInst2_LFInst_7_U19  ( .A1(SubCellInst2_LFInst_7_n33 ), .A2(
        SubCellInst2_LFInst_7_n32 ), .ZN(SubCellInst2_LFInst_7_n34 ) );
  NOR2_X1 SubCellInst2_LFInst_7_U18  ( .A1(PermutationOutput2[30]), .A2(
        PermutationOutput2[31]), .ZN(SubCellInst2_LFInst_7_n32 ) );
  NAND2_X1 SubCellInst2_LFInst_7_U17  ( .A1(SubCellInst2_LFInst_7_n31 ), 
        .A2(SubCellInst2_LFInst_7_n30 ), .ZN(Output[29]) );
  NAND2_X1 SubCellInst2_LFInst_7_U16  ( .A1(PermutationOutput2[28]), .A2(
        SubCellInst2_LFInst_7_n29 ), .ZN(SubCellInst2_LFInst_7_n30 ) );
  NAND2_X1 SubCellInst2_LFInst_7_U15  ( .A1(PermutationOutput2[30]), .A2(
        SubCellInst2_LFInst_7_n28 ), .ZN(SubCellInst2_LFInst_7_n31 ) );
  NAND2_X1 SubCellInst2_LFInst_7_U14  ( .A1(PermutationOutput2[31]), .A2(
        SubCellInst2_LFInst_7_n33 ), .ZN(SubCellInst2_LFInst_7_n28 ) );
  NAND2_X1 SubCellInst2_LFInst_7_U13  ( .A1(SubCellInst2_LFInst_7_n27 ), 
        .A2(SubCellInst2_LFInst_7_n26 ), .ZN(Output[30]) );
  NAND2_X1 SubCellInst2_LFInst_7_U12  ( .A1(SubCellInst2_LFInst_7_n25 ), 
        .A2(PermutationOutput2[29]), .ZN(SubCellInst2_LFInst_7_n27 ) );
  NAND2_X1 SubCellInst2_LFInst_7_U11  ( .A1(SubCellInst2_LFInst_7_n24 ), 
        .A2(SubCellInst2_LFInst_7_n23 ), .ZN(SubCellInst2_LFInst_7_n25 ) );
  NAND2_X1 SubCellInst2_LFInst_7_U10  ( .A1(PermutationOutput2[28]), .A2(
        PermutationOutput2[31]), .ZN(SubCellInst2_LFInst_7_n24 ) );
  NAND2_X1 SubCellInst2_LFInst_7_U9  ( .A1(SubCellInst2_LFInst_7_n26 ), .A2(
        SubCellInst2_LFInst_7_n22 ), .ZN(Output[31]) );
  OR2_X1 SubCellInst2_LFInst_7_U8  ( .A1(PermutationOutput2[29]), .A2(
        SubCellInst2_LFInst_7_n35 ), .ZN(SubCellInst2_LFInst_7_n22 ) );
  NOR2_X1 SubCellInst2_LFInst_7_U7  ( .A1(SubCellInst2_LFInst_7_n23 ), .A2(
        SubCellInst2_LFInst_7_n29 ), .ZN(SubCellInst2_LFInst_7_n35 ) );
  INV_X1 SubCellInst2_LFInst_7_U6  ( .A(PermutationOutput2[30]), .ZN(
        SubCellInst2_LFInst_7_n23 ) );
  NAND2_X1 SubCellInst2_LFInst_7_U5  ( .A1(SubCellInst2_LFInst_7_n29 ), .A2(
        SubCellInst2_LFInst_7_n33 ), .ZN(SubCellInst2_LFInst_7_n26 ) );
  INV_X1 SubCellInst2_LFInst_7_U4  ( .A(PermutationOutput2[28]), .ZN(
        SubCellInst2_LFInst_7_n33 ) );
  INV_X1 SubCellInst2_LFInst_7_U3  ( .A(PermutationOutput2[31]), .ZN(
        SubCellInst2_LFInst_7_n29 ) );
  NOR2_X1 SubCellInst2_LFInst_8_U21  ( .A1(SubCellInst2_LFInst_8_n36 ), .A2(
        SubCellInst2_LFInst_8_n35 ), .ZN(Output[32]) );
  NOR2_X1 SubCellInst2_LFInst_8_U20  ( .A1(PermutationOutput2[33]), .A2(
        SubCellInst2_LFInst_8_n34 ), .ZN(SubCellInst2_LFInst_8_n36 ) );
  NOR2_X1 SubCellInst2_LFInst_8_U19  ( .A1(SubCellInst2_LFInst_8_n33 ), .A2(
        SubCellInst2_LFInst_8_n32 ), .ZN(SubCellInst2_LFInst_8_n34 ) );
  NOR2_X1 SubCellInst2_LFInst_8_U18  ( .A1(PermutationOutput2[34]), .A2(
        PermutationOutput2[35]), .ZN(SubCellInst2_LFInst_8_n32 ) );
  NAND2_X1 SubCellInst2_LFInst_8_U17  ( .A1(SubCellInst2_LFInst_8_n31 ), 
        .A2(SubCellInst2_LFInst_8_n30 ), .ZN(Output[33]) );
  NAND2_X1 SubCellInst2_LFInst_8_U16  ( .A1(PermutationOutput2[32]), .A2(
        SubCellInst2_LFInst_8_n29 ), .ZN(SubCellInst2_LFInst_8_n30 ) );
  NAND2_X1 SubCellInst2_LFInst_8_U15  ( .A1(PermutationOutput2[34]), .A2(
        SubCellInst2_LFInst_8_n28 ), .ZN(SubCellInst2_LFInst_8_n31 ) );
  NAND2_X1 SubCellInst2_LFInst_8_U14  ( .A1(PermutationOutput2[35]), .A2(
        SubCellInst2_LFInst_8_n33 ), .ZN(SubCellInst2_LFInst_8_n28 ) );
  NAND2_X1 SubCellInst2_LFInst_8_U13  ( .A1(SubCellInst2_LFInst_8_n27 ), 
        .A2(SubCellInst2_LFInst_8_n26 ), .ZN(Output[34]) );
  NAND2_X1 SubCellInst2_LFInst_8_U12  ( .A1(SubCellInst2_LFInst_8_n25 ), 
        .A2(PermutationOutput2[33]), .ZN(SubCellInst2_LFInst_8_n27 ) );
  NAND2_X1 SubCellInst2_LFInst_8_U11  ( .A1(SubCellInst2_LFInst_8_n24 ), 
        .A2(SubCellInst2_LFInst_8_n23 ), .ZN(SubCellInst2_LFInst_8_n25 ) );
  NAND2_X1 SubCellInst2_LFInst_8_U10  ( .A1(PermutationOutput2[32]), .A2(
        PermutationOutput2[35]), .ZN(SubCellInst2_LFInst_8_n24 ) );
  NAND2_X1 SubCellInst2_LFInst_8_U9  ( .A1(SubCellInst2_LFInst_8_n26 ), .A2(
        SubCellInst2_LFInst_8_n22 ), .ZN(Output[35]) );
  OR2_X1 SubCellInst2_LFInst_8_U8  ( .A1(PermutationOutput2[33]), .A2(
        SubCellInst2_LFInst_8_n35 ), .ZN(SubCellInst2_LFInst_8_n22 ) );
  NOR2_X1 SubCellInst2_LFInst_8_U7  ( .A1(SubCellInst2_LFInst_8_n23 ), .A2(
        SubCellInst2_LFInst_8_n29 ), .ZN(SubCellInst2_LFInst_8_n35 ) );
  INV_X1 SubCellInst2_LFInst_8_U6  ( .A(PermutationOutput2[34]), .ZN(
        SubCellInst2_LFInst_8_n23 ) );
  NAND2_X1 SubCellInst2_LFInst_8_U5  ( .A1(SubCellInst2_LFInst_8_n29 ), .A2(
        SubCellInst2_LFInst_8_n33 ), .ZN(SubCellInst2_LFInst_8_n26 ) );
  INV_X1 SubCellInst2_LFInst_8_U4  ( .A(PermutationOutput2[32]), .ZN(
        SubCellInst2_LFInst_8_n33 ) );
  INV_X1 SubCellInst2_LFInst_8_U3  ( .A(PermutationOutput2[35]), .ZN(
        SubCellInst2_LFInst_8_n29 ) );
  NOR2_X1 SubCellInst2_LFInst_9_U21  ( .A1(SubCellInst2_LFInst_9_n36 ), .A2(
        SubCellInst2_LFInst_9_n35 ), .ZN(Output[36]) );
  NOR2_X1 SubCellInst2_LFInst_9_U20  ( .A1(PermutationOutput2[37]), .A2(
        SubCellInst2_LFInst_9_n34 ), .ZN(SubCellInst2_LFInst_9_n36 ) );
  NOR2_X1 SubCellInst2_LFInst_9_U19  ( .A1(SubCellInst2_LFInst_9_n33 ), .A2(
        SubCellInst2_LFInst_9_n32 ), .ZN(SubCellInst2_LFInst_9_n34 ) );
  NOR2_X1 SubCellInst2_LFInst_9_U18  ( .A1(PermutationOutput2[38]), .A2(
        PermutationOutput2[39]), .ZN(SubCellInst2_LFInst_9_n32 ) );
  NAND2_X1 SubCellInst2_LFInst_9_U17  ( .A1(SubCellInst2_LFInst_9_n31 ), 
        .A2(SubCellInst2_LFInst_9_n30 ), .ZN(Output[37]) );
  NAND2_X1 SubCellInst2_LFInst_9_U16  ( .A1(PermutationOutput2[36]), .A2(
        SubCellInst2_LFInst_9_n29 ), .ZN(SubCellInst2_LFInst_9_n30 ) );
  NAND2_X1 SubCellInst2_LFInst_9_U15  ( .A1(PermutationOutput2[38]), .A2(
        SubCellInst2_LFInst_9_n28 ), .ZN(SubCellInst2_LFInst_9_n31 ) );
  NAND2_X1 SubCellInst2_LFInst_9_U14  ( .A1(PermutationOutput2[39]), .A2(
        SubCellInst2_LFInst_9_n33 ), .ZN(SubCellInst2_LFInst_9_n28 ) );
  NAND2_X1 SubCellInst2_LFInst_9_U13  ( .A1(SubCellInst2_LFInst_9_n27 ), 
        .A2(SubCellInst2_LFInst_9_n26 ), .ZN(Output[38]) );
  NAND2_X1 SubCellInst2_LFInst_9_U12  ( .A1(SubCellInst2_LFInst_9_n25 ), 
        .A2(PermutationOutput2[37]), .ZN(SubCellInst2_LFInst_9_n27 ) );
  NAND2_X1 SubCellInst2_LFInst_9_U11  ( .A1(SubCellInst2_LFInst_9_n24 ), 
        .A2(SubCellInst2_LFInst_9_n23 ), .ZN(SubCellInst2_LFInst_9_n25 ) );
  NAND2_X1 SubCellInst2_LFInst_9_U10  ( .A1(PermutationOutput2[36]), .A2(
        PermutationOutput2[39]), .ZN(SubCellInst2_LFInst_9_n24 ) );
  NAND2_X1 SubCellInst2_LFInst_9_U9  ( .A1(SubCellInst2_LFInst_9_n26 ), .A2(
        SubCellInst2_LFInst_9_n22 ), .ZN(Output[39]) );
  OR2_X1 SubCellInst2_LFInst_9_U8  ( .A1(PermutationOutput2[37]), .A2(
        SubCellInst2_LFInst_9_n35 ), .ZN(SubCellInst2_LFInst_9_n22 ) );
  NOR2_X1 SubCellInst2_LFInst_9_U7  ( .A1(SubCellInst2_LFInst_9_n23 ), .A2(
        SubCellInst2_LFInst_9_n29 ), .ZN(SubCellInst2_LFInst_9_n35 ) );
  INV_X1 SubCellInst2_LFInst_9_U6  ( .A(PermutationOutput2[38]), .ZN(
        SubCellInst2_LFInst_9_n23 ) );
  NAND2_X1 SubCellInst2_LFInst_9_U5  ( .A1(SubCellInst2_LFInst_9_n29 ), .A2(
        SubCellInst2_LFInst_9_n33 ), .ZN(SubCellInst2_LFInst_9_n26 ) );
  INV_X1 SubCellInst2_LFInst_9_U4  ( .A(PermutationOutput2[36]), .ZN(
        SubCellInst2_LFInst_9_n33 ) );
  INV_X1 SubCellInst2_LFInst_9_U3  ( .A(PermutationOutput2[39]), .ZN(
        SubCellInst2_LFInst_9_n29 ) );
  NOR2_X1 SubCellInst2_LFInst_10_U21  ( .A1(SubCellInst2_LFInst_10_n36 ), 
        .A2(SubCellInst2_LFInst_10_n35 ), .ZN(Output[40]) );
  NOR2_X1 SubCellInst2_LFInst_10_U20  ( .A1(PermutationOutput2[41]), .A2(
        SubCellInst2_LFInst_10_n34 ), .ZN(SubCellInst2_LFInst_10_n36 ) );
  NOR2_X1 SubCellInst2_LFInst_10_U19  ( .A1(SubCellInst2_LFInst_10_n33 ), 
        .A2(SubCellInst2_LFInst_10_n32 ), .ZN(SubCellInst2_LFInst_10_n34 )
         );
  NOR2_X1 SubCellInst2_LFInst_10_U18  ( .A1(PermutationOutput2[42]), .A2(
        PermutationOutput2[43]), .ZN(SubCellInst2_LFInst_10_n32 ) );
  NAND2_X1 SubCellInst2_LFInst_10_U17  ( .A1(SubCellInst2_LFInst_10_n31 ), 
        .A2(SubCellInst2_LFInst_10_n30 ), .ZN(Output[41]) );
  NAND2_X1 SubCellInst2_LFInst_10_U16  ( .A1(PermutationOutput2[40]), .A2(
        SubCellInst2_LFInst_10_n29 ), .ZN(SubCellInst2_LFInst_10_n30 ) );
  NAND2_X1 SubCellInst2_LFInst_10_U15  ( .A1(PermutationOutput2[42]), .A2(
        SubCellInst2_LFInst_10_n28 ), .ZN(SubCellInst2_LFInst_10_n31 ) );
  NAND2_X1 SubCellInst2_LFInst_10_U14  ( .A1(PermutationOutput2[43]), .A2(
        SubCellInst2_LFInst_10_n33 ), .ZN(SubCellInst2_LFInst_10_n28 ) );
  NAND2_X1 SubCellInst2_LFInst_10_U13  ( .A1(SubCellInst2_LFInst_10_n27 ), 
        .A2(SubCellInst2_LFInst_10_n26 ), .ZN(Output[42]) );
  NAND2_X1 SubCellInst2_LFInst_10_U12  ( .A1(SubCellInst2_LFInst_10_n25 ), 
        .A2(PermutationOutput2[41]), .ZN(SubCellInst2_LFInst_10_n27 ) );
  NAND2_X1 SubCellInst2_LFInst_10_U11  ( .A1(SubCellInst2_LFInst_10_n24 ), 
        .A2(SubCellInst2_LFInst_10_n23 ), .ZN(SubCellInst2_LFInst_10_n25 )
         );
  NAND2_X1 SubCellInst2_LFInst_10_U10  ( .A1(PermutationOutput2[40]), .A2(
        PermutationOutput2[43]), .ZN(SubCellInst2_LFInst_10_n24 ) );
  NAND2_X1 SubCellInst2_LFInst_10_U9  ( .A1(SubCellInst2_LFInst_10_n26 ), 
        .A2(SubCellInst2_LFInst_10_n22 ), .ZN(Output[43]) );
  OR2_X1 SubCellInst2_LFInst_10_U8  ( .A1(PermutationOutput2[41]), .A2(
        SubCellInst2_LFInst_10_n35 ), .ZN(SubCellInst2_LFInst_10_n22 ) );
  NOR2_X1 SubCellInst2_LFInst_10_U7  ( .A1(SubCellInst2_LFInst_10_n23 ), 
        .A2(SubCellInst2_LFInst_10_n29 ), .ZN(SubCellInst2_LFInst_10_n35 )
         );
  INV_X1 SubCellInst2_LFInst_10_U6  ( .A(PermutationOutput2[42]), .ZN(
        SubCellInst2_LFInst_10_n23 ) );
  NAND2_X1 SubCellInst2_LFInst_10_U5  ( .A1(SubCellInst2_LFInst_10_n29 ), 
        .A2(SubCellInst2_LFInst_10_n33 ), .ZN(SubCellInst2_LFInst_10_n26 )
         );
  INV_X1 SubCellInst2_LFInst_10_U4  ( .A(PermutationOutput2[40]), .ZN(
        SubCellInst2_LFInst_10_n33 ) );
  INV_X1 SubCellInst2_LFInst_10_U3  ( .A(PermutationOutput2[43]), .ZN(
        SubCellInst2_LFInst_10_n29 ) );
  NOR2_X1 SubCellInst2_LFInst_11_U21  ( .A1(SubCellInst2_LFInst_11_n36 ), 
        .A2(SubCellInst2_LFInst_11_n35 ), .ZN(Output[44]) );
  NOR2_X1 SubCellInst2_LFInst_11_U20  ( .A1(PermutationOutput2[45]), .A2(
        SubCellInst2_LFInst_11_n34 ), .ZN(SubCellInst2_LFInst_11_n36 ) );
  NOR2_X1 SubCellInst2_LFInst_11_U19  ( .A1(SubCellInst2_LFInst_11_n33 ), 
        .A2(SubCellInst2_LFInst_11_n32 ), .ZN(SubCellInst2_LFInst_11_n34 )
         );
  NOR2_X1 SubCellInst2_LFInst_11_U18  ( .A1(PermutationOutput2[46]), .A2(
        PermutationOutput2[47]), .ZN(SubCellInst2_LFInst_11_n32 ) );
  NAND2_X1 SubCellInst2_LFInst_11_U17  ( .A1(SubCellInst2_LFInst_11_n31 ), 
        .A2(SubCellInst2_LFInst_11_n30 ), .ZN(Output[45]) );
  NAND2_X1 SubCellInst2_LFInst_11_U16  ( .A1(PermutationOutput2[44]), .A2(
        SubCellInst2_LFInst_11_n29 ), .ZN(SubCellInst2_LFInst_11_n30 ) );
  NAND2_X1 SubCellInst2_LFInst_11_U15  ( .A1(PermutationOutput2[46]), .A2(
        SubCellInst2_LFInst_11_n28 ), .ZN(SubCellInst2_LFInst_11_n31 ) );
  NAND2_X1 SubCellInst2_LFInst_11_U14  ( .A1(PermutationOutput2[47]), .A2(
        SubCellInst2_LFInst_11_n33 ), .ZN(SubCellInst2_LFInst_11_n28 ) );
  NAND2_X1 SubCellInst2_LFInst_11_U13  ( .A1(SubCellInst2_LFInst_11_n27 ), 
        .A2(SubCellInst2_LFInst_11_n26 ), .ZN(Output[46]) );
  NAND2_X1 SubCellInst2_LFInst_11_U12  ( .A1(SubCellInst2_LFInst_11_n25 ), 
        .A2(PermutationOutput2[45]), .ZN(SubCellInst2_LFInst_11_n27 ) );
  NAND2_X1 SubCellInst2_LFInst_11_U11  ( .A1(SubCellInst2_LFInst_11_n24 ), 
        .A2(SubCellInst2_LFInst_11_n23 ), .ZN(SubCellInst2_LFInst_11_n25 )
         );
  NAND2_X1 SubCellInst2_LFInst_11_U10  ( .A1(PermutationOutput2[44]), .A2(
        PermutationOutput2[47]), .ZN(SubCellInst2_LFInst_11_n24 ) );
  NAND2_X1 SubCellInst2_LFInst_11_U9  ( .A1(SubCellInst2_LFInst_11_n26 ), 
        .A2(SubCellInst2_LFInst_11_n22 ), .ZN(Output[47]) );
  OR2_X1 SubCellInst2_LFInst_11_U8  ( .A1(PermutationOutput2[45]), .A2(
        SubCellInst2_LFInst_11_n35 ), .ZN(SubCellInst2_LFInst_11_n22 ) );
  NOR2_X1 SubCellInst2_LFInst_11_U7  ( .A1(SubCellInst2_LFInst_11_n23 ), 
        .A2(SubCellInst2_LFInst_11_n29 ), .ZN(SubCellInst2_LFInst_11_n35 )
         );
  INV_X1 SubCellInst2_LFInst_11_U6  ( .A(PermutationOutput2[46]), .ZN(
        SubCellInst2_LFInst_11_n23 ) );
  NAND2_X1 SubCellInst2_LFInst_11_U5  ( .A1(SubCellInst2_LFInst_11_n29 ), 
        .A2(SubCellInst2_LFInst_11_n33 ), .ZN(SubCellInst2_LFInst_11_n26 )
         );
  INV_X1 SubCellInst2_LFInst_11_U4  ( .A(PermutationOutput2[44]), .ZN(
        SubCellInst2_LFInst_11_n33 ) );
  INV_X1 SubCellInst2_LFInst_11_U3  ( .A(PermutationOutput2[47]), .ZN(
        SubCellInst2_LFInst_11_n29 ) );
  NOR2_X1 SubCellInst2_LFInst_12_U21  ( .A1(SubCellInst2_LFInst_12_n36 ), 
        .A2(SubCellInst2_LFInst_12_n35 ), .ZN(Output[48]) );
  NOR2_X1 SubCellInst2_LFInst_12_U20  ( .A1(PermutationOutput2[49]), .A2(
        SubCellInst2_LFInst_12_n34 ), .ZN(SubCellInst2_LFInst_12_n36 ) );
  NOR2_X1 SubCellInst2_LFInst_12_U19  ( .A1(SubCellInst2_LFInst_12_n33 ), 
        .A2(SubCellInst2_LFInst_12_n32 ), .ZN(SubCellInst2_LFInst_12_n34 )
         );
  NOR2_X1 SubCellInst2_LFInst_12_U18  ( .A1(PermutationOutput2[50]), .A2(
        PermutationOutput2[51]), .ZN(SubCellInst2_LFInst_12_n32 ) );
  NAND2_X1 SubCellInst2_LFInst_12_U17  ( .A1(SubCellInst2_LFInst_12_n31 ), 
        .A2(SubCellInst2_LFInst_12_n30 ), .ZN(Output[49]) );
  NAND2_X1 SubCellInst2_LFInst_12_U16  ( .A1(PermutationOutput2[48]), .A2(
        SubCellInst2_LFInst_12_n29 ), .ZN(SubCellInst2_LFInst_12_n30 ) );
  NAND2_X1 SubCellInst2_LFInst_12_U15  ( .A1(PermutationOutput2[50]), .A2(
        SubCellInst2_LFInst_12_n28 ), .ZN(SubCellInst2_LFInst_12_n31 ) );
  NAND2_X1 SubCellInst2_LFInst_12_U14  ( .A1(PermutationOutput2[51]), .A2(
        SubCellInst2_LFInst_12_n33 ), .ZN(SubCellInst2_LFInst_12_n28 ) );
  NAND2_X1 SubCellInst2_LFInst_12_U13  ( .A1(SubCellInst2_LFInst_12_n27 ), 
        .A2(SubCellInst2_LFInst_12_n26 ), .ZN(Output[50]) );
  NAND2_X1 SubCellInst2_LFInst_12_U12  ( .A1(SubCellInst2_LFInst_12_n25 ), 
        .A2(PermutationOutput2[49]), .ZN(SubCellInst2_LFInst_12_n27 ) );
  NAND2_X1 SubCellInst2_LFInst_12_U11  ( .A1(SubCellInst2_LFInst_12_n24 ), 
        .A2(SubCellInst2_LFInst_12_n23 ), .ZN(SubCellInst2_LFInst_12_n25 )
         );
  NAND2_X1 SubCellInst2_LFInst_12_U10  ( .A1(PermutationOutput2[48]), .A2(
        PermutationOutput2[51]), .ZN(SubCellInst2_LFInst_12_n24 ) );
  NAND2_X1 SubCellInst2_LFInst_12_U9  ( .A1(SubCellInst2_LFInst_12_n26 ), 
        .A2(SubCellInst2_LFInst_12_n22 ), .ZN(Output[51]) );
  OR2_X1 SubCellInst2_LFInst_12_U8  ( .A1(PermutationOutput2[49]), .A2(
        SubCellInst2_LFInst_12_n35 ), .ZN(SubCellInst2_LFInst_12_n22 ) );
  NOR2_X1 SubCellInst2_LFInst_12_U7  ( .A1(SubCellInst2_LFInst_12_n23 ), 
        .A2(SubCellInst2_LFInst_12_n29 ), .ZN(SubCellInst2_LFInst_12_n35 )
         );
  INV_X1 SubCellInst2_LFInst_12_U6  ( .A(PermutationOutput2[50]), .ZN(
        SubCellInst2_LFInst_12_n23 ) );
  NAND2_X1 SubCellInst2_LFInst_12_U5  ( .A1(SubCellInst2_LFInst_12_n29 ), 
        .A2(SubCellInst2_LFInst_12_n33 ), .ZN(SubCellInst2_LFInst_12_n26 )
         );
  INV_X1 SubCellInst2_LFInst_12_U4  ( .A(PermutationOutput2[48]), .ZN(
        SubCellInst2_LFInst_12_n33 ) );
  INV_X1 SubCellInst2_LFInst_12_U3  ( .A(PermutationOutput2[51]), .ZN(
        SubCellInst2_LFInst_12_n29 ) );
  NOR2_X1 SubCellInst2_LFInst_13_U21  ( .A1(SubCellInst2_LFInst_13_n36 ), 
        .A2(SubCellInst2_LFInst_13_n35 ), .ZN(Output[52]) );
  NOR2_X1 SubCellInst2_LFInst_13_U20  ( .A1(PermutationOutput2[53]), .A2(
        SubCellInst2_LFInst_13_n34 ), .ZN(SubCellInst2_LFInst_13_n36 ) );
  NOR2_X1 SubCellInst2_LFInst_13_U19  ( .A1(SubCellInst2_LFInst_13_n33 ), 
        .A2(SubCellInst2_LFInst_13_n32 ), .ZN(SubCellInst2_LFInst_13_n34 )
         );
  NOR2_X1 SubCellInst2_LFInst_13_U18  ( .A1(PermutationOutput2[54]), .A2(
        PermutationOutput2[55]), .ZN(SubCellInst2_LFInst_13_n32 ) );
  NAND2_X1 SubCellInst2_LFInst_13_U17  ( .A1(SubCellInst2_LFInst_13_n31 ), 
        .A2(SubCellInst2_LFInst_13_n30 ), .ZN(Output[53]) );
  NAND2_X1 SubCellInst2_LFInst_13_U16  ( .A1(PermutationOutput2[52]), .A2(
        SubCellInst2_LFInst_13_n29 ), .ZN(SubCellInst2_LFInst_13_n30 ) );
  NAND2_X1 SubCellInst2_LFInst_13_U15  ( .A1(PermutationOutput2[54]), .A2(
        SubCellInst2_LFInst_13_n28 ), .ZN(SubCellInst2_LFInst_13_n31 ) );
  NAND2_X1 SubCellInst2_LFInst_13_U14  ( .A1(PermutationOutput2[55]), .A2(
        SubCellInst2_LFInst_13_n33 ), .ZN(SubCellInst2_LFInst_13_n28 ) );
  NAND2_X1 SubCellInst2_LFInst_13_U13  ( .A1(SubCellInst2_LFInst_13_n27 ), 
        .A2(SubCellInst2_LFInst_13_n26 ), .ZN(Output[54]) );
  NAND2_X1 SubCellInst2_LFInst_13_U12  ( .A1(SubCellInst2_LFInst_13_n25 ), 
        .A2(PermutationOutput2[53]), .ZN(SubCellInst2_LFInst_13_n27 ) );
  NAND2_X1 SubCellInst2_LFInst_13_U11  ( .A1(SubCellInst2_LFInst_13_n24 ), 
        .A2(SubCellInst2_LFInst_13_n23 ), .ZN(SubCellInst2_LFInst_13_n25 )
         );
  NAND2_X1 SubCellInst2_LFInst_13_U10  ( .A1(PermutationOutput2[52]), .A2(
        PermutationOutput2[55]), .ZN(SubCellInst2_LFInst_13_n24 ) );
  NAND2_X1 SubCellInst2_LFInst_13_U9  ( .A1(SubCellInst2_LFInst_13_n26 ), 
        .A2(SubCellInst2_LFInst_13_n22 ), .ZN(Output[55]) );
  OR2_X1 SubCellInst2_LFInst_13_U8  ( .A1(PermutationOutput2[53]), .A2(
        SubCellInst2_LFInst_13_n35 ), .ZN(SubCellInst2_LFInst_13_n22 ) );
  NOR2_X1 SubCellInst2_LFInst_13_U7  ( .A1(SubCellInst2_LFInst_13_n23 ), 
        .A2(SubCellInst2_LFInst_13_n29 ), .ZN(SubCellInst2_LFInst_13_n35 )
         );
  INV_X1 SubCellInst2_LFInst_13_U6  ( .A(PermutationOutput2[54]), .ZN(
        SubCellInst2_LFInst_13_n23 ) );
  NAND2_X1 SubCellInst2_LFInst_13_U5  ( .A1(SubCellInst2_LFInst_13_n29 ), 
        .A2(SubCellInst2_LFInst_13_n33 ), .ZN(SubCellInst2_LFInst_13_n26 )
         );
  INV_X1 SubCellInst2_LFInst_13_U4  ( .A(PermutationOutput2[52]), .ZN(
        SubCellInst2_LFInst_13_n33 ) );
  INV_X1 SubCellInst2_LFInst_13_U3  ( .A(PermutationOutput2[55]), .ZN(
        SubCellInst2_LFInst_13_n29 ) );
  NOR2_X1 SubCellInst2_LFInst_14_U21  ( .A1(SubCellInst2_LFInst_14_n36 ), 
        .A2(SubCellInst2_LFInst_14_n35 ), .ZN(Output[56]) );
  NOR2_X1 SubCellInst2_LFInst_14_U20  ( .A1(PermutationOutput2[57]), .A2(
        SubCellInst2_LFInst_14_n34 ), .ZN(SubCellInst2_LFInst_14_n36 ) );
  NOR2_X1 SubCellInst2_LFInst_14_U19  ( .A1(SubCellInst2_LFInst_14_n33 ), 
        .A2(SubCellInst2_LFInst_14_n32 ), .ZN(SubCellInst2_LFInst_14_n34 )
         );
  NOR2_X1 SubCellInst2_LFInst_14_U18  ( .A1(PermutationOutput2[58]), .A2(
        PermutationOutput2[59]), .ZN(SubCellInst2_LFInst_14_n32 ) );
  NAND2_X1 SubCellInst2_LFInst_14_U17  ( .A1(SubCellInst2_LFInst_14_n31 ), 
        .A2(SubCellInst2_LFInst_14_n30 ), .ZN(Output[57]) );
  NAND2_X1 SubCellInst2_LFInst_14_U16  ( .A1(PermutationOutput2[56]), .A2(
        SubCellInst2_LFInst_14_n29 ), .ZN(SubCellInst2_LFInst_14_n30 ) );
  NAND2_X1 SubCellInst2_LFInst_14_U15  ( .A1(PermutationOutput2[58]), .A2(
        SubCellInst2_LFInst_14_n28 ), .ZN(SubCellInst2_LFInst_14_n31 ) );
  NAND2_X1 SubCellInst2_LFInst_14_U14  ( .A1(PermutationOutput2[59]), .A2(
        SubCellInst2_LFInst_14_n33 ), .ZN(SubCellInst2_LFInst_14_n28 ) );
  NAND2_X1 SubCellInst2_LFInst_14_U13  ( .A1(SubCellInst2_LFInst_14_n27 ), 
        .A2(SubCellInst2_LFInst_14_n26 ), .ZN(Output[58]) );
  NAND2_X1 SubCellInst2_LFInst_14_U12  ( .A1(SubCellInst2_LFInst_14_n25 ), 
        .A2(PermutationOutput2[57]), .ZN(SubCellInst2_LFInst_14_n27 ) );
  NAND2_X1 SubCellInst2_LFInst_14_U11  ( .A1(SubCellInst2_LFInst_14_n24 ), 
        .A2(SubCellInst2_LFInst_14_n23 ), .ZN(SubCellInst2_LFInst_14_n25 )
         );
  NAND2_X1 SubCellInst2_LFInst_14_U10  ( .A1(PermutationOutput2[56]), .A2(
        PermutationOutput2[59]), .ZN(SubCellInst2_LFInst_14_n24 ) );
  NAND2_X1 SubCellInst2_LFInst_14_U9  ( .A1(SubCellInst2_LFInst_14_n26 ), 
        .A2(SubCellInst2_LFInst_14_n22 ), .ZN(Output[59]) );
  OR2_X1 SubCellInst2_LFInst_14_U8  ( .A1(PermutationOutput2[57]), .A2(
        SubCellInst2_LFInst_14_n35 ), .ZN(SubCellInst2_LFInst_14_n22 ) );
  NOR2_X1 SubCellInst2_LFInst_14_U7  ( .A1(SubCellInst2_LFInst_14_n23 ), 
        .A2(SubCellInst2_LFInst_14_n29 ), .ZN(SubCellInst2_LFInst_14_n35 )
         );
  INV_X1 SubCellInst2_LFInst_14_U6  ( .A(PermutationOutput2[58]), .ZN(
        SubCellInst2_LFInst_14_n23 ) );
  NAND2_X1 SubCellInst2_LFInst_14_U5  ( .A1(SubCellInst2_LFInst_14_n29 ), 
        .A2(SubCellInst2_LFInst_14_n33 ), .ZN(SubCellInst2_LFInst_14_n26 )
         );
  INV_X1 SubCellInst2_LFInst_14_U4  ( .A(PermutationOutput2[56]), .ZN(
        SubCellInst2_LFInst_14_n33 ) );
  INV_X1 SubCellInst2_LFInst_14_U3  ( .A(PermutationOutput2[59]), .ZN(
        SubCellInst2_LFInst_14_n29 ) );
  NOR2_X1 SubCellInst2_LFInst_15_U21  ( .A1(SubCellInst2_LFInst_15_n36 ), 
        .A2(SubCellInst2_LFInst_15_n35 ), .ZN(Output[60]) );
  NOR2_X1 SubCellInst2_LFInst_15_U20  ( .A1(PermutationOutput2[61]), .A2(
        SubCellInst2_LFInst_15_n34 ), .ZN(SubCellInst2_LFInst_15_n36 ) );
  NOR2_X1 SubCellInst2_LFInst_15_U19  ( .A1(SubCellInst2_LFInst_15_n33 ), 
        .A2(SubCellInst2_LFInst_15_n32 ), .ZN(SubCellInst2_LFInst_15_n34 )
         );
  NOR2_X1 SubCellInst2_LFInst_15_U18  ( .A1(PermutationOutput2[62]), .A2(
        PermutationOutput2[63]), .ZN(SubCellInst2_LFInst_15_n32 ) );
  NAND2_X1 SubCellInst2_LFInst_15_U17  ( .A1(SubCellInst2_LFInst_15_n31 ), 
        .A2(SubCellInst2_LFInst_15_n30 ), .ZN(Output[61]) );
  NAND2_X1 SubCellInst2_LFInst_15_U16  ( .A1(PermutationOutput2[60]), .A2(
        SubCellInst2_LFInst_15_n29 ), .ZN(SubCellInst2_LFInst_15_n30 ) );
  NAND2_X1 SubCellInst2_LFInst_15_U15  ( .A1(PermutationOutput2[62]), .A2(
        SubCellInst2_LFInst_15_n28 ), .ZN(SubCellInst2_LFInst_15_n31 ) );
  NAND2_X1 SubCellInst2_LFInst_15_U14  ( .A1(PermutationOutput2[63]), .A2(
        SubCellInst2_LFInst_15_n33 ), .ZN(SubCellInst2_LFInst_15_n28 ) );
  NAND2_X1 SubCellInst2_LFInst_15_U13  ( .A1(SubCellInst2_LFInst_15_n27 ), 
        .A2(SubCellInst2_LFInst_15_n26 ), .ZN(Output[62]) );
  NAND2_X1 SubCellInst2_LFInst_15_U12  ( .A1(SubCellInst2_LFInst_15_n25 ), 
        .A2(PermutationOutput2[61]), .ZN(SubCellInst2_LFInst_15_n27 ) );
  NAND2_X1 SubCellInst2_LFInst_15_U11  ( .A1(SubCellInst2_LFInst_15_n24 ), 
        .A2(SubCellInst2_LFInst_15_n23 ), .ZN(SubCellInst2_LFInst_15_n25 )
         );
  NAND2_X1 SubCellInst2_LFInst_15_U10  ( .A1(PermutationOutput2[60]), .A2(
        PermutationOutput2[63]), .ZN(SubCellInst2_LFInst_15_n24 ) );
  NAND2_X1 SubCellInst2_LFInst_15_U9  ( .A1(SubCellInst2_LFInst_15_n26 ), 
        .A2(SubCellInst2_LFInst_15_n22 ), .ZN(Output[63]) );
  OR2_X1 SubCellInst2_LFInst_15_U8  ( .A1(PermutationOutput2[61]), .A2(
        SubCellInst2_LFInst_15_n35 ), .ZN(SubCellInst2_LFInst_15_n22 ) );
  NOR2_X1 SubCellInst2_LFInst_15_U7  ( .A1(SubCellInst2_LFInst_15_n23 ), 
        .A2(SubCellInst2_LFInst_15_n29 ), .ZN(SubCellInst2_LFInst_15_n35 )
         );
  INV_X1 SubCellInst2_LFInst_15_U6  ( .A(PermutationOutput2[62]), .ZN(
        SubCellInst2_LFInst_15_n23 ) );
  NAND2_X1 SubCellInst2_LFInst_15_U5  ( .A1(SubCellInst2_LFInst_15_n29 ), 
        .A2(SubCellInst2_LFInst_15_n33 ), .ZN(SubCellInst2_LFInst_15_n26 )
         );
  INV_X1 SubCellInst2_LFInst_15_U4  ( .A(PermutationOutput2[60]), .ZN(
        SubCellInst2_LFInst_15_n33 ) );
  INV_X1 SubCellInst2_LFInst_15_U3  ( .A(PermutationOutput2[63]), .ZN(
        SubCellInst2_LFInst_15_n29 ) );
endmodule

