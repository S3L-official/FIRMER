module LED64Enc ( clk, rst, Plaintext, Key, Ciphertext, ErrorFlag );
  input [63:0] Plaintext;
  input [63:0] Key;
  output [63:0] Ciphertext;
  (* FIRMER="clock" *)input clk;
  (* FIRMER="control" *)input rst;
  output ErrorFlag;
  wire   n149, \AddKeyXOR_XORInst_0_0_n2 , \AddKeyXOR_XORInst_0_2_n2 ,
         \AddKeyXOR_XORInst_1_2_n2 , \AddKeyXOR_XORInst_2_2_n2 ,
         \AddKeyXOR_XORInst_3_2_n2 , \AddKeyXOR_XORInst_4_2_n2 ,
         \AddKeyXOR_XORInst_5_2_n2 , \AddKeyXOR_XORInst_6_2_n2 ,
         \AddKeyXOR_XORInst_7_2_n2 , \AddKeyXOR_XORInst_8_2_n2 ,
         \AddKeyXOR_XORInst_9_2_n2 , \AddKeyXOR_XORInst_10_2_n2 ,
         \AddKeyXOR_XORInst_11_2_n2 , \AddKeyXOR_XORInst_12_2_n2 ,
         \AddKeyXOR_XORInst_13_2_n2 , \AddKeyXOR_XORInst_14_2_n2 ,
         \AddKeyXOR_XORInst_15_2_n2 , \SubCellInst_LFInst_0_LFInst_0_n9 ,
         \SubCellInst_LFInst_0_LFInst_0_n8 ,
         \SubCellInst_LFInst_0_LFInst_0_n7 ,
         \SubCellInst_LFInst_0_LFInst_0_n10 ,
         \SubCellInst_LFInst_0_LFInst_1_n18 ,
         \SubCellInst_LFInst_0_LFInst_1_n17 ,
         \SubCellInst_LFInst_0_LFInst_1_n16 ,
         \SubCellInst_LFInst_0_LFInst_1_n15 ,
         \SubCellInst_LFInst_0_LFInst_1_n14 ,
         \SubCellInst_LFInst_0_LFInst_1_n13 ,
         \SubCellInst_LFInst_0_LFInst_1_n12 ,
         \SubCellInst_LFInst_0_LFInst_1_n11 ,
         \SubCellInst_LFInst_0_LFInst_1_n10 ,
         \SubCellInst_LFInst_0_LFInst_2_n22 ,
         \SubCellInst_LFInst_0_LFInst_2_n21 ,
         \SubCellInst_LFInst_0_LFInst_2_n20 ,
         \SubCellInst_LFInst_0_LFInst_2_n19 ,
         \SubCellInst_LFInst_0_LFInst_2_n18 ,
         \SubCellInst_LFInst_0_LFInst_2_n17 ,
         \SubCellInst_LFInst_0_LFInst_2_n16 ,
         \SubCellInst_LFInst_0_LFInst_2_n15 ,
         \SubCellInst_LFInst_0_LFInst_3_n16 ,
         \SubCellInst_LFInst_0_LFInst_3_n15 ,
         \SubCellInst_LFInst_0_LFInst_3_n14 ,
         \SubCellInst_LFInst_0_LFInst_3_n13 ,
         \SubCellInst_LFInst_0_LFInst_3_n12 ,
         \SubCellInst_LFInst_0_LFInst_3_n11 ,
         \SubCellInst_LFInst_1_LFInst_0_n10 ,
         \SubCellInst_LFInst_1_LFInst_0_n9 ,
         \SubCellInst_LFInst_1_LFInst_0_n8 ,
         \SubCellInst_LFInst_1_LFInst_0_n7 ,
         \SubCellInst_LFInst_1_LFInst_1_n18 ,
         \SubCellInst_LFInst_1_LFInst_1_n17 ,
         \SubCellInst_LFInst_1_LFInst_1_n16 ,
         \SubCellInst_LFInst_1_LFInst_1_n15 ,
         \SubCellInst_LFInst_1_LFInst_1_n14 ,
         \SubCellInst_LFInst_1_LFInst_1_n13 ,
         \SubCellInst_LFInst_1_LFInst_1_n12 ,
         \SubCellInst_LFInst_1_LFInst_1_n11 ,
         \SubCellInst_LFInst_1_LFInst_1_n10 ,
         \SubCellInst_LFInst_1_LFInst_2_n22 ,
         \SubCellInst_LFInst_1_LFInst_2_n21 ,
         \SubCellInst_LFInst_1_LFInst_2_n20 ,
         \SubCellInst_LFInst_1_LFInst_2_n19 ,
         \SubCellInst_LFInst_1_LFInst_2_n18 ,
         \SubCellInst_LFInst_1_LFInst_2_n17 ,
         \SubCellInst_LFInst_1_LFInst_2_n16 ,
         \SubCellInst_LFInst_1_LFInst_2_n15 ,
         \SubCellInst_LFInst_1_LFInst_3_n16 ,
         \SubCellInst_LFInst_1_LFInst_3_n15 ,
         \SubCellInst_LFInst_1_LFInst_3_n14 ,
         \SubCellInst_LFInst_1_LFInst_3_n13 ,
         \SubCellInst_LFInst_1_LFInst_3_n12 ,
         \SubCellInst_LFInst_1_LFInst_3_n11 ,
         \SubCellInst_LFInst_2_LFInst_0_n10 ,
         \SubCellInst_LFInst_2_LFInst_0_n9 ,
         \SubCellInst_LFInst_2_LFInst_0_n8 ,
         \SubCellInst_LFInst_2_LFInst_0_n7 ,
         \SubCellInst_LFInst_2_LFInst_1_n18 ,
         \SubCellInst_LFInst_2_LFInst_1_n17 ,
         \SubCellInst_LFInst_2_LFInst_1_n16 ,
         \SubCellInst_LFInst_2_LFInst_1_n15 ,
         \SubCellInst_LFInst_2_LFInst_1_n14 ,
         \SubCellInst_LFInst_2_LFInst_1_n13 ,
         \SubCellInst_LFInst_2_LFInst_1_n12 ,
         \SubCellInst_LFInst_2_LFInst_1_n11 ,
         \SubCellInst_LFInst_2_LFInst_1_n10 ,
         \SubCellInst_LFInst_2_LFInst_2_n22 ,
         \SubCellInst_LFInst_2_LFInst_2_n21 ,
         \SubCellInst_LFInst_2_LFInst_2_n20 ,
         \SubCellInst_LFInst_2_LFInst_2_n19 ,
         \SubCellInst_LFInst_2_LFInst_2_n18 ,
         \SubCellInst_LFInst_2_LFInst_2_n17 ,
         \SubCellInst_LFInst_2_LFInst_2_n16 ,
         \SubCellInst_LFInst_2_LFInst_2_n15 ,
         \SubCellInst_LFInst_2_LFInst_3_n16 ,
         \SubCellInst_LFInst_2_LFInst_3_n15 ,
         \SubCellInst_LFInst_2_LFInst_3_n14 ,
         \SubCellInst_LFInst_2_LFInst_3_n13 ,
         \SubCellInst_LFInst_2_LFInst_3_n12 ,
         \SubCellInst_LFInst_2_LFInst_3_n11 ,
         \SubCellInst_LFInst_3_LFInst_0_n10 ,
         \SubCellInst_LFInst_3_LFInst_0_n9 ,
         \SubCellInst_LFInst_3_LFInst_0_n8 ,
         \SubCellInst_LFInst_3_LFInst_0_n7 ,
         \SubCellInst_LFInst_3_LFInst_1_n18 ,
         \SubCellInst_LFInst_3_LFInst_1_n17 ,
         \SubCellInst_LFInst_3_LFInst_1_n16 ,
         \SubCellInst_LFInst_3_LFInst_1_n15 ,
         \SubCellInst_LFInst_3_LFInst_1_n14 ,
         \SubCellInst_LFInst_3_LFInst_1_n13 ,
         \SubCellInst_LFInst_3_LFInst_1_n12 ,
         \SubCellInst_LFInst_3_LFInst_1_n11 ,
         \SubCellInst_LFInst_3_LFInst_1_n10 ,
         \SubCellInst_LFInst_3_LFInst_2_n22 ,
         \SubCellInst_LFInst_3_LFInst_2_n21 ,
         \SubCellInst_LFInst_3_LFInst_2_n20 ,
         \SubCellInst_LFInst_3_LFInst_2_n19 ,
         \SubCellInst_LFInst_3_LFInst_2_n18 ,
         \SubCellInst_LFInst_3_LFInst_2_n17 ,
         \SubCellInst_LFInst_3_LFInst_2_n16 ,
         \SubCellInst_LFInst_3_LFInst_2_n15 ,
         \SubCellInst_LFInst_3_LFInst_3_n16 ,
         \SubCellInst_LFInst_3_LFInst_3_n15 ,
         \SubCellInst_LFInst_3_LFInst_3_n14 ,
         \SubCellInst_LFInst_3_LFInst_3_n13 ,
         \SubCellInst_LFInst_3_LFInst_3_n12 ,
         \SubCellInst_LFInst_3_LFInst_3_n11 ,
         \SubCellInst_LFInst_4_LFInst_0_n9 ,
         \SubCellInst_LFInst_4_LFInst_0_n8 ,
         \SubCellInst_LFInst_4_LFInst_0_n7 ,
         \SubCellInst_LFInst_4_LFInst_0_n10 ,
         \SubCellInst_LFInst_4_LFInst_1_n18 ,
         \SubCellInst_LFInst_4_LFInst_1_n17 ,
         \SubCellInst_LFInst_4_LFInst_1_n16 ,
         \SubCellInst_LFInst_4_LFInst_1_n15 ,
         \SubCellInst_LFInst_4_LFInst_1_n14 ,
         \SubCellInst_LFInst_4_LFInst_1_n13 ,
         \SubCellInst_LFInst_4_LFInst_1_n12 ,
         \SubCellInst_LFInst_4_LFInst_1_n11 ,
         \SubCellInst_LFInst_4_LFInst_1_n10 ,
         \SubCellInst_LFInst_4_LFInst_2_n22 ,
         \SubCellInst_LFInst_4_LFInst_2_n21 ,
         \SubCellInst_LFInst_4_LFInst_2_n20 ,
         \SubCellInst_LFInst_4_LFInst_2_n19 ,
         \SubCellInst_LFInst_4_LFInst_2_n18 ,
         \SubCellInst_LFInst_4_LFInst_2_n17 ,
         \SubCellInst_LFInst_4_LFInst_2_n16 ,
         \SubCellInst_LFInst_4_LFInst_2_n15 ,
         \SubCellInst_LFInst_4_LFInst_3_n16 ,
         \SubCellInst_LFInst_4_LFInst_3_n15 ,
         \SubCellInst_LFInst_4_LFInst_3_n14 ,
         \SubCellInst_LFInst_4_LFInst_3_n13 ,
         \SubCellInst_LFInst_4_LFInst_3_n12 ,
         \SubCellInst_LFInst_4_LFInst_3_n11 ,
         \SubCellInst_LFInst_5_LFInst_0_n10 ,
         \SubCellInst_LFInst_5_LFInst_0_n9 ,
         \SubCellInst_LFInst_5_LFInst_0_n8 ,
         \SubCellInst_LFInst_5_LFInst_0_n7 ,
         \SubCellInst_LFInst_5_LFInst_1_n18 ,
         \SubCellInst_LFInst_5_LFInst_1_n17 ,
         \SubCellInst_LFInst_5_LFInst_1_n16 ,
         \SubCellInst_LFInst_5_LFInst_1_n15 ,
         \SubCellInst_LFInst_5_LFInst_1_n14 ,
         \SubCellInst_LFInst_5_LFInst_1_n13 ,
         \SubCellInst_LFInst_5_LFInst_1_n12 ,
         \SubCellInst_LFInst_5_LFInst_1_n11 ,
         \SubCellInst_LFInst_5_LFInst_1_n10 ,
         \SubCellInst_LFInst_5_LFInst_2_n22 ,
         \SubCellInst_LFInst_5_LFInst_2_n21 ,
         \SubCellInst_LFInst_5_LFInst_2_n20 ,
         \SubCellInst_LFInst_5_LFInst_2_n19 ,
         \SubCellInst_LFInst_5_LFInst_2_n18 ,
         \SubCellInst_LFInst_5_LFInst_2_n17 ,
         \SubCellInst_LFInst_5_LFInst_2_n16 ,
         \SubCellInst_LFInst_5_LFInst_2_n15 ,
         \SubCellInst_LFInst_5_LFInst_3_n16 ,
         \SubCellInst_LFInst_5_LFInst_3_n15 ,
         \SubCellInst_LFInst_5_LFInst_3_n14 ,
         \SubCellInst_LFInst_5_LFInst_3_n13 ,
         \SubCellInst_LFInst_5_LFInst_3_n12 ,
         \SubCellInst_LFInst_5_LFInst_3_n11 ,
         \SubCellInst_LFInst_6_LFInst_0_n10 ,
         \SubCellInst_LFInst_6_LFInst_0_n9 ,
         \SubCellInst_LFInst_6_LFInst_0_n8 ,
         \SubCellInst_LFInst_6_LFInst_0_n7 ,
         \SubCellInst_LFInst_6_LFInst_1_n18 ,
         \SubCellInst_LFInst_6_LFInst_1_n17 ,
         \SubCellInst_LFInst_6_LFInst_1_n16 ,
         \SubCellInst_LFInst_6_LFInst_1_n15 ,
         \SubCellInst_LFInst_6_LFInst_1_n14 ,
         \SubCellInst_LFInst_6_LFInst_1_n13 ,
         \SubCellInst_LFInst_6_LFInst_1_n12 ,
         \SubCellInst_LFInst_6_LFInst_1_n11 ,
         \SubCellInst_LFInst_6_LFInst_1_n10 ,
         \SubCellInst_LFInst_6_LFInst_2_n22 ,
         \SubCellInst_LFInst_6_LFInst_2_n21 ,
         \SubCellInst_LFInst_6_LFInst_2_n20 ,
         \SubCellInst_LFInst_6_LFInst_2_n19 ,
         \SubCellInst_LFInst_6_LFInst_2_n18 ,
         \SubCellInst_LFInst_6_LFInst_2_n17 ,
         \SubCellInst_LFInst_6_LFInst_2_n16 ,
         \SubCellInst_LFInst_6_LFInst_2_n15 ,
         \SubCellInst_LFInst_6_LFInst_3_n16 ,
         \SubCellInst_LFInst_6_LFInst_3_n15 ,
         \SubCellInst_LFInst_6_LFInst_3_n14 ,
         \SubCellInst_LFInst_6_LFInst_3_n13 ,
         \SubCellInst_LFInst_6_LFInst_3_n12 ,
         \SubCellInst_LFInst_6_LFInst_3_n11 ,
         \SubCellInst_LFInst_7_LFInst_0_n10 ,
         \SubCellInst_LFInst_7_LFInst_0_n9 ,
         \SubCellInst_LFInst_7_LFInst_0_n8 ,
         \SubCellInst_LFInst_7_LFInst_0_n7 ,
         \SubCellInst_LFInst_7_LFInst_1_n18 ,
         \SubCellInst_LFInst_7_LFInst_1_n17 ,
         \SubCellInst_LFInst_7_LFInst_1_n16 ,
         \SubCellInst_LFInst_7_LFInst_1_n15 ,
         \SubCellInst_LFInst_7_LFInst_1_n14 ,
         \SubCellInst_LFInst_7_LFInst_1_n13 ,
         \SubCellInst_LFInst_7_LFInst_1_n12 ,
         \SubCellInst_LFInst_7_LFInst_1_n11 ,
         \SubCellInst_LFInst_7_LFInst_1_n10 ,
         \SubCellInst_LFInst_7_LFInst_2_n22 ,
         \SubCellInst_LFInst_7_LFInst_2_n21 ,
         \SubCellInst_LFInst_7_LFInst_2_n20 ,
         \SubCellInst_LFInst_7_LFInst_2_n19 ,
         \SubCellInst_LFInst_7_LFInst_2_n18 ,
         \SubCellInst_LFInst_7_LFInst_2_n17 ,
         \SubCellInst_LFInst_7_LFInst_2_n16 ,
         \SubCellInst_LFInst_7_LFInst_2_n15 ,
         \SubCellInst_LFInst_7_LFInst_3_n16 ,
         \SubCellInst_LFInst_7_LFInst_3_n15 ,
         \SubCellInst_LFInst_7_LFInst_3_n14 ,
         \SubCellInst_LFInst_7_LFInst_3_n13 ,
         \SubCellInst_LFInst_7_LFInst_3_n12 ,
         \SubCellInst_LFInst_7_LFInst_3_n11 ,
         \SubCellInst_LFInst_8_LFInst_0_n10 ,
         \SubCellInst_LFInst_8_LFInst_0_n9 ,
         \SubCellInst_LFInst_8_LFInst_0_n8 ,
         \SubCellInst_LFInst_8_LFInst_0_n7 ,
         \SubCellInst_LFInst_8_LFInst_1_n18 ,
         \SubCellInst_LFInst_8_LFInst_1_n17 ,
         \SubCellInst_LFInst_8_LFInst_1_n16 ,
         \SubCellInst_LFInst_8_LFInst_1_n15 ,
         \SubCellInst_LFInst_8_LFInst_1_n14 ,
         \SubCellInst_LFInst_8_LFInst_1_n13 ,
         \SubCellInst_LFInst_8_LFInst_1_n12 ,
         \SubCellInst_LFInst_8_LFInst_1_n11 ,
         \SubCellInst_LFInst_8_LFInst_1_n10 ,
         \SubCellInst_LFInst_8_LFInst_2_n22 ,
         \SubCellInst_LFInst_8_LFInst_2_n21 ,
         \SubCellInst_LFInst_8_LFInst_2_n20 ,
         \SubCellInst_LFInst_8_LFInst_2_n19 ,
         \SubCellInst_LFInst_8_LFInst_2_n18 ,
         \SubCellInst_LFInst_8_LFInst_2_n17 ,
         \SubCellInst_LFInst_8_LFInst_2_n16 ,
         \SubCellInst_LFInst_8_LFInst_2_n15 ,
         \SubCellInst_LFInst_8_LFInst_3_n16 ,
         \SubCellInst_LFInst_8_LFInst_3_n15 ,
         \SubCellInst_LFInst_8_LFInst_3_n14 ,
         \SubCellInst_LFInst_8_LFInst_3_n13 ,
         \SubCellInst_LFInst_8_LFInst_3_n12 ,
         \SubCellInst_LFInst_8_LFInst_3_n11 ,
         \SubCellInst_LFInst_9_LFInst_0_n10 ,
         \SubCellInst_LFInst_9_LFInst_0_n9 ,
         \SubCellInst_LFInst_9_LFInst_0_n8 ,
         \SubCellInst_LFInst_9_LFInst_0_n7 ,
         \SubCellInst_LFInst_9_LFInst_1_n18 ,
         \SubCellInst_LFInst_9_LFInst_1_n17 ,
         \SubCellInst_LFInst_9_LFInst_1_n16 ,
         \SubCellInst_LFInst_9_LFInst_1_n15 ,
         \SubCellInst_LFInst_9_LFInst_1_n14 ,
         \SubCellInst_LFInst_9_LFInst_1_n13 ,
         \SubCellInst_LFInst_9_LFInst_1_n12 ,
         \SubCellInst_LFInst_9_LFInst_1_n11 ,
         \SubCellInst_LFInst_9_LFInst_1_n10 ,
         \SubCellInst_LFInst_9_LFInst_2_n22 ,
         \SubCellInst_LFInst_9_LFInst_2_n21 ,
         \SubCellInst_LFInst_9_LFInst_2_n20 ,
         \SubCellInst_LFInst_9_LFInst_2_n19 ,
         \SubCellInst_LFInst_9_LFInst_2_n18 ,
         \SubCellInst_LFInst_9_LFInst_2_n17 ,
         \SubCellInst_LFInst_9_LFInst_2_n16 ,
         \SubCellInst_LFInst_9_LFInst_2_n15 ,
         \SubCellInst_LFInst_9_LFInst_3_n16 ,
         \SubCellInst_LFInst_9_LFInst_3_n15 ,
         \SubCellInst_LFInst_9_LFInst_3_n14 ,
         \SubCellInst_LFInst_9_LFInst_3_n13 ,
         \SubCellInst_LFInst_9_LFInst_3_n12 ,
         \SubCellInst_LFInst_9_LFInst_3_n11 ,
         \SubCellInst_LFInst_10_LFInst_0_n10 ,
         \SubCellInst_LFInst_10_LFInst_0_n9 ,
         \SubCellInst_LFInst_10_LFInst_0_n8 ,
         \SubCellInst_LFInst_10_LFInst_0_n7 ,
         \SubCellInst_LFInst_10_LFInst_1_n18 ,
         \SubCellInst_LFInst_10_LFInst_1_n17 ,
         \SubCellInst_LFInst_10_LFInst_1_n16 ,
         \SubCellInst_LFInst_10_LFInst_1_n15 ,
         \SubCellInst_LFInst_10_LFInst_1_n14 ,
         \SubCellInst_LFInst_10_LFInst_1_n13 ,
         \SubCellInst_LFInst_10_LFInst_1_n12 ,
         \SubCellInst_LFInst_10_LFInst_1_n11 ,
         \SubCellInst_LFInst_10_LFInst_1_n10 ,
         \SubCellInst_LFInst_10_LFInst_2_n22 ,
         \SubCellInst_LFInst_10_LFInst_2_n21 ,
         \SubCellInst_LFInst_10_LFInst_2_n20 ,
         \SubCellInst_LFInst_10_LFInst_2_n19 ,
         \SubCellInst_LFInst_10_LFInst_2_n18 ,
         \SubCellInst_LFInst_10_LFInst_2_n17 ,
         \SubCellInst_LFInst_10_LFInst_2_n16 ,
         \SubCellInst_LFInst_10_LFInst_2_n15 ,
         \SubCellInst_LFInst_10_LFInst_3_n16 ,
         \SubCellInst_LFInst_10_LFInst_3_n15 ,
         \SubCellInst_LFInst_10_LFInst_3_n14 ,
         \SubCellInst_LFInst_10_LFInst_3_n13 ,
         \SubCellInst_LFInst_10_LFInst_3_n12 ,
         \SubCellInst_LFInst_10_LFInst_3_n11 ,
         \SubCellInst_LFInst_11_LFInst_0_n10 ,
         \SubCellInst_LFInst_11_LFInst_0_n9 ,
         \SubCellInst_LFInst_11_LFInst_0_n8 ,
         \SubCellInst_LFInst_11_LFInst_0_n7 ,
         \SubCellInst_LFInst_11_LFInst_1_n18 ,
         \SubCellInst_LFInst_11_LFInst_1_n17 ,
         \SubCellInst_LFInst_11_LFInst_1_n16 ,
         \SubCellInst_LFInst_11_LFInst_1_n15 ,
         \SubCellInst_LFInst_11_LFInst_1_n14 ,
         \SubCellInst_LFInst_11_LFInst_1_n13 ,
         \SubCellInst_LFInst_11_LFInst_1_n12 ,
         \SubCellInst_LFInst_11_LFInst_1_n11 ,
         \SubCellInst_LFInst_11_LFInst_1_n10 ,
         \SubCellInst_LFInst_11_LFInst_2_n22 ,
         \SubCellInst_LFInst_11_LFInst_2_n21 ,
         \SubCellInst_LFInst_11_LFInst_2_n20 ,
         \SubCellInst_LFInst_11_LFInst_2_n19 ,
         \SubCellInst_LFInst_11_LFInst_2_n18 ,
         \SubCellInst_LFInst_11_LFInst_2_n17 ,
         \SubCellInst_LFInst_11_LFInst_2_n16 ,
         \SubCellInst_LFInst_11_LFInst_2_n15 ,
         \SubCellInst_LFInst_11_LFInst_3_n16 ,
         \SubCellInst_LFInst_11_LFInst_3_n15 ,
         \SubCellInst_LFInst_11_LFInst_3_n14 ,
         \SubCellInst_LFInst_11_LFInst_3_n13 ,
         \SubCellInst_LFInst_11_LFInst_3_n12 ,
         \SubCellInst_LFInst_11_LFInst_3_n11 ,
         \SubCellInst_LFInst_12_LFInst_0_n10 ,
         \SubCellInst_LFInst_12_LFInst_0_n9 ,
         \SubCellInst_LFInst_12_LFInst_0_n8 ,
         \SubCellInst_LFInst_12_LFInst_0_n7 ,
         \SubCellInst_LFInst_12_LFInst_1_n18 ,
         \SubCellInst_LFInst_12_LFInst_1_n17 ,
         \SubCellInst_LFInst_12_LFInst_1_n16 ,
         \SubCellInst_LFInst_12_LFInst_1_n15 ,
         \SubCellInst_LFInst_12_LFInst_1_n14 ,
         \SubCellInst_LFInst_12_LFInst_1_n13 ,
         \SubCellInst_LFInst_12_LFInst_1_n12 ,
         \SubCellInst_LFInst_12_LFInst_1_n11 ,
         \SubCellInst_LFInst_12_LFInst_1_n10 ,
         \SubCellInst_LFInst_12_LFInst_2_n22 ,
         \SubCellInst_LFInst_12_LFInst_2_n21 ,
         \SubCellInst_LFInst_12_LFInst_2_n20 ,
         \SubCellInst_LFInst_12_LFInst_2_n19 ,
         \SubCellInst_LFInst_12_LFInst_2_n18 ,
         \SubCellInst_LFInst_12_LFInst_2_n17 ,
         \SubCellInst_LFInst_12_LFInst_2_n16 ,
         \SubCellInst_LFInst_12_LFInst_2_n15 ,
         \SubCellInst_LFInst_12_LFInst_3_n16 ,
         \SubCellInst_LFInst_12_LFInst_3_n15 ,
         \SubCellInst_LFInst_12_LFInst_3_n14 ,
         \SubCellInst_LFInst_12_LFInst_3_n13 ,
         \SubCellInst_LFInst_12_LFInst_3_n12 ,
         \SubCellInst_LFInst_12_LFInst_3_n11 ,
         \SubCellInst_LFInst_13_LFInst_0_n10 ,
         \SubCellInst_LFInst_13_LFInst_0_n9 ,
         \SubCellInst_LFInst_13_LFInst_0_n8 ,
         \SubCellInst_LFInst_13_LFInst_0_n7 ,
         \SubCellInst_LFInst_13_LFInst_1_n18 ,
         \SubCellInst_LFInst_13_LFInst_1_n17 ,
         \SubCellInst_LFInst_13_LFInst_1_n16 ,
         \SubCellInst_LFInst_13_LFInst_1_n15 ,
         \SubCellInst_LFInst_13_LFInst_1_n14 ,
         \SubCellInst_LFInst_13_LFInst_1_n13 ,
         \SubCellInst_LFInst_13_LFInst_1_n12 ,
         \SubCellInst_LFInst_13_LFInst_1_n11 ,
         \SubCellInst_LFInst_13_LFInst_1_n10 ,
         \SubCellInst_LFInst_13_LFInst_2_n22 ,
         \SubCellInst_LFInst_13_LFInst_2_n21 ,
         \SubCellInst_LFInst_13_LFInst_2_n20 ,
         \SubCellInst_LFInst_13_LFInst_2_n19 ,
         \SubCellInst_LFInst_13_LFInst_2_n18 ,
         \SubCellInst_LFInst_13_LFInst_2_n17 ,
         \SubCellInst_LFInst_13_LFInst_2_n16 ,
         \SubCellInst_LFInst_13_LFInst_2_n15 ,
         \SubCellInst_LFInst_13_LFInst_3_n16 ,
         \SubCellInst_LFInst_13_LFInst_3_n15 ,
         \SubCellInst_LFInst_13_LFInst_3_n14 ,
         \SubCellInst_LFInst_13_LFInst_3_n13 ,
         \SubCellInst_LFInst_13_LFInst_3_n12 ,
         \SubCellInst_LFInst_13_LFInst_3_n11 ,
         \SubCellInst_LFInst_14_LFInst_0_n10 ,
         \SubCellInst_LFInst_14_LFInst_0_n9 ,
         \SubCellInst_LFInst_14_LFInst_0_n8 ,
         \SubCellInst_LFInst_14_LFInst_0_n7 ,
         \SubCellInst_LFInst_14_LFInst_1_n18 ,
         \SubCellInst_LFInst_14_LFInst_1_n17 ,
         \SubCellInst_LFInst_14_LFInst_1_n16 ,
         \SubCellInst_LFInst_14_LFInst_1_n15 ,
         \SubCellInst_LFInst_14_LFInst_1_n14 ,
         \SubCellInst_LFInst_14_LFInst_1_n13 ,
         \SubCellInst_LFInst_14_LFInst_1_n12 ,
         \SubCellInst_LFInst_14_LFInst_1_n11 ,
         \SubCellInst_LFInst_14_LFInst_1_n10 ,
         \SubCellInst_LFInst_14_LFInst_2_n22 ,
         \SubCellInst_LFInst_14_LFInst_2_n21 ,
         \SubCellInst_LFInst_14_LFInst_2_n20 ,
         \SubCellInst_LFInst_14_LFInst_2_n19 ,
         \SubCellInst_LFInst_14_LFInst_2_n18 ,
         \SubCellInst_LFInst_14_LFInst_2_n17 ,
         \SubCellInst_LFInst_14_LFInst_2_n16 ,
         \SubCellInst_LFInst_14_LFInst_2_n15 ,
         \SubCellInst_LFInst_14_LFInst_3_n16 ,
         \SubCellInst_LFInst_14_LFInst_3_n15 ,
         \SubCellInst_LFInst_14_LFInst_3_n14 ,
         \SubCellInst_LFInst_14_LFInst_3_n13 ,
         \SubCellInst_LFInst_14_LFInst_3_n12 ,
         \SubCellInst_LFInst_14_LFInst_3_n11 ,
         \SubCellInst_LFInst_15_LFInst_0_n10 ,
         \SubCellInst_LFInst_15_LFInst_0_n9 ,
         \SubCellInst_LFInst_15_LFInst_0_n8 ,
         \SubCellInst_LFInst_15_LFInst_0_n7 ,
         \SubCellInst_LFInst_15_LFInst_1_n18 ,
         \SubCellInst_LFInst_15_LFInst_1_n17 ,
         \SubCellInst_LFInst_15_LFInst_1_n16 ,
         \SubCellInst_LFInst_15_LFInst_1_n15 ,
         \SubCellInst_LFInst_15_LFInst_1_n14 ,
         \SubCellInst_LFInst_15_LFInst_1_n13 ,
         \SubCellInst_LFInst_15_LFInst_1_n12 ,
         \SubCellInst_LFInst_15_LFInst_1_n11 ,
         \SubCellInst_LFInst_15_LFInst_1_n10 ,
         \SubCellInst_LFInst_15_LFInst_2_n22 ,
         \SubCellInst_LFInst_15_LFInst_2_n21 ,
         \SubCellInst_LFInst_15_LFInst_2_n20 ,
         \SubCellInst_LFInst_15_LFInst_2_n19 ,
         \SubCellInst_LFInst_15_LFInst_2_n18 ,
         \SubCellInst_LFInst_15_LFInst_2_n17 ,
         \SubCellInst_LFInst_15_LFInst_2_n16 ,
         \SubCellInst_LFInst_15_LFInst_2_n15 ,
         \SubCellInst_LFInst_15_LFInst_3_n16 ,
         \SubCellInst_LFInst_15_LFInst_3_n15 ,
         \SubCellInst_LFInst_15_LFInst_3_n14 ,
         \SubCellInst_LFInst_15_LFInst_3_n13 ,
         \SubCellInst_LFInst_15_LFInst_3_n12 ,
         \SubCellInst_LFInst_15_LFInst_3_n11 , \MCInst_MC0_v0_2Inst_0_n2 ,
         \MCInst_MC0_v1_2Inst_0_n2 , \MCInst_MC0_v2_3Inst_0_n4 ,
         \MCInst_MC0_v2_3Inst_0_n3 , \MCInst_MC0_v3_3Inst_0_n2 ,
         \MCInst_MC0_v0_2Inst_1_n2 , \MCInst_MC0_v2_1Inst_1_n2 ,
         \MCInst_MC0_v2_2Inst_1_n4 , \MCInst_MC0_v2_2Inst_1_n3 ,
         \MCInst_MC0_v3_3Inst_1_n2 , \MCInst_MC0_v1_1Inst_2_n2 ,
         \MCInst_MC0_v1_2Inst_2_n2 , \MCInst_MC0_v2_1Inst_2_n2 ,
         \MCInst_MC0_v2_2Inst_2_n2 , \MCInst_MC0_v3_1Inst_2_n2 ,
         \MCInst_MC0_v1_2Inst_3_n4 , \MCInst_MC0_v1_2Inst_3_n3 ,
         \MCInst_MC0_v2_2Inst_3_n2 , \MCInst_MC0_v2_3Inst_3_n2 ,
         \MCInst_MC0_r0Inst_XORInst_0_0_n5 ,
         \MCInst_MC0_r0Inst_XORInst_0_0_n4 ,
         \MCInst_MC0_r0Inst_XORInst_0_1_n5 ,
         \MCInst_MC0_r0Inst_XORInst_0_1_n4 ,
         \MCInst_MC0_r0Inst_XORInst_0_2_n5 ,
         \MCInst_MC0_r0Inst_XORInst_0_2_n4 ,
         \MCInst_MC0_r0Inst_XORInst_0_3_n5 ,
         \MCInst_MC0_r0Inst_XORInst_0_3_n4 ,
         \MCInst_MC0_r1Inst_XORInst_0_0_n5 ,
         \MCInst_MC0_r1Inst_XORInst_0_0_n4 ,
         \MCInst_MC0_r1Inst_XORInst_0_1_n5 ,
         \MCInst_MC0_r1Inst_XORInst_0_1_n4 ,
         \MCInst_MC0_r1Inst_XORInst_0_2_n5 ,
         \MCInst_MC0_r1Inst_XORInst_0_2_n4 ,
         \MCInst_MC0_r1Inst_XORInst_0_3_n5 ,
         \MCInst_MC0_r1Inst_XORInst_0_3_n4 ,
         \MCInst_MC0_r2Inst_XORInst_0_0_n5 ,
         \MCInst_MC0_r2Inst_XORInst_0_0_n4 ,
         \MCInst_MC0_r2Inst_XORInst_0_1_n5 ,
         \MCInst_MC0_r2Inst_XORInst_0_1_n4 ,
         \MCInst_MC0_r2Inst_XORInst_0_2_n5 ,
         \MCInst_MC0_r2Inst_XORInst_0_2_n4 ,
         \MCInst_MC0_r2Inst_XORInst_0_3_n5 ,
         \MCInst_MC0_r2Inst_XORInst_0_3_n4 ,
         \MCInst_MC0_r3Inst_XORInst_0_0_n5 ,
         \MCInst_MC0_r3Inst_XORInst_0_0_n4 ,
         \MCInst_MC0_r3Inst_XORInst_0_1_n5 ,
         \MCInst_MC0_r3Inst_XORInst_0_1_n4 ,
         \MCInst_MC0_r3Inst_XORInst_0_2_n5 ,
         \MCInst_MC0_r3Inst_XORInst_0_2_n4 ,
         \MCInst_MC0_r3Inst_XORInst_0_3_n5 ,
         \MCInst_MC0_r3Inst_XORInst_0_3_n4 , \MCInst_MC1_v0_2Inst_0_n2 ,
         \MCInst_MC1_v1_2Inst_0_n2 , \MCInst_MC1_v2_3Inst_0_n4 ,
         \MCInst_MC1_v2_3Inst_0_n3 , \MCInst_MC1_v3_3Inst_0_n2 ,
         \MCInst_MC1_v0_2Inst_1_n2 , \MCInst_MC1_v2_1Inst_1_n2 ,
         \MCInst_MC1_v2_2Inst_1_n4 , \MCInst_MC1_v2_2Inst_1_n3 ,
         \MCInst_MC1_v3_3Inst_1_n2 , \MCInst_MC1_v1_1Inst_2_n2 ,
         \MCInst_MC1_v1_2Inst_2_n2 , \MCInst_MC1_v2_1Inst_2_n2 ,
         \MCInst_MC1_v2_2Inst_2_n2 , \MCInst_MC1_v3_1Inst_2_n2 ,
         \MCInst_MC1_v1_2Inst_3_n4 , \MCInst_MC1_v1_2Inst_3_n3 ,
         \MCInst_MC1_v2_2Inst_3_n2 , \MCInst_MC1_v2_3Inst_3_n2 ,
         \MCInst_MC1_r0Inst_XORInst_0_0_n5 ,
         \MCInst_MC1_r0Inst_XORInst_0_0_n4 ,
         \MCInst_MC1_r0Inst_XORInst_0_1_n5 ,
         \MCInst_MC1_r0Inst_XORInst_0_1_n4 ,
         \MCInst_MC1_r0Inst_XORInst_0_2_n5 ,
         \MCInst_MC1_r0Inst_XORInst_0_2_n4 ,
         \MCInst_MC1_r0Inst_XORInst_0_3_n5 ,
         \MCInst_MC1_r0Inst_XORInst_0_3_n4 ,
         \MCInst_MC1_r1Inst_XORInst_0_0_n5 ,
         \MCInst_MC1_r1Inst_XORInst_0_0_n4 ,
         \MCInst_MC1_r1Inst_XORInst_0_1_n5 ,
         \MCInst_MC1_r1Inst_XORInst_0_1_n4 ,
         \MCInst_MC1_r1Inst_XORInst_0_2_n5 ,
         \MCInst_MC1_r1Inst_XORInst_0_2_n4 ,
         \MCInst_MC1_r1Inst_XORInst_0_3_n5 ,
         \MCInst_MC1_r1Inst_XORInst_0_3_n4 ,
         \MCInst_MC1_r2Inst_XORInst_0_0_n5 ,
         \MCInst_MC1_r2Inst_XORInst_0_0_n4 ,
         \MCInst_MC1_r2Inst_XORInst_0_1_n5 ,
         \MCInst_MC1_r2Inst_XORInst_0_1_n4 ,
         \MCInst_MC1_r2Inst_XORInst_0_2_n5 ,
         \MCInst_MC1_r2Inst_XORInst_0_2_n4 ,
         \MCInst_MC1_r2Inst_XORInst_0_3_n5 ,
         \MCInst_MC1_r2Inst_XORInst_0_3_n4 ,
         \MCInst_MC1_r3Inst_XORInst_0_0_n5 ,
         \MCInst_MC1_r3Inst_XORInst_0_0_n4 ,
         \MCInst_MC1_r3Inst_XORInst_0_1_n5 ,
         \MCInst_MC1_r3Inst_XORInst_0_1_n4 ,
         \MCInst_MC1_r3Inst_XORInst_0_2_n5 ,
         \MCInst_MC1_r3Inst_XORInst_0_2_n4 ,
         \MCInst_MC1_r3Inst_XORInst_0_3_n5 ,
         \MCInst_MC1_r3Inst_XORInst_0_3_n4 , \MCInst_MC2_v0_2Inst_0_n2 ,
         \MCInst_MC2_v1_2Inst_0_n2 , \MCInst_MC2_v2_3Inst_0_n4 ,
         \MCInst_MC2_v2_3Inst_0_n3 , \MCInst_MC2_v3_3Inst_0_n2 ,
         \MCInst_MC2_v0_2Inst_1_n2 , \MCInst_MC2_v2_1Inst_1_n2 ,
         \MCInst_MC2_v2_2Inst_1_n4 , \MCInst_MC2_v2_2Inst_1_n3 ,
         \MCInst_MC2_v3_3Inst_1_n2 , \MCInst_MC2_v1_1Inst_2_n2 ,
         \MCInst_MC2_v1_2Inst_2_n2 , \MCInst_MC2_v2_1Inst_2_n2 ,
         \MCInst_MC2_v2_2Inst_2_n2 , \MCInst_MC2_v3_1Inst_2_n2 ,
         \MCInst_MC2_v1_2Inst_3_n4 , \MCInst_MC2_v1_2Inst_3_n3 ,
         \MCInst_MC2_v2_2Inst_3_n2 , \MCInst_MC2_v2_3Inst_3_n2 ,
         \MCInst_MC2_r0Inst_XORInst_0_0_n5 ,
         \MCInst_MC2_r0Inst_XORInst_0_0_n4 ,
         \MCInst_MC2_r0Inst_XORInst_0_1_n5 ,
         \MCInst_MC2_r0Inst_XORInst_0_1_n4 ,
         \MCInst_MC2_r0Inst_XORInst_0_2_n5 ,
         \MCInst_MC2_r0Inst_XORInst_0_2_n4 ,
         \MCInst_MC2_r0Inst_XORInst_0_3_n5 ,
         \MCInst_MC2_r0Inst_XORInst_0_3_n4 ,
         \MCInst_MC2_r1Inst_XORInst_0_0_n5 ,
         \MCInst_MC2_r1Inst_XORInst_0_0_n4 ,
         \MCInst_MC2_r1Inst_XORInst_0_1_n5 ,
         \MCInst_MC2_r1Inst_XORInst_0_1_n4 ,
         \MCInst_MC2_r1Inst_XORInst_0_2_n5 ,
         \MCInst_MC2_r1Inst_XORInst_0_2_n4 ,
         \MCInst_MC2_r1Inst_XORInst_0_3_n5 ,
         \MCInst_MC2_r1Inst_XORInst_0_3_n4 ,
         \MCInst_MC2_r2Inst_XORInst_0_0_n5 ,
         \MCInst_MC2_r2Inst_XORInst_0_0_n4 ,
         \MCInst_MC2_r2Inst_XORInst_0_1_n5 ,
         \MCInst_MC2_r2Inst_XORInst_0_1_n4 ,
         \MCInst_MC2_r2Inst_XORInst_0_2_n5 ,
         \MCInst_MC2_r2Inst_XORInst_0_2_n4 ,
         \MCInst_MC2_r2Inst_XORInst_0_3_n5 ,
         \MCInst_MC2_r2Inst_XORInst_0_3_n4 ,
         \MCInst_MC2_r3Inst_XORInst_0_0_n5 ,
         \MCInst_MC2_r3Inst_XORInst_0_0_n4 ,
         \MCInst_MC2_r3Inst_XORInst_0_1_n5 ,
         \MCInst_MC2_r3Inst_XORInst_0_1_n4 ,
         \MCInst_MC2_r3Inst_XORInst_0_2_n5 ,
         \MCInst_MC2_r3Inst_XORInst_0_2_n4 ,
         \MCInst_MC2_r3Inst_XORInst_0_3_n5 ,
         \MCInst_MC2_r3Inst_XORInst_0_3_n4 , \MCInst_MC3_v0_2Inst_0_n2 ,
         \MCInst_MC3_v1_2Inst_0_n2 , \MCInst_MC3_v2_3Inst_0_n4 ,
         \MCInst_MC3_v2_3Inst_0_n3 , \MCInst_MC3_v3_3Inst_0_n2 ,
         \MCInst_MC3_v0_2Inst_1_n2 , \MCInst_MC3_v2_1Inst_1_n2 ,
         \MCInst_MC3_v2_2Inst_1_n4 , \MCInst_MC3_v2_2Inst_1_n3 ,
         \MCInst_MC3_v3_3Inst_1_n2 , \MCInst_MC3_v1_1Inst_2_n2 ,
         \MCInst_MC3_v1_2Inst_2_n2 , \MCInst_MC3_v2_1Inst_2_n2 ,
         \MCInst_MC3_v2_2Inst_2_n2 , \MCInst_MC3_v3_1Inst_2_n2 ,
         \MCInst_MC3_v1_2Inst_3_n4 , \MCInst_MC3_v1_2Inst_3_n3 ,
         \MCInst_MC3_v2_2Inst_3_n2 , \MCInst_MC3_v2_3Inst_3_n2 ,
         \MCInst_MC3_r0Inst_XORInst_0_0_n5 ,
         \MCInst_MC3_r0Inst_XORInst_0_0_n4 ,
         \MCInst_MC3_r0Inst_XORInst_0_1_n5 ,
         \MCInst_MC3_r0Inst_XORInst_0_1_n4 ,
         \MCInst_MC3_r0Inst_XORInst_0_2_n5 ,
         \MCInst_MC3_r0Inst_XORInst_0_2_n4 ,
         \MCInst_MC3_r0Inst_XORInst_0_3_n5 ,
         \MCInst_MC3_r0Inst_XORInst_0_3_n4 ,
         \MCInst_MC3_r1Inst_XORInst_0_0_n5 ,
         \MCInst_MC3_r1Inst_XORInst_0_0_n4 ,
         \MCInst_MC3_r1Inst_XORInst_0_1_n5 ,
         \MCInst_MC3_r1Inst_XORInst_0_1_n4 ,
         \MCInst_MC3_r1Inst_XORInst_0_2_n5 ,
         \MCInst_MC3_r1Inst_XORInst_0_2_n4 ,
         \MCInst_MC3_r1Inst_XORInst_0_3_n5 ,
         \MCInst_MC3_r1Inst_XORInst_0_3_n4 ,
         \MCInst_MC3_r2Inst_XORInst_0_0_n5 ,
         \MCInst_MC3_r2Inst_XORInst_0_0_n4 ,
         \MCInst_MC3_r2Inst_XORInst_0_1_n5 ,
         \MCInst_MC3_r2Inst_XORInst_0_1_n4 ,
         \MCInst_MC3_r2Inst_XORInst_0_2_n5 ,
         \MCInst_MC3_r2Inst_XORInst_0_2_n4 ,
         \MCInst_MC3_r2Inst_XORInst_0_3_n5 ,
         \MCInst_MC3_r2Inst_XORInst_0_3_n4 ,
         \MCInst_MC3_r3Inst_XORInst_0_0_n5 ,
         \MCInst_MC3_r3Inst_XORInst_0_0_n4 ,
         \MCInst_MC3_r3Inst_XORInst_0_1_n5 ,
         \MCInst_MC3_r3Inst_XORInst_0_1_n4 ,
         \MCInst_MC3_r3Inst_XORInst_0_2_n5 ,
         \MCInst_MC3_r3Inst_XORInst_0_2_n4 ,
         \MCInst_MC3_r3Inst_XORInst_0_3_n5 ,
         \MCInst_MC3_r3Inst_XORInst_0_3_n4 ,
         \Red_PlaintextInst_LFInst_0_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_0_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_0_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_1_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_1_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_1_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_2_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_2_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_2_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_3_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_3_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_3_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_4_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_4_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_4_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_5_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_5_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_5_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_6_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_6_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_6_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_7_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_7_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_7_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_8_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_8_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_8_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_9_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_9_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_9_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_10_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_10_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_10_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_11_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_11_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_11_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_12_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_12_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_12_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_13_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_13_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_13_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_14_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_14_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_14_LFInst_2_n2 ,
         \Red_PlaintextInst_LFInst_15_LFInst_0_n2 ,
         \Red_PlaintextInst_LFInst_15_LFInst_1_n2 ,
         \Red_PlaintextInst_LFInst_15_LFInst_2_n2 ,
         \Red_MCInst_MC0_v1_0Inst_0_n2 , \Red_MCInst_MC0_v2_2Inst_0_n2 ,
         \Red_MCInst_MC0_v2_3Inst_0_n2 , \Red_MCInst_MC0_v3_2Inst_0_n4 ,
         \Red_MCInst_MC0_v3_2Inst_0_n3 , \Red_MCInst_MC0_v0_1Inst_1_n2 ,
         \Red_MCInst_MC0_v1_0Inst_1_n2 , \Red_MCInst_MC0_v1_1Inst_1_n4 ,
         \Red_MCInst_MC0_v1_1Inst_1_n3 , \Red_MCInst_MC0_v3_1Inst_1_n4 ,
         \Red_MCInst_MC0_v3_1Inst_1_n3 , \Red_MCInst_MC0_v0_0Inst_2_n2 ,
         \Red_MCInst_MC0_v0_3Inst_2_n4 , \Red_MCInst_MC0_v0_3Inst_2_n3 ,
         \Red_MCInst_MC0_v1_0Inst_2_n2 , \Red_MCInst_MC0_v1_2Inst_2_n2 ,
         \Red_MCInst_MC0_v1_3Inst_2_n4 , \Red_MCInst_MC0_v1_3Inst_2_n3 ,
         \Red_MCInst_MC0_v2_0Inst_2_n4 , \Red_MCInst_MC0_v2_0Inst_2_n3 ,
         \Red_MCInst_MC0_v3_0Inst_2_n4 , \Red_MCInst_MC0_v3_0Inst_2_n3 ,
         \Red_MCInst_MC0_v3_2Inst_2_n2 ,
         \Red_MCInst_MC0_r0Inst_XORInst_0_0_n5 ,
         \Red_MCInst_MC0_r0Inst_XORInst_0_0_n4 ,
         \Red_MCInst_MC0_r0Inst_XORInst_0_1_n5 ,
         \Red_MCInst_MC0_r0Inst_XORInst_0_1_n4 ,
         \Red_MCInst_MC0_r0Inst_XORInst_0_2_n5 ,
         \Red_MCInst_MC0_r0Inst_XORInst_0_2_n4 ,
         \Red_MCInst_MC0_r1Inst_XORInst_0_0_n5 ,
         \Red_MCInst_MC0_r1Inst_XORInst_0_0_n4 ,
         \Red_MCInst_MC0_r1Inst_XORInst_0_1_n5 ,
         \Red_MCInst_MC0_r1Inst_XORInst_0_1_n4 ,
         \Red_MCInst_MC0_r1Inst_XORInst_0_2_n5 ,
         \Red_MCInst_MC0_r1Inst_XORInst_0_2_n4 ,
         \Red_MCInst_MC0_r2Inst_XORInst_0_0_n5 ,
         \Red_MCInst_MC0_r2Inst_XORInst_0_0_n4 ,
         \Red_MCInst_MC0_r2Inst_XORInst_0_1_n5 ,
         \Red_MCInst_MC0_r2Inst_XORInst_0_1_n4 ,
         \Red_MCInst_MC0_r2Inst_XORInst_0_2_n5 ,
         \Red_MCInst_MC0_r2Inst_XORInst_0_2_n4 ,
         \Red_MCInst_MC0_r3Inst_XORInst_0_0_n5 ,
         \Red_MCInst_MC0_r3Inst_XORInst_0_0_n4 ,
         \Red_MCInst_MC0_r3Inst_XORInst_0_1_n5 ,
         \Red_MCInst_MC0_r3Inst_XORInst_0_1_n4 ,
         \Red_MCInst_MC0_r3Inst_XORInst_0_2_n5 ,
         \Red_MCInst_MC0_r3Inst_XORInst_0_2_n4 ,
         \Red_MCInst_MC1_v1_0Inst_0_n2 , \Red_MCInst_MC1_v2_2Inst_0_n2 ,
         \Red_MCInst_MC1_v2_3Inst_0_n2 , \Red_MCInst_MC1_v3_2Inst_0_n4 ,
         \Red_MCInst_MC1_v3_2Inst_0_n3 , \Red_MCInst_MC1_v0_1Inst_1_n2 ,
         \Red_MCInst_MC1_v1_0Inst_1_n2 , \Red_MCInst_MC1_v1_1Inst_1_n4 ,
         \Red_MCInst_MC1_v1_1Inst_1_n3 , \Red_MCInst_MC1_v3_1Inst_1_n4 ,
         \Red_MCInst_MC1_v3_1Inst_1_n3 , \Red_MCInst_MC1_v0_0Inst_2_n2 ,
         \Red_MCInst_MC1_v0_3Inst_2_n4 , \Red_MCInst_MC1_v0_3Inst_2_n3 ,
         \Red_MCInst_MC1_v1_0Inst_2_n2 , \Red_MCInst_MC1_v1_2Inst_2_n2 ,
         \Red_MCInst_MC1_v1_3Inst_2_n4 , \Red_MCInst_MC1_v1_3Inst_2_n3 ,
         \Red_MCInst_MC1_v2_0Inst_2_n4 , \Red_MCInst_MC1_v2_0Inst_2_n3 ,
         \Red_MCInst_MC1_v3_0Inst_2_n4 , \Red_MCInst_MC1_v3_0Inst_2_n3 ,
         \Red_MCInst_MC1_v3_2Inst_2_n2 ,
         \Red_MCInst_MC1_r0Inst_XORInst_0_0_n5 ,
         \Red_MCInst_MC1_r0Inst_XORInst_0_0_n4 ,
         \Red_MCInst_MC1_r0Inst_XORInst_0_1_n5 ,
         \Red_MCInst_MC1_r0Inst_XORInst_0_1_n4 ,
         \Red_MCInst_MC1_r0Inst_XORInst_0_2_n5 ,
         \Red_MCInst_MC1_r0Inst_XORInst_0_2_n4 ,
         \Red_MCInst_MC1_r1Inst_XORInst_0_0_n5 ,
         \Red_MCInst_MC1_r1Inst_XORInst_0_0_n4 ,
         \Red_MCInst_MC1_r1Inst_XORInst_0_1_n5 ,
         \Red_MCInst_MC1_r1Inst_XORInst_0_1_n4 ,
         \Red_MCInst_MC1_r1Inst_XORInst_0_2_n5 ,
         \Red_MCInst_MC1_r1Inst_XORInst_0_2_n4 ,
         \Red_MCInst_MC1_r2Inst_XORInst_0_0_n5 ,
         \Red_MCInst_MC1_r2Inst_XORInst_0_0_n4 ,
         \Red_MCInst_MC1_r2Inst_XORInst_0_1_n5 ,
         \Red_MCInst_MC1_r2Inst_XORInst_0_1_n4 ,
         \Red_MCInst_MC1_r2Inst_XORInst_0_2_n5 ,
         \Red_MCInst_MC1_r2Inst_XORInst_0_2_n4 ,
         \Red_MCInst_MC1_r3Inst_XORInst_0_0_n5 ,
         \Red_MCInst_MC1_r3Inst_XORInst_0_0_n4 ,
         \Red_MCInst_MC1_r3Inst_XORInst_0_1_n5 ,
         \Red_MCInst_MC1_r3Inst_XORInst_0_1_n4 ,
         \Red_MCInst_MC1_r3Inst_XORInst_0_2_n5 ,
         \Red_MCInst_MC1_r3Inst_XORInst_0_2_n4 ,
         \Red_MCInst_MC2_v1_0Inst_0_n2 , \Red_MCInst_MC2_v2_2Inst_0_n2 ,
         \Red_MCInst_MC2_v2_3Inst_0_n2 , \Red_MCInst_MC2_v3_2Inst_0_n4 ,
         \Red_MCInst_MC2_v3_2Inst_0_n3 , \Red_MCInst_MC2_v0_1Inst_1_n2 ,
         \Red_MCInst_MC2_v1_0Inst_1_n2 , \Red_MCInst_MC2_v1_1Inst_1_n4 ,
         \Red_MCInst_MC2_v1_1Inst_1_n3 , \Red_MCInst_MC2_v3_1Inst_1_n4 ,
         \Red_MCInst_MC2_v3_1Inst_1_n3 , \Red_MCInst_MC2_v0_0Inst_2_n2 ,
         \Red_MCInst_MC2_v0_3Inst_2_n4 , \Red_MCInst_MC2_v0_3Inst_2_n3 ,
         \Red_MCInst_MC2_v1_0Inst_2_n2 , \Red_MCInst_MC2_v1_2Inst_2_n2 ,
         \Red_MCInst_MC2_v1_3Inst_2_n4 , \Red_MCInst_MC2_v1_3Inst_2_n3 ,
         \Red_MCInst_MC2_v2_0Inst_2_n4 , \Red_MCInst_MC2_v2_0Inst_2_n3 ,
         \Red_MCInst_MC2_v3_0Inst_2_n4 , \Red_MCInst_MC2_v3_0Inst_2_n3 ,
         \Red_MCInst_MC2_v3_2Inst_2_n2 ,
         \Red_MCInst_MC2_r0Inst_XORInst_0_0_n5 ,
         \Red_MCInst_MC2_r0Inst_XORInst_0_0_n4 ,
         \Red_MCInst_MC2_r0Inst_XORInst_0_1_n5 ,
         \Red_MCInst_MC2_r0Inst_XORInst_0_1_n4 ,
         \Red_MCInst_MC2_r0Inst_XORInst_0_2_n5 ,
         \Red_MCInst_MC2_r0Inst_XORInst_0_2_n4 ,
         \Red_MCInst_MC2_r1Inst_XORInst_0_0_n5 ,
         \Red_MCInst_MC2_r1Inst_XORInst_0_0_n4 ,
         \Red_MCInst_MC2_r1Inst_XORInst_0_1_n5 ,
         \Red_MCInst_MC2_r1Inst_XORInst_0_1_n4 ,
         \Red_MCInst_MC2_r1Inst_XORInst_0_2_n5 ,
         \Red_MCInst_MC2_r1Inst_XORInst_0_2_n4 ,
         \Red_MCInst_MC2_r2Inst_XORInst_0_0_n5 ,
         \Red_MCInst_MC2_r2Inst_XORInst_0_0_n4 ,
         \Red_MCInst_MC2_r2Inst_XORInst_0_1_n5 ,
         \Red_MCInst_MC2_r2Inst_XORInst_0_1_n4 ,
         \Red_MCInst_MC2_r2Inst_XORInst_0_2_n5 ,
         \Red_MCInst_MC2_r2Inst_XORInst_0_2_n4 ,
         \Red_MCInst_MC2_r3Inst_XORInst_0_0_n5 ,
         \Red_MCInst_MC2_r3Inst_XORInst_0_0_n4 ,
         \Red_MCInst_MC2_r3Inst_XORInst_0_1_n5 ,
         \Red_MCInst_MC2_r3Inst_XORInst_0_1_n4 ,
         \Red_MCInst_MC2_r3Inst_XORInst_0_2_n5 ,
         \Red_MCInst_MC2_r3Inst_XORInst_0_2_n4 ,
         \Red_MCInst_MC3_v1_0Inst_0_n2 , \Red_MCInst_MC3_v2_2Inst_0_n2 ,
         \Red_MCInst_MC3_v2_3Inst_0_n2 , \Red_MCInst_MC3_v3_2Inst_0_n4 ,
         \Red_MCInst_MC3_v3_2Inst_0_n3 , \Red_MCInst_MC3_v0_1Inst_1_n2 ,
         \Red_MCInst_MC3_v1_0Inst_1_n2 , \Red_MCInst_MC3_v1_1Inst_1_n4 ,
         \Red_MCInst_MC3_v1_1Inst_1_n3 , \Red_MCInst_MC3_v3_1Inst_1_n4 ,
         \Red_MCInst_MC3_v3_1Inst_1_n3 , \Red_MCInst_MC3_v0_0Inst_2_n2 ,
         \Red_MCInst_MC3_v0_3Inst_2_n4 , \Red_MCInst_MC3_v0_3Inst_2_n3 ,
         \Red_MCInst_MC3_v1_0Inst_2_n2 , \Red_MCInst_MC3_v1_2Inst_2_n2 ,
         \Red_MCInst_MC3_v1_3Inst_2_n4 , \Red_MCInst_MC3_v1_3Inst_2_n3 ,
         \Red_MCInst_MC3_v2_0Inst_2_n4 , \Red_MCInst_MC3_v2_0Inst_2_n3 ,
         \Red_MCInst_MC3_v3_0Inst_2_n4 , \Red_MCInst_MC3_v3_0Inst_2_n3 ,
         \Red_MCInst_MC3_v3_2Inst_2_n2 ,
         \Red_MCInst_MC3_r0Inst_XORInst_0_0_n5 ,
         \Red_MCInst_MC3_r0Inst_XORInst_0_0_n4 ,
         \Red_MCInst_MC3_r0Inst_XORInst_0_1_n5 ,
         \Red_MCInst_MC3_r0Inst_XORInst_0_1_n4 ,
         \Red_MCInst_MC3_r0Inst_XORInst_0_2_n5 ,
         \Red_MCInst_MC3_r0Inst_XORInst_0_2_n4 ,
         \Red_MCInst_MC3_r1Inst_XORInst_0_0_n5 ,
         \Red_MCInst_MC3_r1Inst_XORInst_0_0_n4 ,
         \Red_MCInst_MC3_r1Inst_XORInst_0_1_n5 ,
         \Red_MCInst_MC3_r1Inst_XORInst_0_1_n4 ,
         \Red_MCInst_MC3_r1Inst_XORInst_0_2_n5 ,
         \Red_MCInst_MC3_r1Inst_XORInst_0_2_n4 ,
         \Red_MCInst_MC3_r2Inst_XORInst_0_0_n5 ,
         \Red_MCInst_MC3_r2Inst_XORInst_0_0_n4 ,
         \Red_MCInst_MC3_r2Inst_XORInst_0_1_n5 ,
         \Red_MCInst_MC3_r2Inst_XORInst_0_1_n4 ,
         \Red_MCInst_MC3_r2Inst_XORInst_0_2_n5 ,
         \Red_MCInst_MC3_r2Inst_XORInst_0_2_n4 ,
         \Red_MCInst_MC3_r3Inst_XORInst_0_0_n5 ,
         \Red_MCInst_MC3_r3Inst_XORInst_0_0_n4 ,
         \Red_MCInst_MC3_r3Inst_XORInst_0_1_n5 ,
         \Red_MCInst_MC3_r3Inst_XORInst_0_1_n4 ,
         \Red_MCInst_MC3_r3Inst_XORInst_0_2_n5 ,
         \Red_MCInst_MC3_r3Inst_XORInst_0_2_n4 ,
         \Red_KeyInst_LFInst_0_LFInst_0_n2 ,
         \Red_KeyInst_LFInst_0_LFInst_1_n2 ,
         \Red_KeyInst_LFInst_0_LFInst_2_n2 ,
         \Red_KeyInst_LFInst_1_LFInst_0_n2 ,
         \Red_KeyInst_LFInst_1_LFInst_1_n2 ,
         \Red_KeyInst_LFInst_1_LFInst_2_n2 ,
         \Red_KeyInst_LFInst_2_LFInst_0_n2 ,
         \Red_KeyInst_LFInst_2_LFInst_1_n2 ,
         \Red_KeyInst_LFInst_2_LFInst_2_n2 ,
         \Red_KeyInst_LFInst_3_LFInst_0_n2 ,
         \Red_KeyInst_LFInst_3_LFInst_1_n2 ,
         \Red_KeyInst_LFInst_3_LFInst_2_n2 ,
         \Red_KeyInst_LFInst_4_LFInst_0_n2 ,
         \Red_KeyInst_LFInst_4_LFInst_1_n2 ,
         \Red_KeyInst_LFInst_4_LFInst_2_n2 ,
         \Red_KeyInst_LFInst_5_LFInst_0_n2 ,
         \Red_KeyInst_LFInst_5_LFInst_1_n2 ,
         \Red_KeyInst_LFInst_5_LFInst_2_n2 ,
         \Red_KeyInst_LFInst_6_LFInst_0_n2 ,
         \Red_KeyInst_LFInst_6_LFInst_1_n2 ,
         \Red_KeyInst_LFInst_6_LFInst_2_n2 ,
         \Red_KeyInst_LFInst_7_LFInst_0_n2 ,
         \Red_KeyInst_LFInst_7_LFInst_1_n2 ,
         \Red_KeyInst_LFInst_7_LFInst_2_n2 ,
         \Red_KeyInst_LFInst_8_LFInst_0_n2 ,
         \Red_KeyInst_LFInst_8_LFInst_1_n2 ,
         \Red_KeyInst_LFInst_8_LFInst_2_n2 ,
         \Red_KeyInst_LFInst_9_LFInst_0_n2 ,
         \Red_KeyInst_LFInst_9_LFInst_1_n2 ,
         \Red_KeyInst_LFInst_9_LFInst_2_n2 ,
         \Red_KeyInst_LFInst_10_LFInst_0_n2 ,
         \Red_KeyInst_LFInst_10_LFInst_1_n2 ,
         \Red_KeyInst_LFInst_10_LFInst_2_n2 ,
         \Red_KeyInst_LFInst_11_LFInst_0_n2 ,
         \Red_KeyInst_LFInst_11_LFInst_1_n2 ,
         \Red_KeyInst_LFInst_11_LFInst_2_n2 ,
         \Red_KeyInst_LFInst_12_LFInst_0_n2 ,
         \Red_KeyInst_LFInst_12_LFInst_1_n2 ,
         \Red_KeyInst_LFInst_12_LFInst_2_n2 ,
         \Red_KeyInst_LFInst_13_LFInst_0_n2 ,
         \Red_KeyInst_LFInst_13_LFInst_1_n2 ,
         \Red_KeyInst_LFInst_13_LFInst_2_n2 ,
         \Red_KeyInst_LFInst_14_LFInst_0_n2 ,
         \Red_KeyInst_LFInst_14_LFInst_1_n2 ,
         \Red_KeyInst_LFInst_14_LFInst_2_n2 ,
         \Red_KeyInst_LFInst_15_LFInst_0_n2 ,
         \Red_KeyInst_LFInst_15_LFInst_1_n2 ,
         \Red_KeyInst_LFInst_15_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_0_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_0_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_0_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_1_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_1_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_1_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_2_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_2_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_2_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_3_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_3_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_3_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_4_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_4_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_4_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_5_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_5_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_5_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_6_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_6_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_6_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_7_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_7_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_7_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_8_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_8_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_8_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_9_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_9_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_9_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_10_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_10_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_10_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_11_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_11_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_11_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_12_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_12_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_12_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_13_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_13_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_13_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_14_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_14_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_14_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_15_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_15_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_15_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_16_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_16_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_16_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_17_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_17_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_17_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_18_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_18_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_18_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_19_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_19_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_19_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_20_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_20_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_20_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_21_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_21_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_21_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_22_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_22_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_22_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_23_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_23_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_23_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_24_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_24_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_24_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_25_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_25_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_25_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_26_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_26_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_26_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_27_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_27_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_27_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_28_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_28_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_28_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_29_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_29_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_29_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_30_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_30_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_30_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_31_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_31_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_31_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_32_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_32_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_32_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_33_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_33_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_33_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_34_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_34_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_34_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_35_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_35_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_35_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_36_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_36_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_36_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_37_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_37_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_37_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_38_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_38_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_38_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_39_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_39_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_39_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_40_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_40_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_40_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_41_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_41_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_41_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_42_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_42_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_42_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_43_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_43_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_43_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_44_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_44_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_44_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_45_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_45_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_45_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_46_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_46_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_46_LFInst_2_n2 ,
         \Red_ToCheckInst_LFInst_47_LFInst_0_n2 ,
         \Red_ToCheckInst_LFInst_47_LFInst_1_n2 ,
         \Red_ToCheckInst_LFInst_47_LFInst_2_n2 , \Check1_CheckInst_0_n95 ,
         \Check1_CheckInst_0_n94 , \Check1_CheckInst_0_n93 ,
         \Check1_CheckInst_0_n92 , \Check1_CheckInst_0_n91 ,
         \Check1_CheckInst_0_n90 , \Check1_CheckInst_0_n89 ,
         \Check1_CheckInst_0_n88 , \Check1_CheckInst_0_n87 ,
         \Check1_CheckInst_0_n86 , \Check1_CheckInst_0_n85 ,
         \Check1_CheckInst_0_n84 , \Check1_CheckInst_0_n83 ,
         \Check1_CheckInst_0_n82 , \Check1_CheckInst_0_n81 ,
         \Check1_CheckInst_0_n80 , \Check1_CheckInst_0_n79 ,
         \Check1_CheckInst_0_n78 , \Check1_CheckInst_0_n77 ,
         \Check1_CheckInst_0_n76 , \Check1_CheckInst_0_n75 ,
         \Check1_CheckInst_0_n74 , \Check1_CheckInst_0_n73 ,
         \Check1_CheckInst_0_n72 , \Check1_CheckInst_0_n71 ,
         \Check1_CheckInst_0_n70 , \Check1_CheckInst_0_n69 ,
         \Check1_CheckInst_0_n68 , \Check1_CheckInst_0_n67 ,
         \Check1_CheckInst_0_n66 , \Check1_CheckInst_0_n65 ,
         \Check1_CheckInst_0_n64 , \Check1_CheckInst_0_n63 ,
         \Check1_CheckInst_0_n62 , \Check1_CheckInst_0_n61 ,
         \Check1_CheckInst_0_n60 , \Check1_CheckInst_0_n59 ,
         \Check1_CheckInst_0_n58 , \Check1_CheckInst_0_n57 ,
         \Check1_CheckInst_0_n56 , \Check1_CheckInst_0_n55 ,
         \Check1_CheckInst_0_n54 , \Check1_CheckInst_0_n53 ,
         \Check1_CheckInst_0_n52 , \Check1_CheckInst_0_n51 ,
         \Check1_CheckInst_0_n50 , \Check1_CheckInst_0_n49 ,
         \Check1_CheckInst_0_n48 , \Check1_CheckInst_0_n47 ,
         \Check1_CheckInst_0_n46 , \Check1_CheckInst_0_n45 ,
         \Check1_CheckInst_0_n44 , \Check1_CheckInst_0_n43 ,
         \Check1_CheckInst_0_n42 , \Check1_CheckInst_0_n41 ,
         \Check1_CheckInst_0_n40 , \Check1_CheckInst_0_n39 ,
         \Check1_CheckInst_0_n38 , \Check1_CheckInst_0_n37 ,
         \Check1_CheckInst_0_n36 , \Check1_CheckInst_0_n35 ,
         \Check1_CheckInst_0_n34 , \Check1_CheckInst_0_n33 ,
         \Check1_CheckInst_0_n32 , \Check1_CheckInst_0_n31 ,
         \Check1_CheckInst_0_n30 , \Check1_CheckInst_0_n29 ,
         \Check1_CheckInst_0_n28 , \Check1_CheckInst_0_n27 ,
         \Check1_CheckInst_0_n26 , \Check1_CheckInst_0_n25 ,
         \Check1_CheckInst_0_n24 , \Check1_CheckInst_0_n23 ,
         \Check1_CheckInst_0_n22 , \Check1_CheckInst_0_n21 ,
         \Check1_CheckInst_0_n20 , \Check1_CheckInst_0_n19 ,
         \Check1_CheckInst_0_n18 , \Check1_CheckInst_1_n96 ,
         \Check1_CheckInst_1_n95 , \Check1_CheckInst_1_n94 ,
         \Check1_CheckInst_1_n93 , \Check1_CheckInst_1_n92 ,
         \Check1_CheckInst_1_n91 , \Check1_CheckInst_1_n90 ,
         \Check1_CheckInst_1_n89 , \Check1_CheckInst_1_n88 ,
         \Check1_CheckInst_1_n87 , \Check1_CheckInst_1_n86 ,
         \Check1_CheckInst_1_n85 , \Check1_CheckInst_1_n84 ,
         \Check1_CheckInst_1_n83 , \Check1_CheckInst_1_n82 ,
         \Check1_CheckInst_1_n81 , \Check1_CheckInst_1_n80 ,
         \Check1_CheckInst_1_n79 , \Check1_CheckInst_1_n78 ,
         \Check1_CheckInst_1_n77 , \Check1_CheckInst_1_n76 ,
         \Check1_CheckInst_1_n75 , \Check1_CheckInst_1_n74 ,
         \Check1_CheckInst_1_n73 , \Check1_CheckInst_1_n72 ,
         \Check1_CheckInst_1_n71 , \Check1_CheckInst_1_n70 ,
         \Check1_CheckInst_1_n69 , \Check1_CheckInst_1_n68 ,
         \Check1_CheckInst_1_n67 , \Check1_CheckInst_1_n66 ,
         \Check1_CheckInst_1_n65 , \Check1_CheckInst_1_n64 ,
         \Check1_CheckInst_1_n63 , \Check1_CheckInst_1_n62 ,
         \Check1_CheckInst_1_n61 , \Check1_CheckInst_1_n60 ,
         \Check1_CheckInst_1_n59 , \Check1_CheckInst_1_n58 ,
         \Check1_CheckInst_1_n57 , \Check1_CheckInst_1_n56 ,
         \Check1_CheckInst_1_n55 , \Check1_CheckInst_1_n54 ,
         \Check1_CheckInst_1_n53 , \Check1_CheckInst_1_n52 ,
         \Check1_CheckInst_1_n51 , \Check1_CheckInst_1_n50 ,
         \Check1_CheckInst_1_n49 , \Check1_CheckInst_1_n48 ,
         \Check1_CheckInst_1_n47 , \Check1_CheckInst_1_n46 ,
         \Check1_CheckInst_1_n45 , \Check1_CheckInst_1_n44 ,
         \Check1_CheckInst_1_n43 , \Check1_CheckInst_1_n42 ,
         \Check1_CheckInst_1_n41 , \Check1_CheckInst_1_n40 ,
         \Check1_CheckInst_1_n39 , \Check1_CheckInst_1_n38 ,
         \Check1_CheckInst_1_n37 , \Check1_CheckInst_1_n36 ,
         \Check1_CheckInst_1_n35 , \Check1_CheckInst_1_n34 ,
         \Check1_CheckInst_1_n33 , \Check1_CheckInst_1_n32 ,
         \Check1_CheckInst_1_n31 , \Check1_CheckInst_1_n30 ,
         \Check1_CheckInst_1_n29 , \Check1_CheckInst_1_n28 ,
         \Check1_CheckInst_1_n27 , \Check1_CheckInst_1_n26 ,
         \Check1_CheckInst_1_n25 , \Check1_CheckInst_1_n24 ,
         \Check1_CheckInst_1_n23 , \Check1_CheckInst_1_n22 ,
         \Check1_CheckInst_1_n21 , \Check1_CheckInst_1_n20 ,
         \Check1_CheckInst_1_n19 , \Check1_CheckInst_2_n96 ,
         \Check1_CheckInst_2_n95 , \Check1_CheckInst_2_n94 ,
         \Check1_CheckInst_2_n93 , \Check1_CheckInst_2_n92 ,
         \Check1_CheckInst_2_n91 , \Check1_CheckInst_2_n90 ,
         \Check1_CheckInst_2_n89 , \Check1_CheckInst_2_n88 ,
         \Check1_CheckInst_2_n87 , \Check1_CheckInst_2_n86 ,
         \Check1_CheckInst_2_n85 , \Check1_CheckInst_2_n84 ,
         \Check1_CheckInst_2_n83 , \Check1_CheckInst_2_n82 ,
         \Check1_CheckInst_2_n81 , \Check1_CheckInst_2_n80 ,
         \Check1_CheckInst_2_n79 , \Check1_CheckInst_2_n78 ,
         \Check1_CheckInst_2_n77 , \Check1_CheckInst_2_n76 ,
         \Check1_CheckInst_2_n75 , \Check1_CheckInst_2_n74 ,
         \Check1_CheckInst_2_n73 , \Check1_CheckInst_2_n72 ,
         \Check1_CheckInst_2_n71 , \Check1_CheckInst_2_n70 ,
         \Check1_CheckInst_2_n69 , \Check1_CheckInst_2_n68 ,
         \Check1_CheckInst_2_n67 , \Check1_CheckInst_2_n66 ,
         \Check1_CheckInst_2_n65 , \Check1_CheckInst_2_n64 ,
         \Check1_CheckInst_2_n63 , \Check1_CheckInst_2_n62 ,
         \Check1_CheckInst_2_n61 , \Check1_CheckInst_2_n60 ,
         \Check1_CheckInst_2_n59 , \Check1_CheckInst_2_n58 ,
         \Check1_CheckInst_2_n57 , \Check1_CheckInst_2_n56 ,
         \Check1_CheckInst_2_n55 , \Check1_CheckInst_2_n54 ,
         \Check1_CheckInst_2_n53 , \Check1_CheckInst_2_n52 ,
         \Check1_CheckInst_2_n51 , \Check1_CheckInst_2_n50 ,
         \Check1_CheckInst_2_n49 , \Check1_CheckInst_2_n48 ,
         \Check1_CheckInst_2_n47 , \Check1_CheckInst_2_n46 ,
         \Check1_CheckInst_2_n45 , \Check1_CheckInst_2_n44 ,
         \Check1_CheckInst_2_n43 , \Check1_CheckInst_2_n42 ,
         \Check1_CheckInst_2_n41 , \Check1_CheckInst_2_n40 ,
         \Check1_CheckInst_2_n39 , \Check1_CheckInst_2_n38 ,
         \Check1_CheckInst_2_n37 , \Check1_CheckInst_2_n36 ,
         \Check1_CheckInst_2_n35 , \Check1_CheckInst_2_n34 ,
         \Check1_CheckInst_2_n33 , \Check1_CheckInst_2_n32 ,
         \Check1_CheckInst_2_n31 , \Check1_CheckInst_2_n30 ,
         \Check1_CheckInst_2_n29 , \Check1_CheckInst_2_n28 ,
         \Check1_CheckInst_2_n27 , \Check1_CheckInst_2_n26 ,
         \Check1_CheckInst_2_n25 , \Check1_CheckInst_2_n24 ,
         \Check1_CheckInst_2_n23 , \Check1_CheckInst_2_n22 ,
         \Check1_CheckInst_2_n21 , \Check1_CheckInst_2_n20 ,
         \Check1_CheckInst_2_n19 ;
  wire   [63:0] AddRoundKeyOutput;
  wire   [47:0] Red_Plaintext;
  wire   [47:0] Red_RoundKey;
  wire   [47:0] Red_AddRoundKeyOutput;
  wire   [47:0] Red_Feedback;
  wire   [143:0] Red_SignaltoCheck;
  wire   [2:0] Error;
  wire   [3:0] \MCInst_MC0_v3_3 ;
  wire   [3:0] \MCInst_MC0_v3_2 ;
  wire   [3:0] \MCInst_MC0_v3_1 ;
  wire   [3:0] \MCInst_MC0_v3_0 ;
  wire   [3:0] \MCInst_MC0_v2_3 ;
  wire   [3:0] \MCInst_MC0_v2_2 ;
  wire   [3:0] \MCInst_MC0_v2_1 ;
  wire   [3:0] \MCInst_MC0_v2_0 ;
  wire   [3:0] \MCInst_MC0_v1_3 ;
  wire   [3:0] \MCInst_MC0_v1_2 ;
  wire   [3:0] \MCInst_MC0_v1_1 ;
  wire   [3:0] \MCInst_MC0_v1_0 ;
  wire   [3:0] \MCInst_MC0_v0_3 ;
  wire   [3:0] \MCInst_MC0_v0_2 ;
  wire   [3:0] \MCInst_MC0_v0_1 ;
  wire   [3:0] \MCInst_MC0_v0_0 ;
  wire   [3:0] \MCInst_MC1_v3_3 ;
  wire   [3:0] \MCInst_MC1_v3_2 ;
  wire   [3:0] \MCInst_MC1_v3_1 ;
  wire   [3:0] \MCInst_MC1_v3_0 ;
  wire   [3:0] \MCInst_MC1_v2_3 ;
  wire   [3:0] \MCInst_MC1_v2_2 ;
  wire   [3:0] \MCInst_MC1_v2_1 ;
  wire   [3:0] \MCInst_MC1_v2_0 ;
  wire   [3:0] \MCInst_MC1_v1_3 ;
  wire   [3:0] \MCInst_MC1_v1_2 ;
  wire   [3:0] \MCInst_MC1_v1_1 ;
  wire   [3:0] \MCInst_MC1_v1_0 ;
  wire   [3:0] \MCInst_MC1_v0_3 ;
  wire   [3:0] \MCInst_MC1_v0_2 ;
  wire   [3:0] \MCInst_MC1_v0_1 ;
  wire   [3:0] \MCInst_MC1_v0_0 ;
  wire   [3:0] \MCInst_MC2_v3_3 ;
  wire   [3:0] \MCInst_MC2_v3_2 ;
  wire   [3:0] \MCInst_MC2_v3_1 ;
  wire   [3:0] \MCInst_MC2_v3_0 ;
  wire   [3:0] \MCInst_MC2_v2_3 ;
  wire   [3:0] \MCInst_MC2_v2_2 ;
  wire   [3:0] \MCInst_MC2_v2_1 ;
  wire   [3:0] \MCInst_MC2_v2_0 ;
  wire   [3:0] \MCInst_MC2_v1_3 ;
  wire   [3:0] \MCInst_MC2_v1_2 ;
  wire   [3:0] \MCInst_MC2_v1_1 ;
  wire   [3:0] \MCInst_MC2_v1_0 ;
  wire   [3:0] \MCInst_MC2_v0_3 ;
  wire   [3:0] \MCInst_MC2_v0_2 ;
  wire   [3:0] \MCInst_MC2_v0_1 ;
  wire   [3:0] \MCInst_MC2_v0_0 ;
  wire   [3:0] \MCInst_MC3_v3_3 ;
  wire   [3:0] \MCInst_MC3_v3_2 ;
  wire   [3:0] \MCInst_MC3_v3_1 ;
  wire   [3:0] \MCInst_MC3_v3_0 ;
  wire   [3:0] \MCInst_MC3_v2_3 ;
  wire   [3:0] \MCInst_MC3_v2_2 ;
  wire   [3:0] \MCInst_MC3_v2_1 ;
  wire   [3:0] \MCInst_MC3_v2_0 ;
  wire   [3:0] \MCInst_MC3_v1_3 ;
  wire   [3:0] \MCInst_MC3_v1_2 ;
  wire   [3:0] \MCInst_MC3_v1_1 ;
  wire   [3:0] \MCInst_MC3_v1_0 ;
  wire   [3:0] \MCInst_MC3_v0_3 ;
  wire   [3:0] \MCInst_MC3_v0_2 ;
  wire   [3:0] \MCInst_MC3_v0_1 ;
  wire   [3:0] \MCInst_MC3_v0_0 ;
  wire   [2:0] \Red_MCInst_MC0_v3_3 ;
  wire   [2:0] \Red_MCInst_MC0_v3_2 ;
  wire   [2:0] \Red_MCInst_MC0_v3_1 ;
  wire   [2:0] \Red_MCInst_MC0_v3_0 ;
  wire   [2:0] \Red_MCInst_MC0_v2_3 ;
  wire   [2:0] \Red_MCInst_MC0_v2_2 ;
  wire   [2:0] \Red_MCInst_MC0_v2_1 ;
  wire   [2:0] \Red_MCInst_MC0_v2_0 ;
  wire   [2:0] \Red_MCInst_MC0_v1_3 ;
  wire   [2:0] \Red_MCInst_MC0_v1_2 ;
  wire   [2:0] \Red_MCInst_MC0_v1_1 ;
  wire   [2:0] \Red_MCInst_MC0_v1_0 ;
  wire   [2:0] \Red_MCInst_MC0_v0_3 ;
  wire   [2:0] \Red_MCInst_MC0_v0_2 ;
  wire   [2:0] \Red_MCInst_MC0_v0_1 ;
  wire   [2:0] \Red_MCInst_MC0_v0_0 ;
  wire   [2:0] \Red_MCInst_MC1_v3_3 ;
  wire   [2:0] \Red_MCInst_MC1_v3_2 ;
  wire   [2:0] \Red_MCInst_MC1_v3_1 ;
  wire   [2:0] \Red_MCInst_MC1_v3_0 ;
  wire   [2:0] \Red_MCInst_MC1_v2_3 ;
  wire   [2:0] \Red_MCInst_MC1_v2_2 ;
  wire   [2:0] \Red_MCInst_MC1_v2_1 ;
  wire   [2:0] \Red_MCInst_MC1_v2_0 ;
  wire   [2:0] \Red_MCInst_MC1_v1_3 ;
  wire   [2:0] \Red_MCInst_MC1_v1_2 ;
  wire   [2:0] \Red_MCInst_MC1_v1_1 ;
  wire   [2:0] \Red_MCInst_MC1_v1_0 ;
  wire   [2:0] \Red_MCInst_MC1_v0_3 ;
  wire   [2:0] \Red_MCInst_MC1_v0_2 ;
  wire   [2:0] \Red_MCInst_MC1_v0_1 ;
  wire   [2:0] \Red_MCInst_MC1_v0_0 ;
  wire   [2:0] \Red_MCInst_MC2_v3_3 ;
  wire   [2:0] \Red_MCInst_MC2_v3_2 ;
  wire   [2:0] \Red_MCInst_MC2_v3_1 ;
  wire   [2:0] \Red_MCInst_MC2_v3_0 ;
  wire   [2:0] \Red_MCInst_MC2_v2_3 ;
  wire   [2:0] \Red_MCInst_MC2_v2_2 ;
  wire   [2:0] \Red_MCInst_MC2_v2_1 ;
  wire   [2:0] \Red_MCInst_MC2_v2_0 ;
  wire   [2:0] \Red_MCInst_MC2_v1_3 ;
  wire   [2:0] \Red_MCInst_MC2_v1_2 ;
  wire   [2:0] \Red_MCInst_MC2_v1_1 ;
  wire   [2:0] \Red_MCInst_MC2_v1_0 ;
  wire   [2:0] \Red_MCInst_MC2_v0_3 ;
  wire   [2:0] \Red_MCInst_MC2_v0_2 ;
  wire   [2:0] \Red_MCInst_MC2_v0_1 ;
  wire   [2:0] \Red_MCInst_MC2_v0_0 ;
  wire   [2:0] \Red_MCInst_MC3_v3_3 ;
  wire   [2:0] \Red_MCInst_MC3_v3_2 ;
  wire   [2:0] \Red_MCInst_MC3_v3_1 ;
  wire   [2:0] \Red_MCInst_MC3_v3_0 ;
  wire   [2:0] \Red_MCInst_MC3_v2_3 ;
  wire   [2:0] \Red_MCInst_MC3_v2_2 ;
  wire   [2:0] \Red_MCInst_MC3_v2_1 ;
  wire   [2:0] \Red_MCInst_MC3_v2_0 ;
  wire   [2:0] \Red_MCInst_MC3_v1_3 ;
  wire   [2:0] \Red_MCInst_MC3_v1_2 ;
  wire   [2:0] \Red_MCInst_MC3_v1_1 ;
  wire   [2:0] \Red_MCInst_MC3_v1_0 ;
  wire   [2:0] \Red_MCInst_MC3_v0_3 ;
  wire   [2:0] \Red_MCInst_MC3_v0_2 ;
  wire   [2:0] \Red_MCInst_MC3_v0_1 ;
  wire   [2:0] \Red_MCInst_MC3_v0_0 ;

  AND2_X1 U7 ( .A1(Error[2]), .A2(Error[0]), .ZN(n149) );
  NAND2_X1 U8 ( .A1(Error[1]), .A2(n149), .ZN(ErrorFlag) );
  INV_X1 \AddKeyXOR_XORInst_0_0_U2  ( .A(\AddKeyXOR_XORInst_0_0_n2 ), .ZN(
        AddRoundKeyOutput[0]) );
  XNOR2_X1 \AddKeyXOR_XORInst_0_0_U1  ( .A(Plaintext[0]), .B(Key[0]), .ZN(
        \AddKeyXOR_XORInst_0_0_n2 ) );
  XOR2_X2 \AddKeyXOR_XORInst_0_1_U1  ( .A(Plaintext[1]), .B(Key[1]), .Z(
        AddRoundKeyOutput[1]) );
  INV_X1 \AddKeyXOR_XORInst_0_2_U2  ( .A(\AddKeyXOR_XORInst_0_2_n2 ), .ZN(
        AddRoundKeyOutput[2]) );
  XNOR2_X1 \AddKeyXOR_XORInst_0_2_U1  ( .A(Plaintext[2]), .B(Key[2]), .ZN(
        \AddKeyXOR_XORInst_0_2_n2 ) );
  XOR2_X1 \AddKeyXOR_XORInst_0_3_U1  ( .A(Plaintext[3]), .B(Key[3]), .Z(
        AddRoundKeyOutput[3]) );
  XOR2_X2 \AddKeyXOR_XORInst_1_0_U1  ( .A(Plaintext[4]), .B(Key[4]), .Z(
        AddRoundKeyOutput[4]) );
  XOR2_X2 \AddKeyXOR_XORInst_1_1_U1  ( .A(Plaintext[5]), .B(Key[5]), .Z(
        AddRoundKeyOutput[5]) );
  INV_X1 \AddKeyXOR_XORInst_1_2_U2  ( .A(\AddKeyXOR_XORInst_1_2_n2 ), .ZN(
        AddRoundKeyOutput[6]) );
  XNOR2_X1 \AddKeyXOR_XORInst_1_2_U1  ( .A(Plaintext[6]), .B(Key[6]), .ZN(
        \AddKeyXOR_XORInst_1_2_n2 ) );
  XOR2_X1 \AddKeyXOR_XORInst_1_3_U1  ( .A(Plaintext[7]), .B(Key[7]), .Z(
        AddRoundKeyOutput[7]) );
  XOR2_X2 \AddKeyXOR_XORInst_2_0_U1  ( .A(Plaintext[8]), .B(Key[8]), .Z(
        AddRoundKeyOutput[8]) );
  XOR2_X2 \AddKeyXOR_XORInst_2_1_U1  ( .A(Plaintext[9]), .B(Key[9]), .Z(
        AddRoundKeyOutput[9]) );
  INV_X1 \AddKeyXOR_XORInst_2_2_U2  ( .A(\AddKeyXOR_XORInst_2_2_n2 ), .ZN(
        AddRoundKeyOutput[10]) );
  XNOR2_X1 \AddKeyXOR_XORInst_2_2_U1  ( .A(Plaintext[10]), .B(Key[10]), .ZN(
        \AddKeyXOR_XORInst_2_2_n2 ) );
  XOR2_X1 \AddKeyXOR_XORInst_2_3_U1  ( .A(Plaintext[11]), .B(Key[11]), .Z(
        AddRoundKeyOutput[11]) );
  XOR2_X2 \AddKeyXOR_XORInst_3_0_U1  ( .A(Plaintext[12]), .B(Key[12]), .Z(
        AddRoundKeyOutput[12]) );
  XOR2_X2 \AddKeyXOR_XORInst_3_1_U1  ( .A(Plaintext[13]), .B(Key[13]), .Z(
        AddRoundKeyOutput[13]) );
  INV_X1 \AddKeyXOR_XORInst_3_2_U2  ( .A(\AddKeyXOR_XORInst_3_2_n2 ), .ZN(
        AddRoundKeyOutput[14]) );
  XNOR2_X1 \AddKeyXOR_XORInst_3_2_U1  ( .A(Plaintext[14]), .B(Key[14]), .ZN(
        \AddKeyXOR_XORInst_3_2_n2 ) );
  XOR2_X1 \AddKeyXOR_XORInst_3_3_U1  ( .A(Plaintext[15]), .B(Key[15]), .Z(
        AddRoundKeyOutput[15]) );
  XOR2_X2 \AddKeyXOR_XORInst_4_0_U1  ( .A(Plaintext[16]), .B(Key[16]), .Z(
        AddRoundKeyOutput[16]) );
  XOR2_X2 \AddKeyXOR_XORInst_4_1_U1  ( .A(Plaintext[17]), .B(Key[17]), .Z(
        AddRoundKeyOutput[17]) );
  INV_X1 \AddKeyXOR_XORInst_4_2_U2  ( .A(\AddKeyXOR_XORInst_4_2_n2 ), .ZN(
        AddRoundKeyOutput[18]) );
  XNOR2_X1 \AddKeyXOR_XORInst_4_2_U1  ( .A(Plaintext[18]), .B(Key[18]), .ZN(
        \AddKeyXOR_XORInst_4_2_n2 ) );
  XOR2_X1 \AddKeyXOR_XORInst_4_3_U1  ( .A(Plaintext[19]), .B(Key[19]), .Z(
        AddRoundKeyOutput[19]) );
  XOR2_X2 \AddKeyXOR_XORInst_5_0_U1  ( .A(Plaintext[20]), .B(Key[20]), .Z(
        AddRoundKeyOutput[20]) );
  XOR2_X2 \AddKeyXOR_XORInst_5_1_U1  ( .A(Plaintext[21]), .B(Key[21]), .Z(
        AddRoundKeyOutput[21]) );
  INV_X1 \AddKeyXOR_XORInst_5_2_U2  ( .A(\AddKeyXOR_XORInst_5_2_n2 ), .ZN(
        AddRoundKeyOutput[22]) );
  XNOR2_X1 \AddKeyXOR_XORInst_5_2_U1  ( .A(Plaintext[22]), .B(Key[22]), .ZN(
        \AddKeyXOR_XORInst_5_2_n2 ) );
  XOR2_X1 \AddKeyXOR_XORInst_5_3_U1  ( .A(Plaintext[23]), .B(Key[23]), .Z(
        AddRoundKeyOutput[23]) );
  XOR2_X2 \AddKeyXOR_XORInst_6_0_U1  ( .A(Plaintext[24]), .B(Key[24]), .Z(
        AddRoundKeyOutput[24]) );
  XOR2_X2 \AddKeyXOR_XORInst_6_1_U1  ( .A(Plaintext[25]), .B(Key[25]), .Z(
        AddRoundKeyOutput[25]) );
  INV_X1 \AddKeyXOR_XORInst_6_2_U2  ( .A(\AddKeyXOR_XORInst_6_2_n2 ), .ZN(
        AddRoundKeyOutput[26]) );
  XNOR2_X1 \AddKeyXOR_XORInst_6_2_U1  ( .A(Plaintext[26]), .B(Key[26]), .ZN(
        \AddKeyXOR_XORInst_6_2_n2 ) );
  XOR2_X1 \AddKeyXOR_XORInst_6_3_U1  ( .A(Plaintext[27]), .B(Key[27]), .Z(
        AddRoundKeyOutput[27]) );
  XOR2_X2 \AddKeyXOR_XORInst_7_0_U1  ( .A(Plaintext[28]), .B(Key[28]), .Z(
        AddRoundKeyOutput[28]) );
  XOR2_X2 \AddKeyXOR_XORInst_7_1_U1  ( .A(Plaintext[29]), .B(Key[29]), .Z(
        AddRoundKeyOutput[29]) );
  INV_X1 \AddKeyXOR_XORInst_7_2_U2  ( .A(\AddKeyXOR_XORInst_7_2_n2 ), .ZN(
        AddRoundKeyOutput[30]) );
  XNOR2_X1 \AddKeyXOR_XORInst_7_2_U1  ( .A(Plaintext[30]), .B(Key[30]), .ZN(
        \AddKeyXOR_XORInst_7_2_n2 ) );
  XOR2_X1 \AddKeyXOR_XORInst_7_3_U1  ( .A(Plaintext[31]), .B(Key[31]), .Z(
        AddRoundKeyOutput[31]) );
  XOR2_X2 \AddKeyXOR_XORInst_8_0_U1  ( .A(Plaintext[32]), .B(Key[32]), .Z(
        AddRoundKeyOutput[32]) );
  XOR2_X2 \AddKeyXOR_XORInst_8_1_U1  ( .A(Plaintext[33]), .B(Key[33]), .Z(
        AddRoundKeyOutput[33]) );
  INV_X1 \AddKeyXOR_XORInst_8_2_U2  ( .A(\AddKeyXOR_XORInst_8_2_n2 ), .ZN(
        AddRoundKeyOutput[34]) );
  XNOR2_X1 \AddKeyXOR_XORInst_8_2_U1  ( .A(Plaintext[34]), .B(Key[34]), .ZN(
        \AddKeyXOR_XORInst_8_2_n2 ) );
  XOR2_X1 \AddKeyXOR_XORInst_8_3_U1  ( .A(Plaintext[35]), .B(Key[35]), .Z(
        AddRoundKeyOutput[35]) );
  XOR2_X2 \AddKeyXOR_XORInst_9_0_U1  ( .A(Plaintext[36]), .B(Key[36]), .Z(
        AddRoundKeyOutput[36]) );
  XOR2_X2 \AddKeyXOR_XORInst_9_1_U1  ( .A(Plaintext[37]), .B(Key[37]), .Z(
        AddRoundKeyOutput[37]) );
  INV_X1 \AddKeyXOR_XORInst_9_2_U2  ( .A(\AddKeyXOR_XORInst_9_2_n2 ), .ZN(
        AddRoundKeyOutput[38]) );
  XNOR2_X1 \AddKeyXOR_XORInst_9_2_U1  ( .A(Plaintext[38]), .B(Key[38]), .ZN(
        \AddKeyXOR_XORInst_9_2_n2 ) );
  XOR2_X1 \AddKeyXOR_XORInst_9_3_U1  ( .A(Plaintext[39]), .B(Key[39]), .Z(
        AddRoundKeyOutput[39]) );
  XOR2_X2 \AddKeyXOR_XORInst_10_0_U1  ( .A(Plaintext[40]), .B(Key[40]), .Z(
        AddRoundKeyOutput[40]) );
  XOR2_X2 \AddKeyXOR_XORInst_10_1_U1  ( .A(Plaintext[41]), .B(Key[41]), .Z(
        AddRoundKeyOutput[41]) );
  INV_X1 \AddKeyXOR_XORInst_10_2_U2  ( .A(\AddKeyXOR_XORInst_10_2_n2 ), .ZN(
        AddRoundKeyOutput[42]) );
  XNOR2_X1 \AddKeyXOR_XORInst_10_2_U1  ( .A(Plaintext[42]), .B(Key[42]), .ZN(
        \AddKeyXOR_XORInst_10_2_n2 ) );
  XOR2_X1 \AddKeyXOR_XORInst_10_3_U1  ( .A(Plaintext[43]), .B(Key[43]), .Z(
        AddRoundKeyOutput[43]) );
  XOR2_X2 \AddKeyXOR_XORInst_11_0_U1  ( .A(Plaintext[44]), .B(Key[44]), .Z(
        AddRoundKeyOutput[44]) );
  XOR2_X2 \AddKeyXOR_XORInst_11_1_U1  ( .A(Plaintext[45]), .B(Key[45]), .Z(
        AddRoundKeyOutput[45]) );
  INV_X1 \AddKeyXOR_XORInst_11_2_U2  ( .A(\AddKeyXOR_XORInst_11_2_n2 ), .ZN(
        AddRoundKeyOutput[46]) );
  XNOR2_X1 \AddKeyXOR_XORInst_11_2_U1  ( .A(Plaintext[46]), .B(Key[46]), .ZN(
        \AddKeyXOR_XORInst_11_2_n2 ) );
  XOR2_X1 \AddKeyXOR_XORInst_11_3_U1  ( .A(Plaintext[47]), .B(Key[47]), .Z(
        AddRoundKeyOutput[47]) );
  XOR2_X2 \AddKeyXOR_XORInst_12_0_U1  ( .A(Plaintext[48]), .B(Key[48]), .Z(
        AddRoundKeyOutput[48]) );
  XOR2_X2 \AddKeyXOR_XORInst_12_1_U1  ( .A(Plaintext[49]), .B(Key[49]), .Z(
        AddRoundKeyOutput[49]) );
  INV_X1 \AddKeyXOR_XORInst_12_2_U2  ( .A(\AddKeyXOR_XORInst_12_2_n2 ), .ZN(
        AddRoundKeyOutput[50]) );
  XNOR2_X1 \AddKeyXOR_XORInst_12_2_U1  ( .A(Plaintext[50]), .B(Key[50]), .ZN(
        \AddKeyXOR_XORInst_12_2_n2 ) );
  XOR2_X1 \AddKeyXOR_XORInst_12_3_U1  ( .A(Plaintext[51]), .B(Key[51]), .Z(
        AddRoundKeyOutput[51]) );
  XOR2_X2 \AddKeyXOR_XORInst_13_0_U1  ( .A(Plaintext[52]), .B(Key[52]), .Z(
        AddRoundKeyOutput[52]) );
  XOR2_X2 \AddKeyXOR_XORInst_13_1_U1  ( .A(Plaintext[53]), .B(Key[53]), .Z(
        AddRoundKeyOutput[53]) );
  INV_X1 \AddKeyXOR_XORInst_13_2_U2  ( .A(\AddKeyXOR_XORInst_13_2_n2 ), .ZN(
        AddRoundKeyOutput[54]) );
  XNOR2_X1 \AddKeyXOR_XORInst_13_2_U1  ( .A(Plaintext[54]), .B(Key[54]), .ZN(
        \AddKeyXOR_XORInst_13_2_n2 ) );
  XOR2_X1 \AddKeyXOR_XORInst_13_3_U1  ( .A(Plaintext[55]), .B(Key[55]), .Z(
        AddRoundKeyOutput[55]) );
  XOR2_X2 \AddKeyXOR_XORInst_14_0_U1  ( .A(Plaintext[56]), .B(Key[56]), .Z(
        AddRoundKeyOutput[56]) );
  XOR2_X2 \AddKeyXOR_XORInst_14_1_U1  ( .A(Plaintext[57]), .B(Key[57]), .Z(
        AddRoundKeyOutput[57]) );
  INV_X1 \AddKeyXOR_XORInst_14_2_U2  ( .A(\AddKeyXOR_XORInst_14_2_n2 ), .ZN(
        AddRoundKeyOutput[58]) );
  XNOR2_X1 \AddKeyXOR_XORInst_14_2_U1  ( .A(Plaintext[58]), .B(Key[58]), .ZN(
        \AddKeyXOR_XORInst_14_2_n2 ) );
  XOR2_X1 \AddKeyXOR_XORInst_14_3_U1  ( .A(Plaintext[59]), .B(Key[59]), .Z(
        AddRoundKeyOutput[59]) );
  XOR2_X2 \AddKeyXOR_XORInst_15_0_U1  ( .A(Plaintext[60]), .B(Key[60]), .Z(
        AddRoundKeyOutput[60]) );
  XOR2_X2 \AddKeyXOR_XORInst_15_1_U1  ( .A(Plaintext[61]), .B(Key[61]), .Z(
        AddRoundKeyOutput[61]) );
  INV_X1 \AddKeyXOR_XORInst_15_2_U2  ( .A(\AddKeyXOR_XORInst_15_2_n2 ), .ZN(
        AddRoundKeyOutput[62]) );
  XNOR2_X1 \AddKeyXOR_XORInst_15_2_U1  ( .A(Plaintext[62]), .B(Key[62]), .ZN(
        \AddKeyXOR_XORInst_15_2_n2 ) );
  XOR2_X1 \AddKeyXOR_XORInst_15_3_U1  ( .A(Plaintext[63]), .B(Key[63]), .Z(
        AddRoundKeyOutput[63]) );
  NAND2_X1 \SubCellInst_LFInst_0_LFInst_0_U7  ( .A1(AddRoundKeyOutput[2]), 
        .A2(\SubCellInst_LFInst_0_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_0_LFInst_0_n8 ) );
  INV_X1 \SubCellInst_LFInst_0_LFInst_0_U6  ( .A(AddRoundKeyOutput[1]), .ZN(
        \SubCellInst_LFInst_0_LFInst_0_n7 ) );
  XOR2_X1 \SubCellInst_LFInst_0_LFInst_0_U5  ( .A(AddRoundKeyOutput[0]), .B(
        AddRoundKeyOutput[3]), .Z(\SubCellInst_LFInst_0_LFInst_0_n9 ) );
  INV_X1 \SubCellInst_LFInst_0_LFInst_0_U4  ( .A(
        \SubCellInst_LFInst_0_LFInst_0_n10 ), .ZN(\MCInst_MC0_v3_2 [3]) );
  XOR2_X1 \SubCellInst_LFInst_0_LFInst_0_U3  ( .A(
        \SubCellInst_LFInst_0_LFInst_0_n9 ), .B(
        \SubCellInst_LFInst_0_LFInst_0_n8 ), .Z(
        \SubCellInst_LFInst_0_LFInst_0_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_0_LFInst_1_U12  ( .A1(
        \SubCellInst_LFInst_0_LFInst_1_n18 ), .A2(
        \SubCellInst_LFInst_0_LFInst_1_n17 ), .ZN(\Red_MCInst_MC0_v3_3 [2]) );
  NAND2_X1 \SubCellInst_LFInst_0_LFInst_1_U11  ( .A1(AddRoundKeyOutput[1]), 
        .A2(\SubCellInst_LFInst_0_LFInst_1_n16 ), .ZN(
        \SubCellInst_LFInst_0_LFInst_1_n17 ) );
  NOR2_X1 \SubCellInst_LFInst_0_LFInst_1_U10  ( .A1(AddRoundKeyOutput[3]), 
        .A2(\SubCellInst_LFInst_0_LFInst_1_n15 ), .ZN(
        \SubCellInst_LFInst_0_LFInst_1_n16 ) );
  AND2_X1 \SubCellInst_LFInst_0_LFInst_1_U9  ( .A1(AddRoundKeyOutput[0]), .A2(
        AddRoundKeyOutput[2]), .ZN(\SubCellInst_LFInst_0_LFInst_1_n15 ) );
  NAND2_X1 \SubCellInst_LFInst_0_LFInst_1_U8  ( .A1(AddRoundKeyOutput[3]), 
        .A2(\SubCellInst_LFInst_0_LFInst_1_n14 ), .ZN(
        \SubCellInst_LFInst_0_LFInst_1_n18 ) );
  NAND2_X1 \SubCellInst_LFInst_0_LFInst_1_U7  ( .A1(
        \SubCellInst_LFInst_0_LFInst_1_n13 ), .A2(
        \SubCellInst_LFInst_0_LFInst_1_n12 ), .ZN(
        \SubCellInst_LFInst_0_LFInst_1_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_0_LFInst_1_U6  ( .A1(AddRoundKeyOutput[0]), 
        .A2(AddRoundKeyOutput[2]), .ZN(\SubCellInst_LFInst_0_LFInst_1_n12 ) );
  NAND2_X1 \SubCellInst_LFInst_0_LFInst_1_U5  ( .A1(
        \SubCellInst_LFInst_0_LFInst_1_n11 ), .A2(
        \SubCellInst_LFInst_0_LFInst_1_n10 ), .ZN(
        \SubCellInst_LFInst_0_LFInst_1_n13 ) );
  NAND2_X1 \SubCellInst_LFInst_0_LFInst_1_U4  ( .A1(AddRoundKeyOutput[0]), 
        .A2(AddRoundKeyOutput[1]), .ZN(\SubCellInst_LFInst_0_LFInst_1_n10 ) );
  INV_X1 \SubCellInst_LFInst_0_LFInst_1_U3  ( .A(AddRoundKeyOutput[2]), .ZN(
        \SubCellInst_LFInst_0_LFInst_1_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_0_LFInst_2_U11  ( .A1(
        \SubCellInst_LFInst_0_LFInst_2_n22 ), .A2(
        \SubCellInst_LFInst_0_LFInst_2_n21 ), .ZN(\MCInst_MC0_v3_0 [3]) );
  NAND2_X1 \SubCellInst_LFInst_0_LFInst_2_U10  ( .A1(AddRoundKeyOutput[2]), 
        .A2(\SubCellInst_LFInst_0_LFInst_2_n20 ), .ZN(
        \SubCellInst_LFInst_0_LFInst_2_n21 ) );
  NOR2_X1 \SubCellInst_LFInst_0_LFInst_2_U9  ( .A1(AddRoundKeyOutput[1]), .A2(
        \SubCellInst_LFInst_0_LFInst_2_n19 ), .ZN(
        \SubCellInst_LFInst_0_LFInst_2_n20 ) );
  INV_X1 \SubCellInst_LFInst_0_LFInst_2_U8  ( .A(AddRoundKeyOutput[3]), .ZN(
        \SubCellInst_LFInst_0_LFInst_2_n19 ) );
  NAND2_X1 \SubCellInst_LFInst_0_LFInst_2_U7  ( .A1(
        \SubCellInst_LFInst_0_LFInst_2_n18 ), .A2(
        \SubCellInst_LFInst_0_LFInst_2_n17 ), .ZN(
        \SubCellInst_LFInst_0_LFInst_2_n22 ) );
  XOR2_X1 \SubCellInst_LFInst_0_LFInst_2_U6  ( .A(
        \SubCellInst_LFInst_0_LFInst_2_n16 ), .B(AddRoundKeyOutput[2]), .Z(
        \SubCellInst_LFInst_0_LFInst_2_n17 ) );
  NAND2_X1 \SubCellInst_LFInst_0_LFInst_2_U5  ( .A1(AddRoundKeyOutput[0]), 
        .A2(AddRoundKeyOutput[1]), .ZN(\SubCellInst_LFInst_0_LFInst_2_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_0_LFInst_2_U4  ( .A1(
        \SubCellInst_LFInst_0_LFInst_2_n15 ), .A2(AddRoundKeyOutput[3]), .ZN(
        \SubCellInst_LFInst_0_LFInst_2_n18 ) );
  XNOR2_X1 \SubCellInst_LFInst_0_LFInst_2_U3  ( .A(AddRoundKeyOutput[0]), .B(
        AddRoundKeyOutput[1]), .ZN(\SubCellInst_LFInst_0_LFInst_2_n15 ) );
  NAND2_X1 \SubCellInst_LFInst_0_LFInst_3_U9  ( .A1(
        \SubCellInst_LFInst_0_LFInst_3_n16 ), .A2(
        \SubCellInst_LFInst_0_LFInst_3_n15 ), .ZN(\Red_MCInst_MC0_v3_1 [2]) );
  NAND2_X1 \SubCellInst_LFInst_0_LFInst_3_U8  ( .A1(AddRoundKeyOutput[1]), 
        .A2(\SubCellInst_LFInst_0_LFInst_3_n14 ), .ZN(
        \SubCellInst_LFInst_0_LFInst_3_n15 ) );
  XOR2_X1 \SubCellInst_LFInst_0_LFInst_3_U7  ( .A(AddRoundKeyOutput[3]), .B(
        AddRoundKeyOutput[2]), .Z(\SubCellInst_LFInst_0_LFInst_3_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_0_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_0_LFInst_3_n13 ), .A2(
        \SubCellInst_LFInst_0_LFInst_3_n12 ), .ZN(
        \SubCellInst_LFInst_0_LFInst_3_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_0_LFInst_3_U5  ( .A1(AddRoundKeyOutput[0]), 
        .A2(AddRoundKeyOutput[2]), .ZN(\SubCellInst_LFInst_0_LFInst_3_n12 ) );
  XNOR2_X1 \SubCellInst_LFInst_0_LFInst_3_U4  ( .A(AddRoundKeyOutput[0]), .B(
        \SubCellInst_LFInst_0_LFInst_3_n11 ), .ZN(
        \SubCellInst_LFInst_0_LFInst_3_n13 ) );
  OR2_X1 \SubCellInst_LFInst_0_LFInst_3_U3  ( .A1(AddRoundKeyOutput[3]), .A2(
        AddRoundKeyOutput[1]), .ZN(\SubCellInst_LFInst_0_LFInst_3_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_1_LFInst_0_U7  ( .A1(AddRoundKeyOutput[6]), 
        .A2(\SubCellInst_LFInst_1_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_1_LFInst_0_n8 ) );
  INV_X1 \SubCellInst_LFInst_1_LFInst_0_U6  ( .A(AddRoundKeyOutput[5]), .ZN(
        \SubCellInst_LFInst_1_LFInst_0_n7 ) );
  XOR2_X1 \SubCellInst_LFInst_1_LFInst_0_U5  ( .A(AddRoundKeyOutput[4]), .B(
        AddRoundKeyOutput[7]), .Z(\SubCellInst_LFInst_1_LFInst_0_n9 ) );
  INV_X1 \SubCellInst_LFInst_1_LFInst_0_U4  ( .A(
        \SubCellInst_LFInst_1_LFInst_0_n10 ), .ZN(\MCInst_MC3_v3_2 [3]) );
  XOR2_X1 \SubCellInst_LFInst_1_LFInst_0_U3  ( .A(
        \SubCellInst_LFInst_1_LFInst_0_n9 ), .B(
        \SubCellInst_LFInst_1_LFInst_0_n8 ), .Z(
        \SubCellInst_LFInst_1_LFInst_0_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_1_LFInst_1_U12  ( .A1(
        \SubCellInst_LFInst_1_LFInst_1_n18 ), .A2(
        \SubCellInst_LFInst_1_LFInst_1_n17 ), .ZN(\Red_MCInst_MC3_v3_3 [2]) );
  NAND2_X1 \SubCellInst_LFInst_1_LFInst_1_U11  ( .A1(AddRoundKeyOutput[5]), 
        .A2(\SubCellInst_LFInst_1_LFInst_1_n16 ), .ZN(
        \SubCellInst_LFInst_1_LFInst_1_n17 ) );
  NOR2_X1 \SubCellInst_LFInst_1_LFInst_1_U10  ( .A1(AddRoundKeyOutput[7]), 
        .A2(\SubCellInst_LFInst_1_LFInst_1_n15 ), .ZN(
        \SubCellInst_LFInst_1_LFInst_1_n16 ) );
  AND2_X1 \SubCellInst_LFInst_1_LFInst_1_U9  ( .A1(AddRoundKeyOutput[4]), .A2(
        AddRoundKeyOutput[6]), .ZN(\SubCellInst_LFInst_1_LFInst_1_n15 ) );
  NAND2_X1 \SubCellInst_LFInst_1_LFInst_1_U8  ( .A1(AddRoundKeyOutput[7]), 
        .A2(\SubCellInst_LFInst_1_LFInst_1_n14 ), .ZN(
        \SubCellInst_LFInst_1_LFInst_1_n18 ) );
  NAND2_X1 \SubCellInst_LFInst_1_LFInst_1_U7  ( .A1(
        \SubCellInst_LFInst_1_LFInst_1_n13 ), .A2(
        \SubCellInst_LFInst_1_LFInst_1_n12 ), .ZN(
        \SubCellInst_LFInst_1_LFInst_1_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_1_LFInst_1_U6  ( .A1(AddRoundKeyOutput[4]), 
        .A2(AddRoundKeyOutput[6]), .ZN(\SubCellInst_LFInst_1_LFInst_1_n12 ) );
  NAND2_X1 \SubCellInst_LFInst_1_LFInst_1_U5  ( .A1(
        \SubCellInst_LFInst_1_LFInst_1_n11 ), .A2(
        \SubCellInst_LFInst_1_LFInst_1_n10 ), .ZN(
        \SubCellInst_LFInst_1_LFInst_1_n13 ) );
  NAND2_X1 \SubCellInst_LFInst_1_LFInst_1_U4  ( .A1(AddRoundKeyOutput[4]), 
        .A2(AddRoundKeyOutput[5]), .ZN(\SubCellInst_LFInst_1_LFInst_1_n10 ) );
  INV_X1 \SubCellInst_LFInst_1_LFInst_1_U3  ( .A(AddRoundKeyOutput[6]), .ZN(
        \SubCellInst_LFInst_1_LFInst_1_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_1_LFInst_2_U11  ( .A1(
        \SubCellInst_LFInst_1_LFInst_2_n22 ), .A2(
        \SubCellInst_LFInst_1_LFInst_2_n21 ), .ZN(\MCInst_MC3_v3_0 [3]) );
  NAND2_X1 \SubCellInst_LFInst_1_LFInst_2_U10  ( .A1(AddRoundKeyOutput[6]), 
        .A2(\SubCellInst_LFInst_1_LFInst_2_n20 ), .ZN(
        \SubCellInst_LFInst_1_LFInst_2_n21 ) );
  NOR2_X1 \SubCellInst_LFInst_1_LFInst_2_U9  ( .A1(AddRoundKeyOutput[5]), .A2(
        \SubCellInst_LFInst_1_LFInst_2_n19 ), .ZN(
        \SubCellInst_LFInst_1_LFInst_2_n20 ) );
  INV_X1 \SubCellInst_LFInst_1_LFInst_2_U8  ( .A(AddRoundKeyOutput[7]), .ZN(
        \SubCellInst_LFInst_1_LFInst_2_n19 ) );
  NAND2_X1 \SubCellInst_LFInst_1_LFInst_2_U7  ( .A1(
        \SubCellInst_LFInst_1_LFInst_2_n18 ), .A2(
        \SubCellInst_LFInst_1_LFInst_2_n17 ), .ZN(
        \SubCellInst_LFInst_1_LFInst_2_n22 ) );
  XOR2_X1 \SubCellInst_LFInst_1_LFInst_2_U6  ( .A(
        \SubCellInst_LFInst_1_LFInst_2_n16 ), .B(AddRoundKeyOutput[6]), .Z(
        \SubCellInst_LFInst_1_LFInst_2_n17 ) );
  NAND2_X1 \SubCellInst_LFInst_1_LFInst_2_U5  ( .A1(AddRoundKeyOutput[4]), 
        .A2(AddRoundKeyOutput[5]), .ZN(\SubCellInst_LFInst_1_LFInst_2_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_1_LFInst_2_U4  ( .A1(
        \SubCellInst_LFInst_1_LFInst_2_n15 ), .A2(AddRoundKeyOutput[7]), .ZN(
        \SubCellInst_LFInst_1_LFInst_2_n18 ) );
  XNOR2_X1 \SubCellInst_LFInst_1_LFInst_2_U3  ( .A(AddRoundKeyOutput[4]), .B(
        AddRoundKeyOutput[5]), .ZN(\SubCellInst_LFInst_1_LFInst_2_n15 ) );
  NAND2_X1 \SubCellInst_LFInst_1_LFInst_3_U9  ( .A1(
        \SubCellInst_LFInst_1_LFInst_3_n16 ), .A2(
        \SubCellInst_LFInst_1_LFInst_3_n15 ), .ZN(\Red_MCInst_MC3_v3_1 [2]) );
  NAND2_X1 \SubCellInst_LFInst_1_LFInst_3_U8  ( .A1(AddRoundKeyOutput[5]), 
        .A2(\SubCellInst_LFInst_1_LFInst_3_n14 ), .ZN(
        \SubCellInst_LFInst_1_LFInst_3_n15 ) );
  XOR2_X1 \SubCellInst_LFInst_1_LFInst_3_U7  ( .A(AddRoundKeyOutput[7]), .B(
        AddRoundKeyOutput[6]), .Z(\SubCellInst_LFInst_1_LFInst_3_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_1_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_1_LFInst_3_n13 ), .A2(
        \SubCellInst_LFInst_1_LFInst_3_n12 ), .ZN(
        \SubCellInst_LFInst_1_LFInst_3_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_1_LFInst_3_U5  ( .A1(AddRoundKeyOutput[4]), 
        .A2(AddRoundKeyOutput[6]), .ZN(\SubCellInst_LFInst_1_LFInst_3_n12 ) );
  XNOR2_X1 \SubCellInst_LFInst_1_LFInst_3_U4  ( .A(AddRoundKeyOutput[4]), .B(
        \SubCellInst_LFInst_1_LFInst_3_n11 ), .ZN(
        \SubCellInst_LFInst_1_LFInst_3_n13 ) );
  OR2_X1 \SubCellInst_LFInst_1_LFInst_3_U3  ( .A1(AddRoundKeyOutput[7]), .A2(
        AddRoundKeyOutput[5]), .ZN(\SubCellInst_LFInst_1_LFInst_3_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_2_LFInst_0_U7  ( .A1(AddRoundKeyOutput[10]), 
        .A2(\SubCellInst_LFInst_2_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_2_LFInst_0_n8 ) );
  INV_X1 \SubCellInst_LFInst_2_LFInst_0_U6  ( .A(AddRoundKeyOutput[9]), .ZN(
        \SubCellInst_LFInst_2_LFInst_0_n7 ) );
  XOR2_X1 \SubCellInst_LFInst_2_LFInst_0_U5  ( .A(AddRoundKeyOutput[8]), .B(
        AddRoundKeyOutput[11]), .Z(\SubCellInst_LFInst_2_LFInst_0_n9 ) );
  INV_X1 \SubCellInst_LFInst_2_LFInst_0_U4  ( .A(
        \SubCellInst_LFInst_2_LFInst_0_n10 ), .ZN(\MCInst_MC2_v3_2 [3]) );
  XOR2_X1 \SubCellInst_LFInst_2_LFInst_0_U3  ( .A(
        \SubCellInst_LFInst_2_LFInst_0_n9 ), .B(
        \SubCellInst_LFInst_2_LFInst_0_n8 ), .Z(
        \SubCellInst_LFInst_2_LFInst_0_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_2_LFInst_1_U12  ( .A1(
        \SubCellInst_LFInst_2_LFInst_1_n18 ), .A2(
        \SubCellInst_LFInst_2_LFInst_1_n17 ), .ZN(\Red_MCInst_MC2_v3_3 [2]) );
  NAND2_X1 \SubCellInst_LFInst_2_LFInst_1_U11  ( .A1(AddRoundKeyOutput[9]), 
        .A2(\SubCellInst_LFInst_2_LFInst_1_n16 ), .ZN(
        \SubCellInst_LFInst_2_LFInst_1_n17 ) );
  NOR2_X1 \SubCellInst_LFInst_2_LFInst_1_U10  ( .A1(AddRoundKeyOutput[11]), 
        .A2(\SubCellInst_LFInst_2_LFInst_1_n15 ), .ZN(
        \SubCellInst_LFInst_2_LFInst_1_n16 ) );
  AND2_X1 \SubCellInst_LFInst_2_LFInst_1_U9  ( .A1(AddRoundKeyOutput[8]), .A2(
        AddRoundKeyOutput[10]), .ZN(\SubCellInst_LFInst_2_LFInst_1_n15 ) );
  NAND2_X1 \SubCellInst_LFInst_2_LFInst_1_U8  ( .A1(AddRoundKeyOutput[11]), 
        .A2(\SubCellInst_LFInst_2_LFInst_1_n14 ), .ZN(
        \SubCellInst_LFInst_2_LFInst_1_n18 ) );
  NAND2_X1 \SubCellInst_LFInst_2_LFInst_1_U7  ( .A1(
        \SubCellInst_LFInst_2_LFInst_1_n13 ), .A2(
        \SubCellInst_LFInst_2_LFInst_1_n12 ), .ZN(
        \SubCellInst_LFInst_2_LFInst_1_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_2_LFInst_1_U6  ( .A1(AddRoundKeyOutput[8]), 
        .A2(AddRoundKeyOutput[10]), .ZN(\SubCellInst_LFInst_2_LFInst_1_n12 )
         );
  NAND2_X1 \SubCellInst_LFInst_2_LFInst_1_U5  ( .A1(
        \SubCellInst_LFInst_2_LFInst_1_n11 ), .A2(
        \SubCellInst_LFInst_2_LFInst_1_n10 ), .ZN(
        \SubCellInst_LFInst_2_LFInst_1_n13 ) );
  NAND2_X1 \SubCellInst_LFInst_2_LFInst_1_U4  ( .A1(AddRoundKeyOutput[8]), 
        .A2(AddRoundKeyOutput[9]), .ZN(\SubCellInst_LFInst_2_LFInst_1_n10 ) );
  INV_X1 \SubCellInst_LFInst_2_LFInst_1_U3  ( .A(AddRoundKeyOutput[10]), .ZN(
        \SubCellInst_LFInst_2_LFInst_1_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_2_LFInst_2_U11  ( .A1(
        \SubCellInst_LFInst_2_LFInst_2_n22 ), .A2(
        \SubCellInst_LFInst_2_LFInst_2_n21 ), .ZN(\MCInst_MC2_v3_0 [3]) );
  NAND2_X1 \SubCellInst_LFInst_2_LFInst_2_U10  ( .A1(AddRoundKeyOutput[10]), 
        .A2(\SubCellInst_LFInst_2_LFInst_2_n20 ), .ZN(
        \SubCellInst_LFInst_2_LFInst_2_n21 ) );
  NOR2_X1 \SubCellInst_LFInst_2_LFInst_2_U9  ( .A1(AddRoundKeyOutput[9]), .A2(
        \SubCellInst_LFInst_2_LFInst_2_n19 ), .ZN(
        \SubCellInst_LFInst_2_LFInst_2_n20 ) );
  INV_X1 \SubCellInst_LFInst_2_LFInst_2_U8  ( .A(AddRoundKeyOutput[11]), .ZN(
        \SubCellInst_LFInst_2_LFInst_2_n19 ) );
  NAND2_X1 \SubCellInst_LFInst_2_LFInst_2_U7  ( .A1(
        \SubCellInst_LFInst_2_LFInst_2_n18 ), .A2(
        \SubCellInst_LFInst_2_LFInst_2_n17 ), .ZN(
        \SubCellInst_LFInst_2_LFInst_2_n22 ) );
  XOR2_X1 \SubCellInst_LFInst_2_LFInst_2_U6  ( .A(
        \SubCellInst_LFInst_2_LFInst_2_n16 ), .B(AddRoundKeyOutput[10]), .Z(
        \SubCellInst_LFInst_2_LFInst_2_n17 ) );
  NAND2_X1 \SubCellInst_LFInst_2_LFInst_2_U5  ( .A1(AddRoundKeyOutput[8]), 
        .A2(AddRoundKeyOutput[9]), .ZN(\SubCellInst_LFInst_2_LFInst_2_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_2_LFInst_2_U4  ( .A1(
        \SubCellInst_LFInst_2_LFInst_2_n15 ), .A2(AddRoundKeyOutput[11]), .ZN(
        \SubCellInst_LFInst_2_LFInst_2_n18 ) );
  XNOR2_X1 \SubCellInst_LFInst_2_LFInst_2_U3  ( .A(AddRoundKeyOutput[8]), .B(
        AddRoundKeyOutput[9]), .ZN(\SubCellInst_LFInst_2_LFInst_2_n15 ) );
  NAND2_X1 \SubCellInst_LFInst_2_LFInst_3_U9  ( .A1(
        \SubCellInst_LFInst_2_LFInst_3_n16 ), .A2(
        \SubCellInst_LFInst_2_LFInst_3_n15 ), .ZN(\Red_MCInst_MC2_v3_1 [2]) );
  NAND2_X1 \SubCellInst_LFInst_2_LFInst_3_U8  ( .A1(AddRoundKeyOutput[9]), 
        .A2(\SubCellInst_LFInst_2_LFInst_3_n14 ), .ZN(
        \SubCellInst_LFInst_2_LFInst_3_n15 ) );
  XOR2_X1 \SubCellInst_LFInst_2_LFInst_3_U7  ( .A(AddRoundKeyOutput[11]), .B(
        AddRoundKeyOutput[10]), .Z(\SubCellInst_LFInst_2_LFInst_3_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_2_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_2_LFInst_3_n13 ), .A2(
        \SubCellInst_LFInst_2_LFInst_3_n12 ), .ZN(
        \SubCellInst_LFInst_2_LFInst_3_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_2_LFInst_3_U5  ( .A1(AddRoundKeyOutput[8]), 
        .A2(AddRoundKeyOutput[10]), .ZN(\SubCellInst_LFInst_2_LFInst_3_n12 )
         );
  XNOR2_X1 \SubCellInst_LFInst_2_LFInst_3_U4  ( .A(AddRoundKeyOutput[8]), .B(
        \SubCellInst_LFInst_2_LFInst_3_n11 ), .ZN(
        \SubCellInst_LFInst_2_LFInst_3_n13 ) );
  OR2_X1 \SubCellInst_LFInst_2_LFInst_3_U3  ( .A1(AddRoundKeyOutput[11]), .A2(
        AddRoundKeyOutput[9]), .ZN(\SubCellInst_LFInst_2_LFInst_3_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_3_LFInst_0_U7  ( .A1(AddRoundKeyOutput[14]), 
        .A2(\SubCellInst_LFInst_3_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_3_LFInst_0_n8 ) );
  INV_X1 \SubCellInst_LFInst_3_LFInst_0_U6  ( .A(AddRoundKeyOutput[13]), .ZN(
        \SubCellInst_LFInst_3_LFInst_0_n7 ) );
  XOR2_X1 \SubCellInst_LFInst_3_LFInst_0_U5  ( .A(AddRoundKeyOutput[12]), .B(
        AddRoundKeyOutput[15]), .Z(\SubCellInst_LFInst_3_LFInst_0_n9 ) );
  INV_X1 \SubCellInst_LFInst_3_LFInst_0_U4  ( .A(
        \SubCellInst_LFInst_3_LFInst_0_n10 ), .ZN(\MCInst_MC1_v3_2 [3]) );
  XOR2_X1 \SubCellInst_LFInst_3_LFInst_0_U3  ( .A(
        \SubCellInst_LFInst_3_LFInst_0_n9 ), .B(
        \SubCellInst_LFInst_3_LFInst_0_n8 ), .Z(
        \SubCellInst_LFInst_3_LFInst_0_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_3_LFInst_1_U12  ( .A1(
        \SubCellInst_LFInst_3_LFInst_1_n18 ), .A2(
        \SubCellInst_LFInst_3_LFInst_1_n17 ), .ZN(\Red_MCInst_MC1_v3_3 [2]) );
  NAND2_X1 \SubCellInst_LFInst_3_LFInst_1_U11  ( .A1(AddRoundKeyOutput[13]), 
        .A2(\SubCellInst_LFInst_3_LFInst_1_n16 ), .ZN(
        \SubCellInst_LFInst_3_LFInst_1_n17 ) );
  NOR2_X1 \SubCellInst_LFInst_3_LFInst_1_U10  ( .A1(AddRoundKeyOutput[15]), 
        .A2(\SubCellInst_LFInst_3_LFInst_1_n15 ), .ZN(
        \SubCellInst_LFInst_3_LFInst_1_n16 ) );
  AND2_X1 \SubCellInst_LFInst_3_LFInst_1_U9  ( .A1(AddRoundKeyOutput[12]), 
        .A2(AddRoundKeyOutput[14]), .ZN(\SubCellInst_LFInst_3_LFInst_1_n15 )
         );
  NAND2_X1 \SubCellInst_LFInst_3_LFInst_1_U8  ( .A1(AddRoundKeyOutput[15]), 
        .A2(\SubCellInst_LFInst_3_LFInst_1_n14 ), .ZN(
        \SubCellInst_LFInst_3_LFInst_1_n18 ) );
  NAND2_X1 \SubCellInst_LFInst_3_LFInst_1_U7  ( .A1(
        \SubCellInst_LFInst_3_LFInst_1_n13 ), .A2(
        \SubCellInst_LFInst_3_LFInst_1_n12 ), .ZN(
        \SubCellInst_LFInst_3_LFInst_1_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_3_LFInst_1_U6  ( .A1(AddRoundKeyOutput[12]), 
        .A2(AddRoundKeyOutput[14]), .ZN(\SubCellInst_LFInst_3_LFInst_1_n12 )
         );
  NAND2_X1 \SubCellInst_LFInst_3_LFInst_1_U5  ( .A1(
        \SubCellInst_LFInst_3_LFInst_1_n11 ), .A2(
        \SubCellInst_LFInst_3_LFInst_1_n10 ), .ZN(
        \SubCellInst_LFInst_3_LFInst_1_n13 ) );
  NAND2_X1 \SubCellInst_LFInst_3_LFInst_1_U4  ( .A1(AddRoundKeyOutput[12]), 
        .A2(AddRoundKeyOutput[13]), .ZN(\SubCellInst_LFInst_3_LFInst_1_n10 )
         );
  INV_X1 \SubCellInst_LFInst_3_LFInst_1_U3  ( .A(AddRoundKeyOutput[14]), .ZN(
        \SubCellInst_LFInst_3_LFInst_1_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_3_LFInst_2_U11  ( .A1(
        \SubCellInst_LFInst_3_LFInst_2_n22 ), .A2(
        \SubCellInst_LFInst_3_LFInst_2_n21 ), .ZN(\MCInst_MC1_v3_0 [3]) );
  NAND2_X1 \SubCellInst_LFInst_3_LFInst_2_U10  ( .A1(AddRoundKeyOutput[14]), 
        .A2(\SubCellInst_LFInst_3_LFInst_2_n20 ), .ZN(
        \SubCellInst_LFInst_3_LFInst_2_n21 ) );
  NOR2_X1 \SubCellInst_LFInst_3_LFInst_2_U9  ( .A1(AddRoundKeyOutput[13]), 
        .A2(\SubCellInst_LFInst_3_LFInst_2_n19 ), .ZN(
        \SubCellInst_LFInst_3_LFInst_2_n20 ) );
  INV_X1 \SubCellInst_LFInst_3_LFInst_2_U8  ( .A(AddRoundKeyOutput[15]), .ZN(
        \SubCellInst_LFInst_3_LFInst_2_n19 ) );
  NAND2_X1 \SubCellInst_LFInst_3_LFInst_2_U7  ( .A1(
        \SubCellInst_LFInst_3_LFInst_2_n18 ), .A2(
        \SubCellInst_LFInst_3_LFInst_2_n17 ), .ZN(
        \SubCellInst_LFInst_3_LFInst_2_n22 ) );
  XOR2_X1 \SubCellInst_LFInst_3_LFInst_2_U6  ( .A(
        \SubCellInst_LFInst_3_LFInst_2_n16 ), .B(AddRoundKeyOutput[14]), .Z(
        \SubCellInst_LFInst_3_LFInst_2_n17 ) );
  NAND2_X1 \SubCellInst_LFInst_3_LFInst_2_U5  ( .A1(AddRoundKeyOutput[12]), 
        .A2(AddRoundKeyOutput[13]), .ZN(\SubCellInst_LFInst_3_LFInst_2_n16 )
         );
  NAND2_X1 \SubCellInst_LFInst_3_LFInst_2_U4  ( .A1(
        \SubCellInst_LFInst_3_LFInst_2_n15 ), .A2(AddRoundKeyOutput[15]), .ZN(
        \SubCellInst_LFInst_3_LFInst_2_n18 ) );
  XNOR2_X1 \SubCellInst_LFInst_3_LFInst_2_U3  ( .A(AddRoundKeyOutput[12]), .B(
        AddRoundKeyOutput[13]), .ZN(\SubCellInst_LFInst_3_LFInst_2_n15 ) );
  NAND2_X1 \SubCellInst_LFInst_3_LFInst_3_U9  ( .A1(
        \SubCellInst_LFInst_3_LFInst_3_n16 ), .A2(
        \SubCellInst_LFInst_3_LFInst_3_n15 ), .ZN(\Red_MCInst_MC1_v3_1 [2]) );
  NAND2_X1 \SubCellInst_LFInst_3_LFInst_3_U8  ( .A1(AddRoundKeyOutput[13]), 
        .A2(\SubCellInst_LFInst_3_LFInst_3_n14 ), .ZN(
        \SubCellInst_LFInst_3_LFInst_3_n15 ) );
  XOR2_X1 \SubCellInst_LFInst_3_LFInst_3_U7  ( .A(AddRoundKeyOutput[15]), .B(
        AddRoundKeyOutput[14]), .Z(\SubCellInst_LFInst_3_LFInst_3_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_3_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_3_LFInst_3_n13 ), .A2(
        \SubCellInst_LFInst_3_LFInst_3_n12 ), .ZN(
        \SubCellInst_LFInst_3_LFInst_3_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_3_LFInst_3_U5  ( .A1(AddRoundKeyOutput[12]), 
        .A2(AddRoundKeyOutput[14]), .ZN(\SubCellInst_LFInst_3_LFInst_3_n12 )
         );
  XNOR2_X1 \SubCellInst_LFInst_3_LFInst_3_U4  ( .A(AddRoundKeyOutput[12]), .B(
        \SubCellInst_LFInst_3_LFInst_3_n11 ), .ZN(
        \SubCellInst_LFInst_3_LFInst_3_n13 ) );
  OR2_X1 \SubCellInst_LFInst_3_LFInst_3_U3  ( .A1(AddRoundKeyOutput[15]), .A2(
        AddRoundKeyOutput[13]), .ZN(\SubCellInst_LFInst_3_LFInst_3_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_4_LFInst_0_U7  ( .A1(AddRoundKeyOutput[18]), 
        .A2(\SubCellInst_LFInst_4_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_4_LFInst_0_n8 ) );
  INV_X1 \SubCellInst_LFInst_4_LFInst_0_U6  ( .A(AddRoundKeyOutput[17]), .ZN(
        \SubCellInst_LFInst_4_LFInst_0_n7 ) );
  XOR2_X1 \SubCellInst_LFInst_4_LFInst_0_U5  ( .A(AddRoundKeyOutput[16]), .B(
        AddRoundKeyOutput[19]), .Z(\SubCellInst_LFInst_4_LFInst_0_n9 ) );
  INV_X2 \SubCellInst_LFInst_4_LFInst_0_U4  ( .A(
        \SubCellInst_LFInst_4_LFInst_0_n10 ), .ZN(\Red_MCInst_MC1_v2_1 [1]) );
  XOR2_X1 \SubCellInst_LFInst_4_LFInst_0_U3  ( .A(
        \SubCellInst_LFInst_4_LFInst_0_n9 ), .B(
        \SubCellInst_LFInst_4_LFInst_0_n8 ), .Z(
        \SubCellInst_LFInst_4_LFInst_0_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_4_LFInst_1_U12  ( .A1(
        \SubCellInst_LFInst_4_LFInst_1_n18 ), .A2(
        \SubCellInst_LFInst_4_LFInst_1_n17 ), .ZN(\MCInst_MC1_v2_0 [2]) );
  NAND2_X1 \SubCellInst_LFInst_4_LFInst_1_U11  ( .A1(AddRoundKeyOutput[17]), 
        .A2(\SubCellInst_LFInst_4_LFInst_1_n16 ), .ZN(
        \SubCellInst_LFInst_4_LFInst_1_n17 ) );
  NOR2_X1 \SubCellInst_LFInst_4_LFInst_1_U10  ( .A1(AddRoundKeyOutput[19]), 
        .A2(\SubCellInst_LFInst_4_LFInst_1_n15 ), .ZN(
        \SubCellInst_LFInst_4_LFInst_1_n16 ) );
  AND2_X1 \SubCellInst_LFInst_4_LFInst_1_U9  ( .A1(AddRoundKeyOutput[16]), 
        .A2(AddRoundKeyOutput[18]), .ZN(\SubCellInst_LFInst_4_LFInst_1_n15 )
         );
  NAND2_X1 \SubCellInst_LFInst_4_LFInst_1_U8  ( .A1(AddRoundKeyOutput[19]), 
        .A2(\SubCellInst_LFInst_4_LFInst_1_n14 ), .ZN(
        \SubCellInst_LFInst_4_LFInst_1_n18 ) );
  NAND2_X1 \SubCellInst_LFInst_4_LFInst_1_U7  ( .A1(
        \SubCellInst_LFInst_4_LFInst_1_n13 ), .A2(
        \SubCellInst_LFInst_4_LFInst_1_n12 ), .ZN(
        \SubCellInst_LFInst_4_LFInst_1_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_4_LFInst_1_U6  ( .A1(AddRoundKeyOutput[16]), 
        .A2(AddRoundKeyOutput[18]), .ZN(\SubCellInst_LFInst_4_LFInst_1_n12 )
         );
  NAND2_X1 \SubCellInst_LFInst_4_LFInst_1_U5  ( .A1(
        \SubCellInst_LFInst_4_LFInst_1_n11 ), .A2(
        \SubCellInst_LFInst_4_LFInst_1_n10 ), .ZN(
        \SubCellInst_LFInst_4_LFInst_1_n13 ) );
  NAND2_X1 \SubCellInst_LFInst_4_LFInst_1_U4  ( .A1(AddRoundKeyOutput[16]), 
        .A2(AddRoundKeyOutput[17]), .ZN(\SubCellInst_LFInst_4_LFInst_1_n10 )
         );
  INV_X1 \SubCellInst_LFInst_4_LFInst_1_U3  ( .A(AddRoundKeyOutput[18]), .ZN(
        \SubCellInst_LFInst_4_LFInst_1_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_4_LFInst_2_U11  ( .A1(
        \SubCellInst_LFInst_4_LFInst_2_n22 ), .A2(
        \SubCellInst_LFInst_4_LFInst_2_n21 ), .ZN(\MCInst_MC1_v2_0 [3]) );
  NAND2_X1 \SubCellInst_LFInst_4_LFInst_2_U10  ( .A1(AddRoundKeyOutput[18]), 
        .A2(\SubCellInst_LFInst_4_LFInst_2_n20 ), .ZN(
        \SubCellInst_LFInst_4_LFInst_2_n21 ) );
  NOR2_X1 \SubCellInst_LFInst_4_LFInst_2_U9  ( .A1(AddRoundKeyOutput[17]), 
        .A2(\SubCellInst_LFInst_4_LFInst_2_n19 ), .ZN(
        \SubCellInst_LFInst_4_LFInst_2_n20 ) );
  INV_X1 \SubCellInst_LFInst_4_LFInst_2_U8  ( .A(AddRoundKeyOutput[19]), .ZN(
        \SubCellInst_LFInst_4_LFInst_2_n19 ) );
  NAND2_X1 \SubCellInst_LFInst_4_LFInst_2_U7  ( .A1(
        \SubCellInst_LFInst_4_LFInst_2_n18 ), .A2(
        \SubCellInst_LFInst_4_LFInst_2_n17 ), .ZN(
        \SubCellInst_LFInst_4_LFInst_2_n22 ) );
  XOR2_X1 \SubCellInst_LFInst_4_LFInst_2_U6  ( .A(
        \SubCellInst_LFInst_4_LFInst_2_n16 ), .B(AddRoundKeyOutput[18]), .Z(
        \SubCellInst_LFInst_4_LFInst_2_n17 ) );
  NAND2_X1 \SubCellInst_LFInst_4_LFInst_2_U5  ( .A1(AddRoundKeyOutput[16]), 
        .A2(AddRoundKeyOutput[17]), .ZN(\SubCellInst_LFInst_4_LFInst_2_n16 )
         );
  NAND2_X1 \SubCellInst_LFInst_4_LFInst_2_U4  ( .A1(
        \SubCellInst_LFInst_4_LFInst_2_n15 ), .A2(AddRoundKeyOutput[19]), .ZN(
        \SubCellInst_LFInst_4_LFInst_2_n18 ) );
  XNOR2_X1 \SubCellInst_LFInst_4_LFInst_2_U3  ( .A(AddRoundKeyOutput[16]), .B(
        AddRoundKeyOutput[17]), .ZN(\SubCellInst_LFInst_4_LFInst_2_n15 ) );
  NAND2_X1 \SubCellInst_LFInst_4_LFInst_3_U9  ( .A1(AddRoundKeyOutput[17]), 
        .A2(\SubCellInst_LFInst_4_LFInst_3_n14 ), .ZN(
        \SubCellInst_LFInst_4_LFInst_3_n15 ) );
  XOR2_X1 \SubCellInst_LFInst_4_LFInst_3_U8  ( .A(AddRoundKeyOutput[19]), .B(
        AddRoundKeyOutput[18]), .Z(\SubCellInst_LFInst_4_LFInst_3_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_4_LFInst_3_U7  ( .A1(
        \SubCellInst_LFInst_4_LFInst_3_n13 ), .A2(
        \SubCellInst_LFInst_4_LFInst_3_n12 ), .ZN(
        \SubCellInst_LFInst_4_LFInst_3_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_4_LFInst_3_U6  ( .A1(AddRoundKeyOutput[16]), 
        .A2(AddRoundKeyOutput[18]), .ZN(\SubCellInst_LFInst_4_LFInst_3_n12 )
         );
  XNOR2_X1 \SubCellInst_LFInst_4_LFInst_3_U5  ( .A(AddRoundKeyOutput[16]), .B(
        \SubCellInst_LFInst_4_LFInst_3_n11 ), .ZN(
        \SubCellInst_LFInst_4_LFInst_3_n13 ) );
  OR2_X1 \SubCellInst_LFInst_4_LFInst_3_U4  ( .A1(AddRoundKeyOutput[19]), .A2(
        AddRoundKeyOutput[17]), .ZN(\SubCellInst_LFInst_4_LFInst_3_n11 ) );
  NAND2_X2 \SubCellInst_LFInst_4_LFInst_3_U3  ( .A1(
        \SubCellInst_LFInst_4_LFInst_3_n16 ), .A2(
        \SubCellInst_LFInst_4_LFInst_3_n15 ), .ZN(\Red_MCInst_MC1_v2_2 [1]) );
  NAND2_X1 \SubCellInst_LFInst_5_LFInst_0_U7  ( .A1(AddRoundKeyOutput[22]), 
        .A2(\SubCellInst_LFInst_5_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_5_LFInst_0_n8 ) );
  INV_X1 \SubCellInst_LFInst_5_LFInst_0_U6  ( .A(AddRoundKeyOutput[21]), .ZN(
        \SubCellInst_LFInst_5_LFInst_0_n7 ) );
  XOR2_X1 \SubCellInst_LFInst_5_LFInst_0_U5  ( .A(AddRoundKeyOutput[20]), .B(
        AddRoundKeyOutput[23]), .Z(\SubCellInst_LFInst_5_LFInst_0_n9 ) );
  INV_X2 \SubCellInst_LFInst_5_LFInst_0_U4  ( .A(
        \SubCellInst_LFInst_5_LFInst_0_n10 ), .ZN(\Red_MCInst_MC0_v2_1 [1]) );
  XOR2_X1 \SubCellInst_LFInst_5_LFInst_0_U3  ( .A(
        \SubCellInst_LFInst_5_LFInst_0_n9 ), .B(
        \SubCellInst_LFInst_5_LFInst_0_n8 ), .Z(
        \SubCellInst_LFInst_5_LFInst_0_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_5_LFInst_1_U12  ( .A1(
        \SubCellInst_LFInst_5_LFInst_1_n18 ), .A2(
        \SubCellInst_LFInst_5_LFInst_1_n17 ), .ZN(\MCInst_MC0_v2_0 [2]) );
  NAND2_X1 \SubCellInst_LFInst_5_LFInst_1_U11  ( .A1(AddRoundKeyOutput[21]), 
        .A2(\SubCellInst_LFInst_5_LFInst_1_n16 ), .ZN(
        \SubCellInst_LFInst_5_LFInst_1_n17 ) );
  NOR2_X1 \SubCellInst_LFInst_5_LFInst_1_U10  ( .A1(AddRoundKeyOutput[23]), 
        .A2(\SubCellInst_LFInst_5_LFInst_1_n15 ), .ZN(
        \SubCellInst_LFInst_5_LFInst_1_n16 ) );
  AND2_X1 \SubCellInst_LFInst_5_LFInst_1_U9  ( .A1(AddRoundKeyOutput[20]), 
        .A2(AddRoundKeyOutput[22]), .ZN(\SubCellInst_LFInst_5_LFInst_1_n15 )
         );
  NAND2_X1 \SubCellInst_LFInst_5_LFInst_1_U8  ( .A1(AddRoundKeyOutput[23]), 
        .A2(\SubCellInst_LFInst_5_LFInst_1_n14 ), .ZN(
        \SubCellInst_LFInst_5_LFInst_1_n18 ) );
  NAND2_X1 \SubCellInst_LFInst_5_LFInst_1_U7  ( .A1(
        \SubCellInst_LFInst_5_LFInst_1_n13 ), .A2(
        \SubCellInst_LFInst_5_LFInst_1_n12 ), .ZN(
        \SubCellInst_LFInst_5_LFInst_1_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_5_LFInst_1_U6  ( .A1(AddRoundKeyOutput[20]), 
        .A2(AddRoundKeyOutput[22]), .ZN(\SubCellInst_LFInst_5_LFInst_1_n12 )
         );
  NAND2_X1 \SubCellInst_LFInst_5_LFInst_1_U5  ( .A1(
        \SubCellInst_LFInst_5_LFInst_1_n11 ), .A2(
        \SubCellInst_LFInst_5_LFInst_1_n10 ), .ZN(
        \SubCellInst_LFInst_5_LFInst_1_n13 ) );
  NAND2_X1 \SubCellInst_LFInst_5_LFInst_1_U4  ( .A1(AddRoundKeyOutput[20]), 
        .A2(AddRoundKeyOutput[21]), .ZN(\SubCellInst_LFInst_5_LFInst_1_n10 )
         );
  INV_X1 \SubCellInst_LFInst_5_LFInst_1_U3  ( .A(AddRoundKeyOutput[22]), .ZN(
        \SubCellInst_LFInst_5_LFInst_1_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_5_LFInst_2_U11  ( .A1(
        \SubCellInst_LFInst_5_LFInst_2_n22 ), .A2(
        \SubCellInst_LFInst_5_LFInst_2_n21 ), .ZN(\MCInst_MC0_v2_0 [3]) );
  NAND2_X1 \SubCellInst_LFInst_5_LFInst_2_U10  ( .A1(AddRoundKeyOutput[22]), 
        .A2(\SubCellInst_LFInst_5_LFInst_2_n20 ), .ZN(
        \SubCellInst_LFInst_5_LFInst_2_n21 ) );
  NOR2_X1 \SubCellInst_LFInst_5_LFInst_2_U9  ( .A1(AddRoundKeyOutput[21]), 
        .A2(\SubCellInst_LFInst_5_LFInst_2_n19 ), .ZN(
        \SubCellInst_LFInst_5_LFInst_2_n20 ) );
  INV_X1 \SubCellInst_LFInst_5_LFInst_2_U8  ( .A(AddRoundKeyOutput[23]), .ZN(
        \SubCellInst_LFInst_5_LFInst_2_n19 ) );
  NAND2_X1 \SubCellInst_LFInst_5_LFInst_2_U7  ( .A1(
        \SubCellInst_LFInst_5_LFInst_2_n18 ), .A2(
        \SubCellInst_LFInst_5_LFInst_2_n17 ), .ZN(
        \SubCellInst_LFInst_5_LFInst_2_n22 ) );
  XOR2_X1 \SubCellInst_LFInst_5_LFInst_2_U6  ( .A(
        \SubCellInst_LFInst_5_LFInst_2_n16 ), .B(AddRoundKeyOutput[22]), .Z(
        \SubCellInst_LFInst_5_LFInst_2_n17 ) );
  NAND2_X1 \SubCellInst_LFInst_5_LFInst_2_U5  ( .A1(AddRoundKeyOutput[20]), 
        .A2(AddRoundKeyOutput[21]), .ZN(\SubCellInst_LFInst_5_LFInst_2_n16 )
         );
  NAND2_X1 \SubCellInst_LFInst_5_LFInst_2_U4  ( .A1(
        \SubCellInst_LFInst_5_LFInst_2_n15 ), .A2(AddRoundKeyOutput[23]), .ZN(
        \SubCellInst_LFInst_5_LFInst_2_n18 ) );
  XNOR2_X1 \SubCellInst_LFInst_5_LFInst_2_U3  ( .A(AddRoundKeyOutput[20]), .B(
        AddRoundKeyOutput[21]), .ZN(\SubCellInst_LFInst_5_LFInst_2_n15 ) );
  NAND2_X1 \SubCellInst_LFInst_5_LFInst_3_U9  ( .A1(AddRoundKeyOutput[21]), 
        .A2(\SubCellInst_LFInst_5_LFInst_3_n14 ), .ZN(
        \SubCellInst_LFInst_5_LFInst_3_n15 ) );
  XOR2_X1 \SubCellInst_LFInst_5_LFInst_3_U8  ( .A(AddRoundKeyOutput[23]), .B(
        AddRoundKeyOutput[22]), .Z(\SubCellInst_LFInst_5_LFInst_3_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_5_LFInst_3_U7  ( .A1(
        \SubCellInst_LFInst_5_LFInst_3_n13 ), .A2(
        \SubCellInst_LFInst_5_LFInst_3_n12 ), .ZN(
        \SubCellInst_LFInst_5_LFInst_3_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_5_LFInst_3_U6  ( .A1(AddRoundKeyOutput[20]), 
        .A2(AddRoundKeyOutput[22]), .ZN(\SubCellInst_LFInst_5_LFInst_3_n12 )
         );
  XNOR2_X1 \SubCellInst_LFInst_5_LFInst_3_U5  ( .A(AddRoundKeyOutput[20]), .B(
        \SubCellInst_LFInst_5_LFInst_3_n11 ), .ZN(
        \SubCellInst_LFInst_5_LFInst_3_n13 ) );
  OR2_X1 \SubCellInst_LFInst_5_LFInst_3_U4  ( .A1(AddRoundKeyOutput[23]), .A2(
        AddRoundKeyOutput[21]), .ZN(\SubCellInst_LFInst_5_LFInst_3_n11 ) );
  NAND2_X2 \SubCellInst_LFInst_5_LFInst_3_U3  ( .A1(
        \SubCellInst_LFInst_5_LFInst_3_n16 ), .A2(
        \SubCellInst_LFInst_5_LFInst_3_n15 ), .ZN(\Red_MCInst_MC0_v2_2 [1]) );
  NAND2_X1 \SubCellInst_LFInst_6_LFInst_0_U7  ( .A1(AddRoundKeyOutput[26]), 
        .A2(\SubCellInst_LFInst_6_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_6_LFInst_0_n8 ) );
  INV_X1 \SubCellInst_LFInst_6_LFInst_0_U6  ( .A(AddRoundKeyOutput[25]), .ZN(
        \SubCellInst_LFInst_6_LFInst_0_n7 ) );
  XOR2_X1 \SubCellInst_LFInst_6_LFInst_0_U5  ( .A(AddRoundKeyOutput[24]), .B(
        AddRoundKeyOutput[27]), .Z(\SubCellInst_LFInst_6_LFInst_0_n9 ) );
  INV_X2 \SubCellInst_LFInst_6_LFInst_0_U4  ( .A(
        \SubCellInst_LFInst_6_LFInst_0_n10 ), .ZN(\Red_MCInst_MC3_v2_1 [1]) );
  XOR2_X1 \SubCellInst_LFInst_6_LFInst_0_U3  ( .A(
        \SubCellInst_LFInst_6_LFInst_0_n9 ), .B(
        \SubCellInst_LFInst_6_LFInst_0_n8 ), .Z(
        \SubCellInst_LFInst_6_LFInst_0_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_6_LFInst_1_U12  ( .A1(
        \SubCellInst_LFInst_6_LFInst_1_n18 ), .A2(
        \SubCellInst_LFInst_6_LFInst_1_n17 ), .ZN(\MCInst_MC3_v2_0 [2]) );
  NAND2_X1 \SubCellInst_LFInst_6_LFInst_1_U11  ( .A1(AddRoundKeyOutput[25]), 
        .A2(\SubCellInst_LFInst_6_LFInst_1_n16 ), .ZN(
        \SubCellInst_LFInst_6_LFInst_1_n17 ) );
  NOR2_X1 \SubCellInst_LFInst_6_LFInst_1_U10  ( .A1(AddRoundKeyOutput[27]), 
        .A2(\SubCellInst_LFInst_6_LFInst_1_n15 ), .ZN(
        \SubCellInst_LFInst_6_LFInst_1_n16 ) );
  AND2_X1 \SubCellInst_LFInst_6_LFInst_1_U9  ( .A1(AddRoundKeyOutput[24]), 
        .A2(AddRoundKeyOutput[26]), .ZN(\SubCellInst_LFInst_6_LFInst_1_n15 )
         );
  NAND2_X1 \SubCellInst_LFInst_6_LFInst_1_U8  ( .A1(AddRoundKeyOutput[27]), 
        .A2(\SubCellInst_LFInst_6_LFInst_1_n14 ), .ZN(
        \SubCellInst_LFInst_6_LFInst_1_n18 ) );
  NAND2_X1 \SubCellInst_LFInst_6_LFInst_1_U7  ( .A1(
        \SubCellInst_LFInst_6_LFInst_1_n13 ), .A2(
        \SubCellInst_LFInst_6_LFInst_1_n12 ), .ZN(
        \SubCellInst_LFInst_6_LFInst_1_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_6_LFInst_1_U6  ( .A1(AddRoundKeyOutput[24]), 
        .A2(AddRoundKeyOutput[26]), .ZN(\SubCellInst_LFInst_6_LFInst_1_n12 )
         );
  NAND2_X1 \SubCellInst_LFInst_6_LFInst_1_U5  ( .A1(
        \SubCellInst_LFInst_6_LFInst_1_n11 ), .A2(
        \SubCellInst_LFInst_6_LFInst_1_n10 ), .ZN(
        \SubCellInst_LFInst_6_LFInst_1_n13 ) );
  NAND2_X1 \SubCellInst_LFInst_6_LFInst_1_U4  ( .A1(AddRoundKeyOutput[24]), 
        .A2(AddRoundKeyOutput[25]), .ZN(\SubCellInst_LFInst_6_LFInst_1_n10 )
         );
  INV_X1 \SubCellInst_LFInst_6_LFInst_1_U3  ( .A(AddRoundKeyOutput[26]), .ZN(
        \SubCellInst_LFInst_6_LFInst_1_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_6_LFInst_2_U11  ( .A1(
        \SubCellInst_LFInst_6_LFInst_2_n22 ), .A2(
        \SubCellInst_LFInst_6_LFInst_2_n21 ), .ZN(\MCInst_MC3_v2_0 [3]) );
  NAND2_X1 \SubCellInst_LFInst_6_LFInst_2_U10  ( .A1(AddRoundKeyOutput[26]), 
        .A2(\SubCellInst_LFInst_6_LFInst_2_n20 ), .ZN(
        \SubCellInst_LFInst_6_LFInst_2_n21 ) );
  NOR2_X1 \SubCellInst_LFInst_6_LFInst_2_U9  ( .A1(AddRoundKeyOutput[25]), 
        .A2(\SubCellInst_LFInst_6_LFInst_2_n19 ), .ZN(
        \SubCellInst_LFInst_6_LFInst_2_n20 ) );
  INV_X1 \SubCellInst_LFInst_6_LFInst_2_U8  ( .A(AddRoundKeyOutput[27]), .ZN(
        \SubCellInst_LFInst_6_LFInst_2_n19 ) );
  NAND2_X1 \SubCellInst_LFInst_6_LFInst_2_U7  ( .A1(
        \SubCellInst_LFInst_6_LFInst_2_n18 ), .A2(
        \SubCellInst_LFInst_6_LFInst_2_n17 ), .ZN(
        \SubCellInst_LFInst_6_LFInst_2_n22 ) );
  XOR2_X1 \SubCellInst_LFInst_6_LFInst_2_U6  ( .A(
        \SubCellInst_LFInst_6_LFInst_2_n16 ), .B(AddRoundKeyOutput[26]), .Z(
        \SubCellInst_LFInst_6_LFInst_2_n17 ) );
  NAND2_X1 \SubCellInst_LFInst_6_LFInst_2_U5  ( .A1(AddRoundKeyOutput[24]), 
        .A2(AddRoundKeyOutput[25]), .ZN(\SubCellInst_LFInst_6_LFInst_2_n16 )
         );
  NAND2_X1 \SubCellInst_LFInst_6_LFInst_2_U4  ( .A1(
        \SubCellInst_LFInst_6_LFInst_2_n15 ), .A2(AddRoundKeyOutput[27]), .ZN(
        \SubCellInst_LFInst_6_LFInst_2_n18 ) );
  XNOR2_X1 \SubCellInst_LFInst_6_LFInst_2_U3  ( .A(AddRoundKeyOutput[24]), .B(
        AddRoundKeyOutput[25]), .ZN(\SubCellInst_LFInst_6_LFInst_2_n15 ) );
  NAND2_X1 \SubCellInst_LFInst_6_LFInst_3_U9  ( .A1(AddRoundKeyOutput[25]), 
        .A2(\SubCellInst_LFInst_6_LFInst_3_n14 ), .ZN(
        \SubCellInst_LFInst_6_LFInst_3_n15 ) );
  XOR2_X1 \SubCellInst_LFInst_6_LFInst_3_U8  ( .A(AddRoundKeyOutput[27]), .B(
        AddRoundKeyOutput[26]), .Z(\SubCellInst_LFInst_6_LFInst_3_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_6_LFInst_3_U7  ( .A1(
        \SubCellInst_LFInst_6_LFInst_3_n13 ), .A2(
        \SubCellInst_LFInst_6_LFInst_3_n12 ), .ZN(
        \SubCellInst_LFInst_6_LFInst_3_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_6_LFInst_3_U6  ( .A1(AddRoundKeyOutput[24]), 
        .A2(AddRoundKeyOutput[26]), .ZN(\SubCellInst_LFInst_6_LFInst_3_n12 )
         );
  XNOR2_X1 \SubCellInst_LFInst_6_LFInst_3_U5  ( .A(AddRoundKeyOutput[24]), .B(
        \SubCellInst_LFInst_6_LFInst_3_n11 ), .ZN(
        \SubCellInst_LFInst_6_LFInst_3_n13 ) );
  OR2_X1 \SubCellInst_LFInst_6_LFInst_3_U4  ( .A1(AddRoundKeyOutput[27]), .A2(
        AddRoundKeyOutput[25]), .ZN(\SubCellInst_LFInst_6_LFInst_3_n11 ) );
  NAND2_X2 \SubCellInst_LFInst_6_LFInst_3_U3  ( .A1(
        \SubCellInst_LFInst_6_LFInst_3_n16 ), .A2(
        \SubCellInst_LFInst_6_LFInst_3_n15 ), .ZN(\Red_MCInst_MC3_v2_2 [1]) );
  NAND2_X1 \SubCellInst_LFInst_7_LFInst_0_U7  ( .A1(AddRoundKeyOutput[30]), 
        .A2(\SubCellInst_LFInst_7_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_7_LFInst_0_n8 ) );
  INV_X1 \SubCellInst_LFInst_7_LFInst_0_U6  ( .A(AddRoundKeyOutput[29]), .ZN(
        \SubCellInst_LFInst_7_LFInst_0_n7 ) );
  XOR2_X1 \SubCellInst_LFInst_7_LFInst_0_U5  ( .A(AddRoundKeyOutput[28]), .B(
        AddRoundKeyOutput[31]), .Z(\SubCellInst_LFInst_7_LFInst_0_n9 ) );
  INV_X2 \SubCellInst_LFInst_7_LFInst_0_U4  ( .A(
        \SubCellInst_LFInst_7_LFInst_0_n10 ), .ZN(\Red_MCInst_MC2_v2_1 [1]) );
  XOR2_X1 \SubCellInst_LFInst_7_LFInst_0_U3  ( .A(
        \SubCellInst_LFInst_7_LFInst_0_n9 ), .B(
        \SubCellInst_LFInst_7_LFInst_0_n8 ), .Z(
        \SubCellInst_LFInst_7_LFInst_0_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_7_LFInst_1_U12  ( .A1(
        \SubCellInst_LFInst_7_LFInst_1_n18 ), .A2(
        \SubCellInst_LFInst_7_LFInst_1_n17 ), .ZN(\MCInst_MC2_v2_0 [2]) );
  NAND2_X1 \SubCellInst_LFInst_7_LFInst_1_U11  ( .A1(AddRoundKeyOutput[29]), 
        .A2(\SubCellInst_LFInst_7_LFInst_1_n16 ), .ZN(
        \SubCellInst_LFInst_7_LFInst_1_n17 ) );
  NOR2_X1 \SubCellInst_LFInst_7_LFInst_1_U10  ( .A1(AddRoundKeyOutput[31]), 
        .A2(\SubCellInst_LFInst_7_LFInst_1_n15 ), .ZN(
        \SubCellInst_LFInst_7_LFInst_1_n16 ) );
  AND2_X1 \SubCellInst_LFInst_7_LFInst_1_U9  ( .A1(AddRoundKeyOutput[28]), 
        .A2(AddRoundKeyOutput[30]), .ZN(\SubCellInst_LFInst_7_LFInst_1_n15 )
         );
  NAND2_X1 \SubCellInst_LFInst_7_LFInst_1_U8  ( .A1(AddRoundKeyOutput[31]), 
        .A2(\SubCellInst_LFInst_7_LFInst_1_n14 ), .ZN(
        \SubCellInst_LFInst_7_LFInst_1_n18 ) );
  NAND2_X1 \SubCellInst_LFInst_7_LFInst_1_U7  ( .A1(
        \SubCellInst_LFInst_7_LFInst_1_n13 ), .A2(
        \SubCellInst_LFInst_7_LFInst_1_n12 ), .ZN(
        \SubCellInst_LFInst_7_LFInst_1_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_7_LFInst_1_U6  ( .A1(AddRoundKeyOutput[28]), 
        .A2(AddRoundKeyOutput[30]), .ZN(\SubCellInst_LFInst_7_LFInst_1_n12 )
         );
  NAND2_X1 \SubCellInst_LFInst_7_LFInst_1_U5  ( .A1(
        \SubCellInst_LFInst_7_LFInst_1_n11 ), .A2(
        \SubCellInst_LFInst_7_LFInst_1_n10 ), .ZN(
        \SubCellInst_LFInst_7_LFInst_1_n13 ) );
  NAND2_X1 \SubCellInst_LFInst_7_LFInst_1_U4  ( .A1(AddRoundKeyOutput[28]), 
        .A2(AddRoundKeyOutput[29]), .ZN(\SubCellInst_LFInst_7_LFInst_1_n10 )
         );
  INV_X1 \SubCellInst_LFInst_7_LFInst_1_U3  ( .A(AddRoundKeyOutput[30]), .ZN(
        \SubCellInst_LFInst_7_LFInst_1_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_7_LFInst_2_U11  ( .A1(
        \SubCellInst_LFInst_7_LFInst_2_n22 ), .A2(
        \SubCellInst_LFInst_7_LFInst_2_n21 ), .ZN(\MCInst_MC2_v2_0 [3]) );
  NAND2_X1 \SubCellInst_LFInst_7_LFInst_2_U10  ( .A1(AddRoundKeyOutput[30]), 
        .A2(\SubCellInst_LFInst_7_LFInst_2_n20 ), .ZN(
        \SubCellInst_LFInst_7_LFInst_2_n21 ) );
  NOR2_X1 \SubCellInst_LFInst_7_LFInst_2_U9  ( .A1(AddRoundKeyOutput[29]), 
        .A2(\SubCellInst_LFInst_7_LFInst_2_n19 ), .ZN(
        \SubCellInst_LFInst_7_LFInst_2_n20 ) );
  INV_X1 \SubCellInst_LFInst_7_LFInst_2_U8  ( .A(AddRoundKeyOutput[31]), .ZN(
        \SubCellInst_LFInst_7_LFInst_2_n19 ) );
  NAND2_X1 \SubCellInst_LFInst_7_LFInst_2_U7  ( .A1(
        \SubCellInst_LFInst_7_LFInst_2_n18 ), .A2(
        \SubCellInst_LFInst_7_LFInst_2_n17 ), .ZN(
        \SubCellInst_LFInst_7_LFInst_2_n22 ) );
  XOR2_X1 \SubCellInst_LFInst_7_LFInst_2_U6  ( .A(
        \SubCellInst_LFInst_7_LFInst_2_n16 ), .B(AddRoundKeyOutput[30]), .Z(
        \SubCellInst_LFInst_7_LFInst_2_n17 ) );
  NAND2_X1 \SubCellInst_LFInst_7_LFInst_2_U5  ( .A1(AddRoundKeyOutput[28]), 
        .A2(AddRoundKeyOutput[29]), .ZN(\SubCellInst_LFInst_7_LFInst_2_n16 )
         );
  NAND2_X1 \SubCellInst_LFInst_7_LFInst_2_U4  ( .A1(
        \SubCellInst_LFInst_7_LFInst_2_n15 ), .A2(AddRoundKeyOutput[31]), .ZN(
        \SubCellInst_LFInst_7_LFInst_2_n18 ) );
  XNOR2_X1 \SubCellInst_LFInst_7_LFInst_2_U3  ( .A(AddRoundKeyOutput[28]), .B(
        AddRoundKeyOutput[29]), .ZN(\SubCellInst_LFInst_7_LFInst_2_n15 ) );
  NAND2_X1 \SubCellInst_LFInst_7_LFInst_3_U9  ( .A1(AddRoundKeyOutput[29]), 
        .A2(\SubCellInst_LFInst_7_LFInst_3_n14 ), .ZN(
        \SubCellInst_LFInst_7_LFInst_3_n15 ) );
  XOR2_X1 \SubCellInst_LFInst_7_LFInst_3_U8  ( .A(AddRoundKeyOutput[31]), .B(
        AddRoundKeyOutput[30]), .Z(\SubCellInst_LFInst_7_LFInst_3_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_7_LFInst_3_U7  ( .A1(
        \SubCellInst_LFInst_7_LFInst_3_n13 ), .A2(
        \SubCellInst_LFInst_7_LFInst_3_n12 ), .ZN(
        \SubCellInst_LFInst_7_LFInst_3_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_7_LFInst_3_U6  ( .A1(AddRoundKeyOutput[28]), 
        .A2(AddRoundKeyOutput[30]), .ZN(\SubCellInst_LFInst_7_LFInst_3_n12 )
         );
  XNOR2_X1 \SubCellInst_LFInst_7_LFInst_3_U5  ( .A(AddRoundKeyOutput[28]), .B(
        \SubCellInst_LFInst_7_LFInst_3_n11 ), .ZN(
        \SubCellInst_LFInst_7_LFInst_3_n13 ) );
  OR2_X1 \SubCellInst_LFInst_7_LFInst_3_U4  ( .A1(AddRoundKeyOutput[31]), .A2(
        AddRoundKeyOutput[29]), .ZN(\SubCellInst_LFInst_7_LFInst_3_n11 ) );
  NAND2_X2 \SubCellInst_LFInst_7_LFInst_3_U3  ( .A1(
        \SubCellInst_LFInst_7_LFInst_3_n16 ), .A2(
        \SubCellInst_LFInst_7_LFInst_3_n15 ), .ZN(\Red_MCInst_MC2_v2_2 [1]) );
  NAND2_X1 \SubCellInst_LFInst_8_LFInst_0_U7  ( .A1(AddRoundKeyOutput[34]), 
        .A2(\SubCellInst_LFInst_8_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_8_LFInst_0_n8 ) );
  INV_X1 \SubCellInst_LFInst_8_LFInst_0_U6  ( .A(AddRoundKeyOutput[33]), .ZN(
        \SubCellInst_LFInst_8_LFInst_0_n7 ) );
  XOR2_X1 \SubCellInst_LFInst_8_LFInst_0_U5  ( .A(AddRoundKeyOutput[32]), .B(
        AddRoundKeyOutput[35]), .Z(\SubCellInst_LFInst_8_LFInst_0_n9 ) );
  INV_X1 \SubCellInst_LFInst_8_LFInst_0_U4  ( .A(
        \SubCellInst_LFInst_8_LFInst_0_n10 ), .ZN(\MCInst_MC2_v1_0 [0]) );
  XOR2_X1 \SubCellInst_LFInst_8_LFInst_0_U3  ( .A(
        \SubCellInst_LFInst_8_LFInst_0_n9 ), .B(
        \SubCellInst_LFInst_8_LFInst_0_n8 ), .Z(
        \SubCellInst_LFInst_8_LFInst_0_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_8_LFInst_1_U12  ( .A1(AddRoundKeyOutput[33]), 
        .A2(\SubCellInst_LFInst_8_LFInst_1_n16 ), .ZN(
        \SubCellInst_LFInst_8_LFInst_1_n17 ) );
  NOR2_X1 \SubCellInst_LFInst_8_LFInst_1_U11  ( .A1(AddRoundKeyOutput[35]), 
        .A2(\SubCellInst_LFInst_8_LFInst_1_n15 ), .ZN(
        \SubCellInst_LFInst_8_LFInst_1_n16 ) );
  AND2_X1 \SubCellInst_LFInst_8_LFInst_1_U10  ( .A1(AddRoundKeyOutput[32]), 
        .A2(AddRoundKeyOutput[34]), .ZN(\SubCellInst_LFInst_8_LFInst_1_n15 )
         );
  NAND2_X1 \SubCellInst_LFInst_8_LFInst_1_U9  ( .A1(AddRoundKeyOutput[35]), 
        .A2(\SubCellInst_LFInst_8_LFInst_1_n14 ), .ZN(
        \SubCellInst_LFInst_8_LFInst_1_n18 ) );
  NAND2_X1 \SubCellInst_LFInst_8_LFInst_1_U8  ( .A1(
        \SubCellInst_LFInst_8_LFInst_1_n13 ), .A2(
        \SubCellInst_LFInst_8_LFInst_1_n12 ), .ZN(
        \SubCellInst_LFInst_8_LFInst_1_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_8_LFInst_1_U7  ( .A1(AddRoundKeyOutput[32]), 
        .A2(AddRoundKeyOutput[34]), .ZN(\SubCellInst_LFInst_8_LFInst_1_n12 )
         );
  NAND2_X1 \SubCellInst_LFInst_8_LFInst_1_U6  ( .A1(
        \SubCellInst_LFInst_8_LFInst_1_n11 ), .A2(
        \SubCellInst_LFInst_8_LFInst_1_n10 ), .ZN(
        \SubCellInst_LFInst_8_LFInst_1_n13 ) );
  NAND2_X1 \SubCellInst_LFInst_8_LFInst_1_U5  ( .A1(AddRoundKeyOutput[32]), 
        .A2(AddRoundKeyOutput[33]), .ZN(\SubCellInst_LFInst_8_LFInst_1_n10 )
         );
  INV_X1 \SubCellInst_LFInst_8_LFInst_1_U4  ( .A(AddRoundKeyOutput[34]), .ZN(
        \SubCellInst_LFInst_8_LFInst_1_n11 ) );
  NAND2_X2 \SubCellInst_LFInst_8_LFInst_1_U3  ( .A1(
        \SubCellInst_LFInst_8_LFInst_1_n18 ), .A2(
        \SubCellInst_LFInst_8_LFInst_1_n17 ), .ZN(\Red_MCInst_MC2_v1_2 [1]) );
  NAND2_X1 \SubCellInst_LFInst_8_LFInst_2_U11  ( .A1(
        \SubCellInst_LFInst_8_LFInst_2_n22 ), .A2(
        \SubCellInst_LFInst_8_LFInst_2_n21 ), .ZN(\MCInst_MC2_v1_3 [3]) );
  NAND2_X1 \SubCellInst_LFInst_8_LFInst_2_U10  ( .A1(AddRoundKeyOutput[34]), 
        .A2(\SubCellInst_LFInst_8_LFInst_2_n20 ), .ZN(
        \SubCellInst_LFInst_8_LFInst_2_n21 ) );
  NOR2_X1 \SubCellInst_LFInst_8_LFInst_2_U9  ( .A1(AddRoundKeyOutput[33]), 
        .A2(\SubCellInst_LFInst_8_LFInst_2_n19 ), .ZN(
        \SubCellInst_LFInst_8_LFInst_2_n20 ) );
  INV_X1 \SubCellInst_LFInst_8_LFInst_2_U8  ( .A(AddRoundKeyOutput[35]), .ZN(
        \SubCellInst_LFInst_8_LFInst_2_n19 ) );
  NAND2_X1 \SubCellInst_LFInst_8_LFInst_2_U7  ( .A1(
        \SubCellInst_LFInst_8_LFInst_2_n18 ), .A2(
        \SubCellInst_LFInst_8_LFInst_2_n17 ), .ZN(
        \SubCellInst_LFInst_8_LFInst_2_n22 ) );
  XOR2_X1 \SubCellInst_LFInst_8_LFInst_2_U6  ( .A(
        \SubCellInst_LFInst_8_LFInst_2_n16 ), .B(AddRoundKeyOutput[34]), .Z(
        \SubCellInst_LFInst_8_LFInst_2_n17 ) );
  NAND2_X1 \SubCellInst_LFInst_8_LFInst_2_U5  ( .A1(AddRoundKeyOutput[32]), 
        .A2(AddRoundKeyOutput[33]), .ZN(\SubCellInst_LFInst_8_LFInst_2_n16 )
         );
  NAND2_X1 \SubCellInst_LFInst_8_LFInst_2_U4  ( .A1(
        \SubCellInst_LFInst_8_LFInst_2_n15 ), .A2(AddRoundKeyOutput[35]), .ZN(
        \SubCellInst_LFInst_8_LFInst_2_n18 ) );
  XNOR2_X1 \SubCellInst_LFInst_8_LFInst_2_U3  ( .A(AddRoundKeyOutput[32]), .B(
        AddRoundKeyOutput[33]), .ZN(\SubCellInst_LFInst_8_LFInst_2_n15 ) );
  NAND2_X1 \SubCellInst_LFInst_8_LFInst_3_U9  ( .A1(
        \SubCellInst_LFInst_8_LFInst_3_n16 ), .A2(
        \SubCellInst_LFInst_8_LFInst_3_n15 ), .ZN(\Red_MCInst_MC2_v1_1 [2]) );
  NAND2_X1 \SubCellInst_LFInst_8_LFInst_3_U8  ( .A1(AddRoundKeyOutput[33]), 
        .A2(\SubCellInst_LFInst_8_LFInst_3_n14 ), .ZN(
        \SubCellInst_LFInst_8_LFInst_3_n15 ) );
  XOR2_X1 \SubCellInst_LFInst_8_LFInst_3_U7  ( .A(AddRoundKeyOutput[35]), .B(
        AddRoundKeyOutput[34]), .Z(\SubCellInst_LFInst_8_LFInst_3_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_8_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_8_LFInst_3_n13 ), .A2(
        \SubCellInst_LFInst_8_LFInst_3_n12 ), .ZN(
        \SubCellInst_LFInst_8_LFInst_3_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_8_LFInst_3_U5  ( .A1(AddRoundKeyOutput[32]), 
        .A2(AddRoundKeyOutput[34]), .ZN(\SubCellInst_LFInst_8_LFInst_3_n12 )
         );
  XNOR2_X1 \SubCellInst_LFInst_8_LFInst_3_U4  ( .A(AddRoundKeyOutput[32]), .B(
        \SubCellInst_LFInst_8_LFInst_3_n11 ), .ZN(
        \SubCellInst_LFInst_8_LFInst_3_n13 ) );
  OR2_X1 \SubCellInst_LFInst_8_LFInst_3_U3  ( .A1(AddRoundKeyOutput[35]), .A2(
        AddRoundKeyOutput[33]), .ZN(\SubCellInst_LFInst_8_LFInst_3_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_9_LFInst_0_U7  ( .A1(AddRoundKeyOutput[38]), 
        .A2(\SubCellInst_LFInst_9_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_9_LFInst_0_n8 ) );
  INV_X1 \SubCellInst_LFInst_9_LFInst_0_U6  ( .A(AddRoundKeyOutput[37]), .ZN(
        \SubCellInst_LFInst_9_LFInst_0_n7 ) );
  XOR2_X1 \SubCellInst_LFInst_9_LFInst_0_U5  ( .A(AddRoundKeyOutput[36]), .B(
        AddRoundKeyOutput[39]), .Z(\SubCellInst_LFInst_9_LFInst_0_n9 ) );
  INV_X1 \SubCellInst_LFInst_9_LFInst_0_U4  ( .A(
        \SubCellInst_LFInst_9_LFInst_0_n10 ), .ZN(\MCInst_MC1_v1_0 [0]) );
  XOR2_X1 \SubCellInst_LFInst_9_LFInst_0_U3  ( .A(
        \SubCellInst_LFInst_9_LFInst_0_n9 ), .B(
        \SubCellInst_LFInst_9_LFInst_0_n8 ), .Z(
        \SubCellInst_LFInst_9_LFInst_0_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_9_LFInst_1_U12  ( .A1(AddRoundKeyOutput[37]), 
        .A2(\SubCellInst_LFInst_9_LFInst_1_n16 ), .ZN(
        \SubCellInst_LFInst_9_LFInst_1_n17 ) );
  NOR2_X1 \SubCellInst_LFInst_9_LFInst_1_U11  ( .A1(AddRoundKeyOutput[39]), 
        .A2(\SubCellInst_LFInst_9_LFInst_1_n15 ), .ZN(
        \SubCellInst_LFInst_9_LFInst_1_n16 ) );
  AND2_X1 \SubCellInst_LFInst_9_LFInst_1_U10  ( .A1(AddRoundKeyOutput[36]), 
        .A2(AddRoundKeyOutput[38]), .ZN(\SubCellInst_LFInst_9_LFInst_1_n15 )
         );
  NAND2_X1 \SubCellInst_LFInst_9_LFInst_1_U9  ( .A1(AddRoundKeyOutput[39]), 
        .A2(\SubCellInst_LFInst_9_LFInst_1_n14 ), .ZN(
        \SubCellInst_LFInst_9_LFInst_1_n18 ) );
  NAND2_X1 \SubCellInst_LFInst_9_LFInst_1_U8  ( .A1(
        \SubCellInst_LFInst_9_LFInst_1_n13 ), .A2(
        \SubCellInst_LFInst_9_LFInst_1_n12 ), .ZN(
        \SubCellInst_LFInst_9_LFInst_1_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_9_LFInst_1_U7  ( .A1(AddRoundKeyOutput[36]), 
        .A2(AddRoundKeyOutput[38]), .ZN(\SubCellInst_LFInst_9_LFInst_1_n12 )
         );
  NAND2_X1 \SubCellInst_LFInst_9_LFInst_1_U6  ( .A1(
        \SubCellInst_LFInst_9_LFInst_1_n11 ), .A2(
        \SubCellInst_LFInst_9_LFInst_1_n10 ), .ZN(
        \SubCellInst_LFInst_9_LFInst_1_n13 ) );
  NAND2_X1 \SubCellInst_LFInst_9_LFInst_1_U5  ( .A1(AddRoundKeyOutput[36]), 
        .A2(AddRoundKeyOutput[37]), .ZN(\SubCellInst_LFInst_9_LFInst_1_n10 )
         );
  INV_X1 \SubCellInst_LFInst_9_LFInst_1_U4  ( .A(AddRoundKeyOutput[38]), .ZN(
        \SubCellInst_LFInst_9_LFInst_1_n11 ) );
  NAND2_X2 \SubCellInst_LFInst_9_LFInst_1_U3  ( .A1(
        \SubCellInst_LFInst_9_LFInst_1_n18 ), .A2(
        \SubCellInst_LFInst_9_LFInst_1_n17 ), .ZN(\Red_MCInst_MC1_v1_2 [1]) );
  NAND2_X1 \SubCellInst_LFInst_9_LFInst_2_U11  ( .A1(
        \SubCellInst_LFInst_9_LFInst_2_n22 ), .A2(
        \SubCellInst_LFInst_9_LFInst_2_n21 ), .ZN(\MCInst_MC1_v1_3 [3]) );
  NAND2_X1 \SubCellInst_LFInst_9_LFInst_2_U10  ( .A1(AddRoundKeyOutput[38]), 
        .A2(\SubCellInst_LFInst_9_LFInst_2_n20 ), .ZN(
        \SubCellInst_LFInst_9_LFInst_2_n21 ) );
  NOR2_X1 \SubCellInst_LFInst_9_LFInst_2_U9  ( .A1(AddRoundKeyOutput[37]), 
        .A2(\SubCellInst_LFInst_9_LFInst_2_n19 ), .ZN(
        \SubCellInst_LFInst_9_LFInst_2_n20 ) );
  INV_X1 \SubCellInst_LFInst_9_LFInst_2_U8  ( .A(AddRoundKeyOutput[39]), .ZN(
        \SubCellInst_LFInst_9_LFInst_2_n19 ) );
  NAND2_X1 \SubCellInst_LFInst_9_LFInst_2_U7  ( .A1(
        \SubCellInst_LFInst_9_LFInst_2_n18 ), .A2(
        \SubCellInst_LFInst_9_LFInst_2_n17 ), .ZN(
        \SubCellInst_LFInst_9_LFInst_2_n22 ) );
  XOR2_X1 \SubCellInst_LFInst_9_LFInst_2_U6  ( .A(
        \SubCellInst_LFInst_9_LFInst_2_n16 ), .B(AddRoundKeyOutput[38]), .Z(
        \SubCellInst_LFInst_9_LFInst_2_n17 ) );
  NAND2_X1 \SubCellInst_LFInst_9_LFInst_2_U5  ( .A1(AddRoundKeyOutput[36]), 
        .A2(AddRoundKeyOutput[37]), .ZN(\SubCellInst_LFInst_9_LFInst_2_n16 )
         );
  NAND2_X1 \SubCellInst_LFInst_9_LFInst_2_U4  ( .A1(
        \SubCellInst_LFInst_9_LFInst_2_n15 ), .A2(AddRoundKeyOutput[39]), .ZN(
        \SubCellInst_LFInst_9_LFInst_2_n18 ) );
  XNOR2_X1 \SubCellInst_LFInst_9_LFInst_2_U3  ( .A(AddRoundKeyOutput[36]), .B(
        AddRoundKeyOutput[37]), .ZN(\SubCellInst_LFInst_9_LFInst_2_n15 ) );
  NAND2_X1 \SubCellInst_LFInst_9_LFInst_3_U9  ( .A1(
        \SubCellInst_LFInst_9_LFInst_3_n16 ), .A2(
        \SubCellInst_LFInst_9_LFInst_3_n15 ), .ZN(\Red_MCInst_MC1_v1_1 [2]) );
  NAND2_X1 \SubCellInst_LFInst_9_LFInst_3_U8  ( .A1(AddRoundKeyOutput[37]), 
        .A2(\SubCellInst_LFInst_9_LFInst_3_n14 ), .ZN(
        \SubCellInst_LFInst_9_LFInst_3_n15 ) );
  XOR2_X1 \SubCellInst_LFInst_9_LFInst_3_U7  ( .A(AddRoundKeyOutput[39]), .B(
        AddRoundKeyOutput[38]), .Z(\SubCellInst_LFInst_9_LFInst_3_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_9_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_9_LFInst_3_n13 ), .A2(
        \SubCellInst_LFInst_9_LFInst_3_n12 ), .ZN(
        \SubCellInst_LFInst_9_LFInst_3_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_9_LFInst_3_U5  ( .A1(AddRoundKeyOutput[36]), 
        .A2(AddRoundKeyOutput[38]), .ZN(\SubCellInst_LFInst_9_LFInst_3_n12 )
         );
  XNOR2_X1 \SubCellInst_LFInst_9_LFInst_3_U4  ( .A(AddRoundKeyOutput[36]), .B(
        \SubCellInst_LFInst_9_LFInst_3_n11 ), .ZN(
        \SubCellInst_LFInst_9_LFInst_3_n13 ) );
  OR2_X1 \SubCellInst_LFInst_9_LFInst_3_U3  ( .A1(AddRoundKeyOutput[39]), .A2(
        AddRoundKeyOutput[37]), .ZN(\SubCellInst_LFInst_9_LFInst_3_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_10_LFInst_0_U7  ( .A1(AddRoundKeyOutput[42]), 
        .A2(\SubCellInst_LFInst_10_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_10_LFInst_0_n8 ) );
  INV_X1 \SubCellInst_LFInst_10_LFInst_0_U6  ( .A(AddRoundKeyOutput[41]), .ZN(
        \SubCellInst_LFInst_10_LFInst_0_n7 ) );
  XOR2_X1 \SubCellInst_LFInst_10_LFInst_0_U5  ( .A(AddRoundKeyOutput[40]), .B(
        AddRoundKeyOutput[43]), .Z(\SubCellInst_LFInst_10_LFInst_0_n9 ) );
  INV_X1 \SubCellInst_LFInst_10_LFInst_0_U4  ( .A(
        \SubCellInst_LFInst_10_LFInst_0_n10 ), .ZN(\MCInst_MC0_v1_0 [0]) );
  XOR2_X1 \SubCellInst_LFInst_10_LFInst_0_U3  ( .A(
        \SubCellInst_LFInst_10_LFInst_0_n9 ), .B(
        \SubCellInst_LFInst_10_LFInst_0_n8 ), .Z(
        \SubCellInst_LFInst_10_LFInst_0_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_10_LFInst_1_U12  ( .A1(AddRoundKeyOutput[41]), 
        .A2(\SubCellInst_LFInst_10_LFInst_1_n16 ), .ZN(
        \SubCellInst_LFInst_10_LFInst_1_n17 ) );
  NOR2_X1 \SubCellInst_LFInst_10_LFInst_1_U11  ( .A1(AddRoundKeyOutput[43]), 
        .A2(\SubCellInst_LFInst_10_LFInst_1_n15 ), .ZN(
        \SubCellInst_LFInst_10_LFInst_1_n16 ) );
  AND2_X1 \SubCellInst_LFInst_10_LFInst_1_U10  ( .A1(AddRoundKeyOutput[40]), 
        .A2(AddRoundKeyOutput[42]), .ZN(\SubCellInst_LFInst_10_LFInst_1_n15 )
         );
  NAND2_X1 \SubCellInst_LFInst_10_LFInst_1_U9  ( .A1(AddRoundKeyOutput[43]), 
        .A2(\SubCellInst_LFInst_10_LFInst_1_n14 ), .ZN(
        \SubCellInst_LFInst_10_LFInst_1_n18 ) );
  NAND2_X1 \SubCellInst_LFInst_10_LFInst_1_U8  ( .A1(
        \SubCellInst_LFInst_10_LFInst_1_n13 ), .A2(
        \SubCellInst_LFInst_10_LFInst_1_n12 ), .ZN(
        \SubCellInst_LFInst_10_LFInst_1_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_10_LFInst_1_U7  ( .A1(AddRoundKeyOutput[40]), 
        .A2(AddRoundKeyOutput[42]), .ZN(\SubCellInst_LFInst_10_LFInst_1_n12 )
         );
  NAND2_X1 \SubCellInst_LFInst_10_LFInst_1_U6  ( .A1(
        \SubCellInst_LFInst_10_LFInst_1_n11 ), .A2(
        \SubCellInst_LFInst_10_LFInst_1_n10 ), .ZN(
        \SubCellInst_LFInst_10_LFInst_1_n13 ) );
  NAND2_X1 \SubCellInst_LFInst_10_LFInst_1_U5  ( .A1(AddRoundKeyOutput[40]), 
        .A2(AddRoundKeyOutput[41]), .ZN(\SubCellInst_LFInst_10_LFInst_1_n10 )
         );
  INV_X1 \SubCellInst_LFInst_10_LFInst_1_U4  ( .A(AddRoundKeyOutput[42]), .ZN(
        \SubCellInst_LFInst_10_LFInst_1_n11 ) );
  NAND2_X2 \SubCellInst_LFInst_10_LFInst_1_U3  ( .A1(
        \SubCellInst_LFInst_10_LFInst_1_n18 ), .A2(
        \SubCellInst_LFInst_10_LFInst_1_n17 ), .ZN(\Red_MCInst_MC0_v1_2 [1])
         );
  NAND2_X1 \SubCellInst_LFInst_10_LFInst_2_U11  ( .A1(
        \SubCellInst_LFInst_10_LFInst_2_n22 ), .A2(
        \SubCellInst_LFInst_10_LFInst_2_n21 ), .ZN(\MCInst_MC0_v1_3 [3]) );
  NAND2_X1 \SubCellInst_LFInst_10_LFInst_2_U10  ( .A1(AddRoundKeyOutput[42]), 
        .A2(\SubCellInst_LFInst_10_LFInst_2_n20 ), .ZN(
        \SubCellInst_LFInst_10_LFInst_2_n21 ) );
  NOR2_X1 \SubCellInst_LFInst_10_LFInst_2_U9  ( .A1(AddRoundKeyOutput[41]), 
        .A2(\SubCellInst_LFInst_10_LFInst_2_n19 ), .ZN(
        \SubCellInst_LFInst_10_LFInst_2_n20 ) );
  INV_X1 \SubCellInst_LFInst_10_LFInst_2_U8  ( .A(AddRoundKeyOutput[43]), .ZN(
        \SubCellInst_LFInst_10_LFInst_2_n19 ) );
  NAND2_X1 \SubCellInst_LFInst_10_LFInst_2_U7  ( .A1(
        \SubCellInst_LFInst_10_LFInst_2_n18 ), .A2(
        \SubCellInst_LFInst_10_LFInst_2_n17 ), .ZN(
        \SubCellInst_LFInst_10_LFInst_2_n22 ) );
  XOR2_X1 \SubCellInst_LFInst_10_LFInst_2_U6  ( .A(
        \SubCellInst_LFInst_10_LFInst_2_n16 ), .B(AddRoundKeyOutput[42]), .Z(
        \SubCellInst_LFInst_10_LFInst_2_n17 ) );
  NAND2_X1 \SubCellInst_LFInst_10_LFInst_2_U5  ( .A1(AddRoundKeyOutput[40]), 
        .A2(AddRoundKeyOutput[41]), .ZN(\SubCellInst_LFInst_10_LFInst_2_n16 )
         );
  NAND2_X1 \SubCellInst_LFInst_10_LFInst_2_U4  ( .A1(
        \SubCellInst_LFInst_10_LFInst_2_n15 ), .A2(AddRoundKeyOutput[43]), 
        .ZN(\SubCellInst_LFInst_10_LFInst_2_n18 ) );
  XNOR2_X1 \SubCellInst_LFInst_10_LFInst_2_U3  ( .A(AddRoundKeyOutput[40]), 
        .B(AddRoundKeyOutput[41]), .ZN(\SubCellInst_LFInst_10_LFInst_2_n15 )
         );
  NAND2_X1 \SubCellInst_LFInst_10_LFInst_3_U9  ( .A1(
        \SubCellInst_LFInst_10_LFInst_3_n16 ), .A2(
        \SubCellInst_LFInst_10_LFInst_3_n15 ), .ZN(\Red_MCInst_MC0_v1_1 [2])
         );
  NAND2_X1 \SubCellInst_LFInst_10_LFInst_3_U8  ( .A1(AddRoundKeyOutput[41]), 
        .A2(\SubCellInst_LFInst_10_LFInst_3_n14 ), .ZN(
        \SubCellInst_LFInst_10_LFInst_3_n15 ) );
  XOR2_X1 \SubCellInst_LFInst_10_LFInst_3_U7  ( .A(AddRoundKeyOutput[43]), .B(
        AddRoundKeyOutput[42]), .Z(\SubCellInst_LFInst_10_LFInst_3_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_10_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_10_LFInst_3_n13 ), .A2(
        \SubCellInst_LFInst_10_LFInst_3_n12 ), .ZN(
        \SubCellInst_LFInst_10_LFInst_3_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_10_LFInst_3_U5  ( .A1(AddRoundKeyOutput[40]), 
        .A2(AddRoundKeyOutput[42]), .ZN(\SubCellInst_LFInst_10_LFInst_3_n12 )
         );
  XNOR2_X1 \SubCellInst_LFInst_10_LFInst_3_U4  ( .A(AddRoundKeyOutput[40]), 
        .B(\SubCellInst_LFInst_10_LFInst_3_n11 ), .ZN(
        \SubCellInst_LFInst_10_LFInst_3_n13 ) );
  OR2_X1 \SubCellInst_LFInst_10_LFInst_3_U3  ( .A1(AddRoundKeyOutput[43]), 
        .A2(AddRoundKeyOutput[41]), .ZN(\SubCellInst_LFInst_10_LFInst_3_n11 )
         );
  NAND2_X1 \SubCellInst_LFInst_11_LFInst_0_U7  ( .A1(AddRoundKeyOutput[46]), 
        .A2(\SubCellInst_LFInst_11_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_11_LFInst_0_n8 ) );
  INV_X1 \SubCellInst_LFInst_11_LFInst_0_U6  ( .A(AddRoundKeyOutput[45]), .ZN(
        \SubCellInst_LFInst_11_LFInst_0_n7 ) );
  XOR2_X1 \SubCellInst_LFInst_11_LFInst_0_U5  ( .A(AddRoundKeyOutput[44]), .B(
        AddRoundKeyOutput[47]), .Z(\SubCellInst_LFInst_11_LFInst_0_n9 ) );
  INV_X1 \SubCellInst_LFInst_11_LFInst_0_U4  ( .A(
        \SubCellInst_LFInst_11_LFInst_0_n10 ), .ZN(\MCInst_MC3_v1_0 [0]) );
  XOR2_X1 \SubCellInst_LFInst_11_LFInst_0_U3  ( .A(
        \SubCellInst_LFInst_11_LFInst_0_n9 ), .B(
        \SubCellInst_LFInst_11_LFInst_0_n8 ), .Z(
        \SubCellInst_LFInst_11_LFInst_0_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_11_LFInst_1_U12  ( .A1(AddRoundKeyOutput[45]), 
        .A2(\SubCellInst_LFInst_11_LFInst_1_n16 ), .ZN(
        \SubCellInst_LFInst_11_LFInst_1_n17 ) );
  NOR2_X1 \SubCellInst_LFInst_11_LFInst_1_U11  ( .A1(AddRoundKeyOutput[47]), 
        .A2(\SubCellInst_LFInst_11_LFInst_1_n15 ), .ZN(
        \SubCellInst_LFInst_11_LFInst_1_n16 ) );
  AND2_X1 \SubCellInst_LFInst_11_LFInst_1_U10  ( .A1(AddRoundKeyOutput[44]), 
        .A2(AddRoundKeyOutput[46]), .ZN(\SubCellInst_LFInst_11_LFInst_1_n15 )
         );
  NAND2_X1 \SubCellInst_LFInst_11_LFInst_1_U9  ( .A1(AddRoundKeyOutput[47]), 
        .A2(\SubCellInst_LFInst_11_LFInst_1_n14 ), .ZN(
        \SubCellInst_LFInst_11_LFInst_1_n18 ) );
  NAND2_X1 \SubCellInst_LFInst_11_LFInst_1_U8  ( .A1(
        \SubCellInst_LFInst_11_LFInst_1_n13 ), .A2(
        \SubCellInst_LFInst_11_LFInst_1_n12 ), .ZN(
        \SubCellInst_LFInst_11_LFInst_1_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_11_LFInst_1_U7  ( .A1(AddRoundKeyOutput[44]), 
        .A2(AddRoundKeyOutput[46]), .ZN(\SubCellInst_LFInst_11_LFInst_1_n12 )
         );
  NAND2_X1 \SubCellInst_LFInst_11_LFInst_1_U6  ( .A1(
        \SubCellInst_LFInst_11_LFInst_1_n11 ), .A2(
        \SubCellInst_LFInst_11_LFInst_1_n10 ), .ZN(
        \SubCellInst_LFInst_11_LFInst_1_n13 ) );
  NAND2_X1 \SubCellInst_LFInst_11_LFInst_1_U5  ( .A1(AddRoundKeyOutput[44]), 
        .A2(AddRoundKeyOutput[45]), .ZN(\SubCellInst_LFInst_11_LFInst_1_n10 )
         );
  INV_X1 \SubCellInst_LFInst_11_LFInst_1_U4  ( .A(AddRoundKeyOutput[46]), .ZN(
        \SubCellInst_LFInst_11_LFInst_1_n11 ) );
  NAND2_X2 \SubCellInst_LFInst_11_LFInst_1_U3  ( .A1(
        \SubCellInst_LFInst_11_LFInst_1_n18 ), .A2(
        \SubCellInst_LFInst_11_LFInst_1_n17 ), .ZN(\Red_MCInst_MC3_v1_2 [1])
         );
  NAND2_X1 \SubCellInst_LFInst_11_LFInst_2_U11  ( .A1(
        \SubCellInst_LFInst_11_LFInst_2_n22 ), .A2(
        \SubCellInst_LFInst_11_LFInst_2_n21 ), .ZN(\MCInst_MC3_v1_3 [3]) );
  NAND2_X1 \SubCellInst_LFInst_11_LFInst_2_U10  ( .A1(AddRoundKeyOutput[46]), 
        .A2(\SubCellInst_LFInst_11_LFInst_2_n20 ), .ZN(
        \SubCellInst_LFInst_11_LFInst_2_n21 ) );
  NOR2_X1 \SubCellInst_LFInst_11_LFInst_2_U9  ( .A1(AddRoundKeyOutput[45]), 
        .A2(\SubCellInst_LFInst_11_LFInst_2_n19 ), .ZN(
        \SubCellInst_LFInst_11_LFInst_2_n20 ) );
  INV_X1 \SubCellInst_LFInst_11_LFInst_2_U8  ( .A(AddRoundKeyOutput[47]), .ZN(
        \SubCellInst_LFInst_11_LFInst_2_n19 ) );
  NAND2_X1 \SubCellInst_LFInst_11_LFInst_2_U7  ( .A1(
        \SubCellInst_LFInst_11_LFInst_2_n18 ), .A2(
        \SubCellInst_LFInst_11_LFInst_2_n17 ), .ZN(
        \SubCellInst_LFInst_11_LFInst_2_n22 ) );
  XOR2_X1 \SubCellInst_LFInst_11_LFInst_2_U6  ( .A(
        \SubCellInst_LFInst_11_LFInst_2_n16 ), .B(AddRoundKeyOutput[46]), .Z(
        \SubCellInst_LFInst_11_LFInst_2_n17 ) );
  NAND2_X1 \SubCellInst_LFInst_11_LFInst_2_U5  ( .A1(AddRoundKeyOutput[44]), 
        .A2(AddRoundKeyOutput[45]), .ZN(\SubCellInst_LFInst_11_LFInst_2_n16 )
         );
  NAND2_X1 \SubCellInst_LFInst_11_LFInst_2_U4  ( .A1(
        \SubCellInst_LFInst_11_LFInst_2_n15 ), .A2(AddRoundKeyOutput[47]), 
        .ZN(\SubCellInst_LFInst_11_LFInst_2_n18 ) );
  XNOR2_X1 \SubCellInst_LFInst_11_LFInst_2_U3  ( .A(AddRoundKeyOutput[44]), 
        .B(AddRoundKeyOutput[45]), .ZN(\SubCellInst_LFInst_11_LFInst_2_n15 )
         );
  NAND2_X1 \SubCellInst_LFInst_11_LFInst_3_U9  ( .A1(
        \SubCellInst_LFInst_11_LFInst_3_n16 ), .A2(
        \SubCellInst_LFInst_11_LFInst_3_n15 ), .ZN(\Red_MCInst_MC3_v1_1 [2])
         );
  NAND2_X1 \SubCellInst_LFInst_11_LFInst_3_U8  ( .A1(AddRoundKeyOutput[45]), 
        .A2(\SubCellInst_LFInst_11_LFInst_3_n14 ), .ZN(
        \SubCellInst_LFInst_11_LFInst_3_n15 ) );
  XOR2_X1 \SubCellInst_LFInst_11_LFInst_3_U7  ( .A(AddRoundKeyOutput[47]), .B(
        AddRoundKeyOutput[46]), .Z(\SubCellInst_LFInst_11_LFInst_3_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_11_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_11_LFInst_3_n13 ), .A2(
        \SubCellInst_LFInst_11_LFInst_3_n12 ), .ZN(
        \SubCellInst_LFInst_11_LFInst_3_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_11_LFInst_3_U5  ( .A1(AddRoundKeyOutput[44]), 
        .A2(AddRoundKeyOutput[46]), .ZN(\SubCellInst_LFInst_11_LFInst_3_n12 )
         );
  XNOR2_X1 \SubCellInst_LFInst_11_LFInst_3_U4  ( .A(AddRoundKeyOutput[44]), 
        .B(\SubCellInst_LFInst_11_LFInst_3_n11 ), .ZN(
        \SubCellInst_LFInst_11_LFInst_3_n13 ) );
  OR2_X1 \SubCellInst_LFInst_11_LFInst_3_U3  ( .A1(AddRoundKeyOutput[47]), 
        .A2(AddRoundKeyOutput[45]), .ZN(\SubCellInst_LFInst_11_LFInst_3_n11 )
         );
  NAND2_X1 \SubCellInst_LFInst_12_LFInst_0_U7  ( .A1(AddRoundKeyOutput[50]), 
        .A2(\SubCellInst_LFInst_12_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_12_LFInst_0_n8 ) );
  INV_X1 \SubCellInst_LFInst_12_LFInst_0_U6  ( .A(AddRoundKeyOutput[49]), .ZN(
        \SubCellInst_LFInst_12_LFInst_0_n7 ) );
  XOR2_X1 \SubCellInst_LFInst_12_LFInst_0_U5  ( .A(AddRoundKeyOutput[48]), .B(
        AddRoundKeyOutput[51]), .Z(\SubCellInst_LFInst_12_LFInst_0_n9 ) );
  INV_X1 \SubCellInst_LFInst_12_LFInst_0_U4  ( .A(
        \SubCellInst_LFInst_12_LFInst_0_n10 ), .ZN(\Red_MCInst_MC3_v0_0 [0])
         );
  XOR2_X1 \SubCellInst_LFInst_12_LFInst_0_U3  ( .A(
        \SubCellInst_LFInst_12_LFInst_0_n9 ), .B(
        \SubCellInst_LFInst_12_LFInst_0_n8 ), .Z(
        \SubCellInst_LFInst_12_LFInst_0_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_12_LFInst_1_U12  ( .A1(
        \SubCellInst_LFInst_12_LFInst_1_n18 ), .A2(
        \SubCellInst_LFInst_12_LFInst_1_n17 ), .ZN(\Red_MCInst_MC3_v0_2 [2])
         );
  NAND2_X1 \SubCellInst_LFInst_12_LFInst_1_U11  ( .A1(AddRoundKeyOutput[49]), 
        .A2(\SubCellInst_LFInst_12_LFInst_1_n16 ), .ZN(
        \SubCellInst_LFInst_12_LFInst_1_n17 ) );
  NOR2_X1 \SubCellInst_LFInst_12_LFInst_1_U10  ( .A1(AddRoundKeyOutput[51]), 
        .A2(\SubCellInst_LFInst_12_LFInst_1_n15 ), .ZN(
        \SubCellInst_LFInst_12_LFInst_1_n16 ) );
  AND2_X1 \SubCellInst_LFInst_12_LFInst_1_U9  ( .A1(AddRoundKeyOutput[48]), 
        .A2(AddRoundKeyOutput[50]), .ZN(\SubCellInst_LFInst_12_LFInst_1_n15 )
         );
  NAND2_X1 \SubCellInst_LFInst_12_LFInst_1_U8  ( .A1(AddRoundKeyOutput[51]), 
        .A2(\SubCellInst_LFInst_12_LFInst_1_n14 ), .ZN(
        \SubCellInst_LFInst_12_LFInst_1_n18 ) );
  NAND2_X1 \SubCellInst_LFInst_12_LFInst_1_U7  ( .A1(
        \SubCellInst_LFInst_12_LFInst_1_n13 ), .A2(
        \SubCellInst_LFInst_12_LFInst_1_n12 ), .ZN(
        \SubCellInst_LFInst_12_LFInst_1_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_12_LFInst_1_U6  ( .A1(AddRoundKeyOutput[48]), 
        .A2(AddRoundKeyOutput[50]), .ZN(\SubCellInst_LFInst_12_LFInst_1_n12 )
         );
  NAND2_X1 \SubCellInst_LFInst_12_LFInst_1_U5  ( .A1(
        \SubCellInst_LFInst_12_LFInst_1_n11 ), .A2(
        \SubCellInst_LFInst_12_LFInst_1_n10 ), .ZN(
        \SubCellInst_LFInst_12_LFInst_1_n13 ) );
  NAND2_X1 \SubCellInst_LFInst_12_LFInst_1_U4  ( .A1(AddRoundKeyOutput[48]), 
        .A2(AddRoundKeyOutput[49]), .ZN(\SubCellInst_LFInst_12_LFInst_1_n10 )
         );
  INV_X1 \SubCellInst_LFInst_12_LFInst_1_U3  ( .A(AddRoundKeyOutput[50]), .ZN(
        \SubCellInst_LFInst_12_LFInst_1_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_12_LFInst_2_U11  ( .A1(
        \SubCellInst_LFInst_12_LFInst_2_n22 ), .A2(
        \SubCellInst_LFInst_12_LFInst_2_n21 ), .ZN(\MCInst_MC3_v0_3 [3]) );
  NAND2_X1 \SubCellInst_LFInst_12_LFInst_2_U10  ( .A1(AddRoundKeyOutput[50]), 
        .A2(\SubCellInst_LFInst_12_LFInst_2_n20 ), .ZN(
        \SubCellInst_LFInst_12_LFInst_2_n21 ) );
  NOR2_X1 \SubCellInst_LFInst_12_LFInst_2_U9  ( .A1(AddRoundKeyOutput[49]), 
        .A2(\SubCellInst_LFInst_12_LFInst_2_n19 ), .ZN(
        \SubCellInst_LFInst_12_LFInst_2_n20 ) );
  INV_X1 \SubCellInst_LFInst_12_LFInst_2_U8  ( .A(AddRoundKeyOutput[51]), .ZN(
        \SubCellInst_LFInst_12_LFInst_2_n19 ) );
  NAND2_X1 \SubCellInst_LFInst_12_LFInst_2_U7  ( .A1(
        \SubCellInst_LFInst_12_LFInst_2_n18 ), .A2(
        \SubCellInst_LFInst_12_LFInst_2_n17 ), .ZN(
        \SubCellInst_LFInst_12_LFInst_2_n22 ) );
  XOR2_X1 \SubCellInst_LFInst_12_LFInst_2_U6  ( .A(
        \SubCellInst_LFInst_12_LFInst_2_n16 ), .B(AddRoundKeyOutput[50]), .Z(
        \SubCellInst_LFInst_12_LFInst_2_n17 ) );
  NAND2_X1 \SubCellInst_LFInst_12_LFInst_2_U5  ( .A1(AddRoundKeyOutput[48]), 
        .A2(AddRoundKeyOutput[49]), .ZN(\SubCellInst_LFInst_12_LFInst_2_n16 )
         );
  NAND2_X1 \SubCellInst_LFInst_12_LFInst_2_U4  ( .A1(
        \SubCellInst_LFInst_12_LFInst_2_n15 ), .A2(AddRoundKeyOutput[51]), 
        .ZN(\SubCellInst_LFInst_12_LFInst_2_n18 ) );
  XNOR2_X1 \SubCellInst_LFInst_12_LFInst_2_U3  ( .A(AddRoundKeyOutput[48]), 
        .B(AddRoundKeyOutput[49]), .ZN(\SubCellInst_LFInst_12_LFInst_2_n15 )
         );
  NAND2_X1 \SubCellInst_LFInst_12_LFInst_3_U9  ( .A1(
        \SubCellInst_LFInst_12_LFInst_3_n16 ), .A2(
        \SubCellInst_LFInst_12_LFInst_3_n15 ), .ZN(\Red_MCInst_MC3_v0_1 [0])
         );
  NAND2_X1 \SubCellInst_LFInst_12_LFInst_3_U8  ( .A1(AddRoundKeyOutput[49]), 
        .A2(\SubCellInst_LFInst_12_LFInst_3_n14 ), .ZN(
        \SubCellInst_LFInst_12_LFInst_3_n15 ) );
  XOR2_X1 \SubCellInst_LFInst_12_LFInst_3_U7  ( .A(AddRoundKeyOutput[51]), .B(
        AddRoundKeyOutput[50]), .Z(\SubCellInst_LFInst_12_LFInst_3_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_12_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_12_LFInst_3_n13 ), .A2(
        \SubCellInst_LFInst_12_LFInst_3_n12 ), .ZN(
        \SubCellInst_LFInst_12_LFInst_3_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_12_LFInst_3_U5  ( .A1(AddRoundKeyOutput[48]), 
        .A2(AddRoundKeyOutput[50]), .ZN(\SubCellInst_LFInst_12_LFInst_3_n12 )
         );
  XNOR2_X1 \SubCellInst_LFInst_12_LFInst_3_U4  ( .A(AddRoundKeyOutput[48]), 
        .B(\SubCellInst_LFInst_12_LFInst_3_n11 ), .ZN(
        \SubCellInst_LFInst_12_LFInst_3_n13 ) );
  OR2_X1 \SubCellInst_LFInst_12_LFInst_3_U3  ( .A1(AddRoundKeyOutput[51]), 
        .A2(AddRoundKeyOutput[49]), .ZN(\SubCellInst_LFInst_12_LFInst_3_n11 )
         );
  NAND2_X1 \SubCellInst_LFInst_13_LFInst_0_U7  ( .A1(AddRoundKeyOutput[54]), 
        .A2(\SubCellInst_LFInst_13_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_13_LFInst_0_n8 ) );
  INV_X1 \SubCellInst_LFInst_13_LFInst_0_U6  ( .A(AddRoundKeyOutput[53]), .ZN(
        \SubCellInst_LFInst_13_LFInst_0_n7 ) );
  XOR2_X1 \SubCellInst_LFInst_13_LFInst_0_U5  ( .A(AddRoundKeyOutput[52]), .B(
        AddRoundKeyOutput[55]), .Z(\SubCellInst_LFInst_13_LFInst_0_n9 ) );
  INV_X1 \SubCellInst_LFInst_13_LFInst_0_U4  ( .A(
        \SubCellInst_LFInst_13_LFInst_0_n10 ), .ZN(\Red_MCInst_MC2_v0_0 [0])
         );
  XOR2_X1 \SubCellInst_LFInst_13_LFInst_0_U3  ( .A(
        \SubCellInst_LFInst_13_LFInst_0_n9 ), .B(
        \SubCellInst_LFInst_13_LFInst_0_n8 ), .Z(
        \SubCellInst_LFInst_13_LFInst_0_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_13_LFInst_1_U12  ( .A1(
        \SubCellInst_LFInst_13_LFInst_1_n18 ), .A2(
        \SubCellInst_LFInst_13_LFInst_1_n17 ), .ZN(\Red_MCInst_MC2_v0_2 [2])
         );
  NAND2_X1 \SubCellInst_LFInst_13_LFInst_1_U11  ( .A1(AddRoundKeyOutput[53]), 
        .A2(\SubCellInst_LFInst_13_LFInst_1_n16 ), .ZN(
        \SubCellInst_LFInst_13_LFInst_1_n17 ) );
  NOR2_X1 \SubCellInst_LFInst_13_LFInst_1_U10  ( .A1(AddRoundKeyOutput[55]), 
        .A2(\SubCellInst_LFInst_13_LFInst_1_n15 ), .ZN(
        \SubCellInst_LFInst_13_LFInst_1_n16 ) );
  AND2_X1 \SubCellInst_LFInst_13_LFInst_1_U9  ( .A1(AddRoundKeyOutput[52]), 
        .A2(AddRoundKeyOutput[54]), .ZN(\SubCellInst_LFInst_13_LFInst_1_n15 )
         );
  NAND2_X1 \SubCellInst_LFInst_13_LFInst_1_U8  ( .A1(AddRoundKeyOutput[55]), 
        .A2(\SubCellInst_LFInst_13_LFInst_1_n14 ), .ZN(
        \SubCellInst_LFInst_13_LFInst_1_n18 ) );
  NAND2_X1 \SubCellInst_LFInst_13_LFInst_1_U7  ( .A1(
        \SubCellInst_LFInst_13_LFInst_1_n13 ), .A2(
        \SubCellInst_LFInst_13_LFInst_1_n12 ), .ZN(
        \SubCellInst_LFInst_13_LFInst_1_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_13_LFInst_1_U6  ( .A1(AddRoundKeyOutput[52]), 
        .A2(AddRoundKeyOutput[54]), .ZN(\SubCellInst_LFInst_13_LFInst_1_n12 )
         );
  NAND2_X1 \SubCellInst_LFInst_13_LFInst_1_U5  ( .A1(
        \SubCellInst_LFInst_13_LFInst_1_n11 ), .A2(
        \SubCellInst_LFInst_13_LFInst_1_n10 ), .ZN(
        \SubCellInst_LFInst_13_LFInst_1_n13 ) );
  NAND2_X1 \SubCellInst_LFInst_13_LFInst_1_U4  ( .A1(AddRoundKeyOutput[52]), 
        .A2(AddRoundKeyOutput[53]), .ZN(\SubCellInst_LFInst_13_LFInst_1_n10 )
         );
  INV_X1 \SubCellInst_LFInst_13_LFInst_1_U3  ( .A(AddRoundKeyOutput[54]), .ZN(
        \SubCellInst_LFInst_13_LFInst_1_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_13_LFInst_2_U11  ( .A1(
        \SubCellInst_LFInst_13_LFInst_2_n22 ), .A2(
        \SubCellInst_LFInst_13_LFInst_2_n21 ), .ZN(\MCInst_MC2_v0_3 [3]) );
  NAND2_X1 \SubCellInst_LFInst_13_LFInst_2_U10  ( .A1(AddRoundKeyOutput[54]), 
        .A2(\SubCellInst_LFInst_13_LFInst_2_n20 ), .ZN(
        \SubCellInst_LFInst_13_LFInst_2_n21 ) );
  NOR2_X1 \SubCellInst_LFInst_13_LFInst_2_U9  ( .A1(AddRoundKeyOutput[53]), 
        .A2(\SubCellInst_LFInst_13_LFInst_2_n19 ), .ZN(
        \SubCellInst_LFInst_13_LFInst_2_n20 ) );
  INV_X1 \SubCellInst_LFInst_13_LFInst_2_U8  ( .A(AddRoundKeyOutput[55]), .ZN(
        \SubCellInst_LFInst_13_LFInst_2_n19 ) );
  NAND2_X1 \SubCellInst_LFInst_13_LFInst_2_U7  ( .A1(
        \SubCellInst_LFInst_13_LFInst_2_n18 ), .A2(
        \SubCellInst_LFInst_13_LFInst_2_n17 ), .ZN(
        \SubCellInst_LFInst_13_LFInst_2_n22 ) );
  XOR2_X1 \SubCellInst_LFInst_13_LFInst_2_U6  ( .A(
        \SubCellInst_LFInst_13_LFInst_2_n16 ), .B(AddRoundKeyOutput[54]), .Z(
        \SubCellInst_LFInst_13_LFInst_2_n17 ) );
  NAND2_X1 \SubCellInst_LFInst_13_LFInst_2_U5  ( .A1(AddRoundKeyOutput[52]), 
        .A2(AddRoundKeyOutput[53]), .ZN(\SubCellInst_LFInst_13_LFInst_2_n16 )
         );
  NAND2_X1 \SubCellInst_LFInst_13_LFInst_2_U4  ( .A1(
        \SubCellInst_LFInst_13_LFInst_2_n15 ), .A2(AddRoundKeyOutput[55]), 
        .ZN(\SubCellInst_LFInst_13_LFInst_2_n18 ) );
  XNOR2_X1 \SubCellInst_LFInst_13_LFInst_2_U3  ( .A(AddRoundKeyOutput[52]), 
        .B(AddRoundKeyOutput[53]), .ZN(\SubCellInst_LFInst_13_LFInst_2_n15 )
         );
  NAND2_X1 \SubCellInst_LFInst_13_LFInst_3_U9  ( .A1(
        \SubCellInst_LFInst_13_LFInst_3_n16 ), .A2(
        \SubCellInst_LFInst_13_LFInst_3_n15 ), .ZN(\Red_MCInst_MC2_v0_1 [0])
         );
  NAND2_X1 \SubCellInst_LFInst_13_LFInst_3_U8  ( .A1(AddRoundKeyOutput[53]), 
        .A2(\SubCellInst_LFInst_13_LFInst_3_n14 ), .ZN(
        \SubCellInst_LFInst_13_LFInst_3_n15 ) );
  XOR2_X1 \SubCellInst_LFInst_13_LFInst_3_U7  ( .A(AddRoundKeyOutput[55]), .B(
        AddRoundKeyOutput[54]), .Z(\SubCellInst_LFInst_13_LFInst_3_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_13_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_13_LFInst_3_n13 ), .A2(
        \SubCellInst_LFInst_13_LFInst_3_n12 ), .ZN(
        \SubCellInst_LFInst_13_LFInst_3_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_13_LFInst_3_U5  ( .A1(AddRoundKeyOutput[52]), 
        .A2(AddRoundKeyOutput[54]), .ZN(\SubCellInst_LFInst_13_LFInst_3_n12 )
         );
  XNOR2_X1 \SubCellInst_LFInst_13_LFInst_3_U4  ( .A(AddRoundKeyOutput[52]), 
        .B(\SubCellInst_LFInst_13_LFInst_3_n11 ), .ZN(
        \SubCellInst_LFInst_13_LFInst_3_n13 ) );
  OR2_X1 \SubCellInst_LFInst_13_LFInst_3_U3  ( .A1(AddRoundKeyOutput[55]), 
        .A2(AddRoundKeyOutput[53]), .ZN(\SubCellInst_LFInst_13_LFInst_3_n11 )
         );
  NAND2_X1 \SubCellInst_LFInst_14_LFInst_0_U7  ( .A1(AddRoundKeyOutput[58]), 
        .A2(\SubCellInst_LFInst_14_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_14_LFInst_0_n8 ) );
  INV_X1 \SubCellInst_LFInst_14_LFInst_0_U6  ( .A(AddRoundKeyOutput[57]), .ZN(
        \SubCellInst_LFInst_14_LFInst_0_n7 ) );
  XOR2_X1 \SubCellInst_LFInst_14_LFInst_0_U5  ( .A(AddRoundKeyOutput[56]), .B(
        AddRoundKeyOutput[59]), .Z(\SubCellInst_LFInst_14_LFInst_0_n9 ) );
  INV_X1 \SubCellInst_LFInst_14_LFInst_0_U4  ( .A(
        \SubCellInst_LFInst_14_LFInst_0_n10 ), .ZN(\Red_MCInst_MC1_v0_0 [0])
         );
  XOR2_X1 \SubCellInst_LFInst_14_LFInst_0_U3  ( .A(
        \SubCellInst_LFInst_14_LFInst_0_n9 ), .B(
        \SubCellInst_LFInst_14_LFInst_0_n8 ), .Z(
        \SubCellInst_LFInst_14_LFInst_0_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_14_LFInst_1_U12  ( .A1(
        \SubCellInst_LFInst_14_LFInst_1_n18 ), .A2(
        \SubCellInst_LFInst_14_LFInst_1_n17 ), .ZN(\Red_MCInst_MC1_v0_2 [2])
         );
  NAND2_X1 \SubCellInst_LFInst_14_LFInst_1_U11  ( .A1(AddRoundKeyOutput[57]), 
        .A2(\SubCellInst_LFInst_14_LFInst_1_n16 ), .ZN(
        \SubCellInst_LFInst_14_LFInst_1_n17 ) );
  NOR2_X1 \SubCellInst_LFInst_14_LFInst_1_U10  ( .A1(AddRoundKeyOutput[59]), 
        .A2(\SubCellInst_LFInst_14_LFInst_1_n15 ), .ZN(
        \SubCellInst_LFInst_14_LFInst_1_n16 ) );
  AND2_X1 \SubCellInst_LFInst_14_LFInst_1_U9  ( .A1(AddRoundKeyOutput[56]), 
        .A2(AddRoundKeyOutput[58]), .ZN(\SubCellInst_LFInst_14_LFInst_1_n15 )
         );
  NAND2_X1 \SubCellInst_LFInst_14_LFInst_1_U8  ( .A1(AddRoundKeyOutput[59]), 
        .A2(\SubCellInst_LFInst_14_LFInst_1_n14 ), .ZN(
        \SubCellInst_LFInst_14_LFInst_1_n18 ) );
  NAND2_X1 \SubCellInst_LFInst_14_LFInst_1_U7  ( .A1(
        \SubCellInst_LFInst_14_LFInst_1_n13 ), .A2(
        \SubCellInst_LFInst_14_LFInst_1_n12 ), .ZN(
        \SubCellInst_LFInst_14_LFInst_1_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_14_LFInst_1_U6  ( .A1(AddRoundKeyOutput[56]), 
        .A2(AddRoundKeyOutput[58]), .ZN(\SubCellInst_LFInst_14_LFInst_1_n12 )
         );
  NAND2_X1 \SubCellInst_LFInst_14_LFInst_1_U5  ( .A1(
        \SubCellInst_LFInst_14_LFInst_1_n11 ), .A2(
        \SubCellInst_LFInst_14_LFInst_1_n10 ), .ZN(
        \SubCellInst_LFInst_14_LFInst_1_n13 ) );
  NAND2_X1 \SubCellInst_LFInst_14_LFInst_1_U4  ( .A1(AddRoundKeyOutput[56]), 
        .A2(AddRoundKeyOutput[57]), .ZN(\SubCellInst_LFInst_14_LFInst_1_n10 )
         );
  INV_X1 \SubCellInst_LFInst_14_LFInst_1_U3  ( .A(AddRoundKeyOutput[58]), .ZN(
        \SubCellInst_LFInst_14_LFInst_1_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_14_LFInst_2_U11  ( .A1(
        \SubCellInst_LFInst_14_LFInst_2_n22 ), .A2(
        \SubCellInst_LFInst_14_LFInst_2_n21 ), .ZN(\MCInst_MC1_v0_3 [3]) );
  NAND2_X1 \SubCellInst_LFInst_14_LFInst_2_U10  ( .A1(AddRoundKeyOutput[58]), 
        .A2(\SubCellInst_LFInst_14_LFInst_2_n20 ), .ZN(
        \SubCellInst_LFInst_14_LFInst_2_n21 ) );
  NOR2_X1 \SubCellInst_LFInst_14_LFInst_2_U9  ( .A1(AddRoundKeyOutput[57]), 
        .A2(\SubCellInst_LFInst_14_LFInst_2_n19 ), .ZN(
        \SubCellInst_LFInst_14_LFInst_2_n20 ) );
  INV_X1 \SubCellInst_LFInst_14_LFInst_2_U8  ( .A(AddRoundKeyOutput[59]), .ZN(
        \SubCellInst_LFInst_14_LFInst_2_n19 ) );
  NAND2_X1 \SubCellInst_LFInst_14_LFInst_2_U7  ( .A1(
        \SubCellInst_LFInst_14_LFInst_2_n18 ), .A2(
        \SubCellInst_LFInst_14_LFInst_2_n17 ), .ZN(
        \SubCellInst_LFInst_14_LFInst_2_n22 ) );
  XOR2_X1 \SubCellInst_LFInst_14_LFInst_2_U6  ( .A(
        \SubCellInst_LFInst_14_LFInst_2_n16 ), .B(AddRoundKeyOutput[58]), .Z(
        \SubCellInst_LFInst_14_LFInst_2_n17 ) );
  NAND2_X1 \SubCellInst_LFInst_14_LFInst_2_U5  ( .A1(AddRoundKeyOutput[56]), 
        .A2(AddRoundKeyOutput[57]), .ZN(\SubCellInst_LFInst_14_LFInst_2_n16 )
         );
  NAND2_X1 \SubCellInst_LFInst_14_LFInst_2_U4  ( .A1(
        \SubCellInst_LFInst_14_LFInst_2_n15 ), .A2(AddRoundKeyOutput[59]), 
        .ZN(\SubCellInst_LFInst_14_LFInst_2_n18 ) );
  XNOR2_X1 \SubCellInst_LFInst_14_LFInst_2_U3  ( .A(AddRoundKeyOutput[56]), 
        .B(AddRoundKeyOutput[57]), .ZN(\SubCellInst_LFInst_14_LFInst_2_n15 )
         );
  NAND2_X1 \SubCellInst_LFInst_14_LFInst_3_U9  ( .A1(
        \SubCellInst_LFInst_14_LFInst_3_n16 ), .A2(
        \SubCellInst_LFInst_14_LFInst_3_n15 ), .ZN(\Red_MCInst_MC1_v0_1 [0])
         );
  NAND2_X1 \SubCellInst_LFInst_14_LFInst_3_U8  ( .A1(AddRoundKeyOutput[57]), 
        .A2(\SubCellInst_LFInst_14_LFInst_3_n14 ), .ZN(
        \SubCellInst_LFInst_14_LFInst_3_n15 ) );
  XOR2_X1 \SubCellInst_LFInst_14_LFInst_3_U7  ( .A(AddRoundKeyOutput[59]), .B(
        AddRoundKeyOutput[58]), .Z(\SubCellInst_LFInst_14_LFInst_3_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_14_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_14_LFInst_3_n13 ), .A2(
        \SubCellInst_LFInst_14_LFInst_3_n12 ), .ZN(
        \SubCellInst_LFInst_14_LFInst_3_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_14_LFInst_3_U5  ( .A1(AddRoundKeyOutput[56]), 
        .A2(AddRoundKeyOutput[58]), .ZN(\SubCellInst_LFInst_14_LFInst_3_n12 )
         );
  XNOR2_X1 \SubCellInst_LFInst_14_LFInst_3_U4  ( .A(AddRoundKeyOutput[56]), 
        .B(\SubCellInst_LFInst_14_LFInst_3_n11 ), .ZN(
        \SubCellInst_LFInst_14_LFInst_3_n13 ) );
  OR2_X1 \SubCellInst_LFInst_14_LFInst_3_U3  ( .A1(AddRoundKeyOutput[59]), 
        .A2(AddRoundKeyOutput[57]), .ZN(\SubCellInst_LFInst_14_LFInst_3_n11 )
         );
  NAND2_X1 \SubCellInst_LFInst_15_LFInst_0_U7  ( .A1(AddRoundKeyOutput[62]), 
        .A2(\SubCellInst_LFInst_15_LFInst_0_n7 ), .ZN(
        \SubCellInst_LFInst_15_LFInst_0_n8 ) );
  INV_X1 \SubCellInst_LFInst_15_LFInst_0_U6  ( .A(AddRoundKeyOutput[61]), .ZN(
        \SubCellInst_LFInst_15_LFInst_0_n7 ) );
  XOR2_X1 \SubCellInst_LFInst_15_LFInst_0_U5  ( .A(AddRoundKeyOutput[60]), .B(
        AddRoundKeyOutput[63]), .Z(\SubCellInst_LFInst_15_LFInst_0_n9 ) );
  INV_X1 \SubCellInst_LFInst_15_LFInst_0_U4  ( .A(
        \SubCellInst_LFInst_15_LFInst_0_n10 ), .ZN(\Red_MCInst_MC0_v0_0 [0])
         );
  XOR2_X1 \SubCellInst_LFInst_15_LFInst_0_U3  ( .A(
        \SubCellInst_LFInst_15_LFInst_0_n9 ), .B(
        \SubCellInst_LFInst_15_LFInst_0_n8 ), .Z(
        \SubCellInst_LFInst_15_LFInst_0_n10 ) );
  NAND2_X1 \SubCellInst_LFInst_15_LFInst_1_U12  ( .A1(
        \SubCellInst_LFInst_15_LFInst_1_n18 ), .A2(
        \SubCellInst_LFInst_15_LFInst_1_n17 ), .ZN(\Red_MCInst_MC0_v0_2 [2])
         );
  NAND2_X1 \SubCellInst_LFInst_15_LFInst_1_U11  ( .A1(AddRoundKeyOutput[61]), 
        .A2(\SubCellInst_LFInst_15_LFInst_1_n16 ), .ZN(
        \SubCellInst_LFInst_15_LFInst_1_n17 ) );
  NOR2_X1 \SubCellInst_LFInst_15_LFInst_1_U10  ( .A1(AddRoundKeyOutput[63]), 
        .A2(\SubCellInst_LFInst_15_LFInst_1_n15 ), .ZN(
        \SubCellInst_LFInst_15_LFInst_1_n16 ) );
  AND2_X1 \SubCellInst_LFInst_15_LFInst_1_U9  ( .A1(AddRoundKeyOutput[60]), 
        .A2(AddRoundKeyOutput[62]), .ZN(\SubCellInst_LFInst_15_LFInst_1_n15 )
         );
  NAND2_X1 \SubCellInst_LFInst_15_LFInst_1_U8  ( .A1(AddRoundKeyOutput[63]), 
        .A2(\SubCellInst_LFInst_15_LFInst_1_n14 ), .ZN(
        \SubCellInst_LFInst_15_LFInst_1_n18 ) );
  NAND2_X1 \SubCellInst_LFInst_15_LFInst_1_U7  ( .A1(
        \SubCellInst_LFInst_15_LFInst_1_n13 ), .A2(
        \SubCellInst_LFInst_15_LFInst_1_n12 ), .ZN(
        \SubCellInst_LFInst_15_LFInst_1_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_15_LFInst_1_U6  ( .A1(AddRoundKeyOutput[60]), 
        .A2(AddRoundKeyOutput[62]), .ZN(\SubCellInst_LFInst_15_LFInst_1_n12 )
         );
  NAND2_X1 \SubCellInst_LFInst_15_LFInst_1_U5  ( .A1(
        \SubCellInst_LFInst_15_LFInst_1_n11 ), .A2(
        \SubCellInst_LFInst_15_LFInst_1_n10 ), .ZN(
        \SubCellInst_LFInst_15_LFInst_1_n13 ) );
  NAND2_X1 \SubCellInst_LFInst_15_LFInst_1_U4  ( .A1(AddRoundKeyOutput[60]), 
        .A2(AddRoundKeyOutput[61]), .ZN(\SubCellInst_LFInst_15_LFInst_1_n10 )
         );
  INV_X1 \SubCellInst_LFInst_15_LFInst_1_U3  ( .A(AddRoundKeyOutput[62]), .ZN(
        \SubCellInst_LFInst_15_LFInst_1_n11 ) );
  NAND2_X1 \SubCellInst_LFInst_15_LFInst_2_U11  ( .A1(
        \SubCellInst_LFInst_15_LFInst_2_n22 ), .A2(
        \SubCellInst_LFInst_15_LFInst_2_n21 ), .ZN(\MCInst_MC0_v0_3 [3]) );
  NAND2_X1 \SubCellInst_LFInst_15_LFInst_2_U10  ( .A1(AddRoundKeyOutput[62]), 
        .A2(\SubCellInst_LFInst_15_LFInst_2_n20 ), .ZN(
        \SubCellInst_LFInst_15_LFInst_2_n21 ) );
  NOR2_X1 \SubCellInst_LFInst_15_LFInst_2_U9  ( .A1(AddRoundKeyOutput[61]), 
        .A2(\SubCellInst_LFInst_15_LFInst_2_n19 ), .ZN(
        \SubCellInst_LFInst_15_LFInst_2_n20 ) );
  INV_X1 \SubCellInst_LFInst_15_LFInst_2_U8  ( .A(AddRoundKeyOutput[63]), .ZN(
        \SubCellInst_LFInst_15_LFInst_2_n19 ) );
  NAND2_X1 \SubCellInst_LFInst_15_LFInst_2_U7  ( .A1(
        \SubCellInst_LFInst_15_LFInst_2_n18 ), .A2(
        \SubCellInst_LFInst_15_LFInst_2_n17 ), .ZN(
        \SubCellInst_LFInst_15_LFInst_2_n22 ) );
  XOR2_X1 \SubCellInst_LFInst_15_LFInst_2_U6  ( .A(
        \SubCellInst_LFInst_15_LFInst_2_n16 ), .B(AddRoundKeyOutput[62]), .Z(
        \SubCellInst_LFInst_15_LFInst_2_n17 ) );
  NAND2_X1 \SubCellInst_LFInst_15_LFInst_2_U5  ( .A1(AddRoundKeyOutput[60]), 
        .A2(AddRoundKeyOutput[61]), .ZN(\SubCellInst_LFInst_15_LFInst_2_n16 )
         );
  NAND2_X1 \SubCellInst_LFInst_15_LFInst_2_U4  ( .A1(
        \SubCellInst_LFInst_15_LFInst_2_n15 ), .A2(AddRoundKeyOutput[63]), 
        .ZN(\SubCellInst_LFInst_15_LFInst_2_n18 ) );
  XNOR2_X1 \SubCellInst_LFInst_15_LFInst_2_U3  ( .A(AddRoundKeyOutput[60]), 
        .B(AddRoundKeyOutput[61]), .ZN(\SubCellInst_LFInst_15_LFInst_2_n15 )
         );
  NAND2_X1 \SubCellInst_LFInst_15_LFInst_3_U9  ( .A1(
        \SubCellInst_LFInst_15_LFInst_3_n16 ), .A2(
        \SubCellInst_LFInst_15_LFInst_3_n15 ), .ZN(\Red_MCInst_MC0_v0_1 [0])
         );
  NAND2_X1 \SubCellInst_LFInst_15_LFInst_3_U8  ( .A1(AddRoundKeyOutput[61]), 
        .A2(\SubCellInst_LFInst_15_LFInst_3_n14 ), .ZN(
        \SubCellInst_LFInst_15_LFInst_3_n15 ) );
  XOR2_X1 \SubCellInst_LFInst_15_LFInst_3_U7  ( .A(AddRoundKeyOutput[63]), .B(
        AddRoundKeyOutput[62]), .Z(\SubCellInst_LFInst_15_LFInst_3_n14 ) );
  NAND2_X1 \SubCellInst_LFInst_15_LFInst_3_U6  ( .A1(
        \SubCellInst_LFInst_15_LFInst_3_n13 ), .A2(
        \SubCellInst_LFInst_15_LFInst_3_n12 ), .ZN(
        \SubCellInst_LFInst_15_LFInst_3_n16 ) );
  NAND2_X1 \SubCellInst_LFInst_15_LFInst_3_U5  ( .A1(AddRoundKeyOutput[60]), 
        .A2(AddRoundKeyOutput[62]), .ZN(\SubCellInst_LFInst_15_LFInst_3_n12 )
         );
  XNOR2_X1 \SubCellInst_LFInst_15_LFInst_3_U4  ( .A(AddRoundKeyOutput[60]), 
        .B(\SubCellInst_LFInst_15_LFInst_3_n11 ), .ZN(
        \SubCellInst_LFInst_15_LFInst_3_n13 ) );
  OR2_X1 \SubCellInst_LFInst_15_LFInst_3_U3  ( .A1(AddRoundKeyOutput[63]), 
        .A2(AddRoundKeyOutput[61]), .ZN(\SubCellInst_LFInst_15_LFInst_3_n11 )
         );
  XNOR2_X1 \MCInst_MC0_v0_2Inst_0_U4  ( .A(\MCInst_MC0_v0_2Inst_0_n2 ), .B(
        \Red_MCInst_MC0_v0_2 [2]), .ZN(\MCInst_MC0_v0_2 [0]) );
  XNOR2_X1 \MCInst_MC0_v0_2Inst_0_U3  ( .A(\Red_MCInst_MC0_v0_1 [0]), .B(
        \Red_MCInst_MC0_v0_0 [0]), .ZN(\MCInst_MC0_v0_2Inst_0_n2 ) );
  XOR2_X1 \MCInst_MC0_v1_1Inst_0_U3  ( .A(\MCInst_MC0_v1_3 [3]), .B(
        \Red_MCInst_MC0_v1_1 [2]), .Z(\MCInst_MC0_v1_1 [0]) );
  XNOR2_X1 \MCInst_MC0_v1_2Inst_0_U4  ( .A(\MCInst_MC0_v1_2Inst_0_n2 ), .B(
        \MCInst_MC0_v1_3 [3]), .ZN(\MCInst_MC0_v1_2 [0]) );
  XNOR2_X1 \MCInst_MC0_v1_2Inst_0_U3  ( .A(\Red_MCInst_MC0_v1_1 [2]), .B(
        \Red_MCInst_MC0_v1_2 [1]), .ZN(\MCInst_MC0_v1_2Inst_0_n2 ) );
  XOR2_X1 \MCInst_MC0_v2_1Inst_0_U3  ( .A(\Red_MCInst_MC0_v2_1 [1]), .B(
        \MCInst_MC0_v2_0 [3]), .Z(\MCInst_MC0_v2_1 [0]) );
  XOR2_X1 \MCInst_MC0_v2_2Inst_0_U3  ( .A(\MCInst_MC0_v2_0 [2]), .B(
        \Red_MCInst_MC0_v2_2 [1]), .Z(\MCInst_MC0_v2_2 [0]) );
  XNOR2_X1 \MCInst_MC0_v2_3Inst_0_U5  ( .A(\MCInst_MC0_v2_3Inst_0_n4 ), .B(
        \MCInst_MC0_v2_3Inst_0_n3 ), .ZN(\MCInst_MC0_v2_3 [0]) );
  XNOR2_X1 \MCInst_MC0_v2_3Inst_0_U4  ( .A(\MCInst_MC0_v2_0 [2]), .B(
        \Red_MCInst_MC0_v2_1 [1]), .ZN(\MCInst_MC0_v2_3Inst_0_n3 ) );
  XOR2_X1 \MCInst_MC0_v2_3Inst_0_U3  ( .A(\MCInst_MC0_v2_0 [3]), .B(
        \Red_MCInst_MC0_v2_2 [1]), .Z(\MCInst_MC0_v2_3Inst_0_n4 ) );
  XOR2_X1 \MCInst_MC0_v3_1Inst_0_U3  ( .A(\MCInst_MC0_v3_0 [3]), .B(
        \Red_MCInst_MC0_v3_1 [2]), .Z(\MCInst_MC0_v3_1 [0]) );
  XOR2_X1 \MCInst_MC0_v3_2Inst_0_U3  ( .A(\MCInst_MC0_v3_2 [3]), .B(
        \Red_MCInst_MC0_v3_3 [2]), .Z(\MCInst_MC0_v3_2 [0]) );
  XNOR2_X1 \MCInst_MC0_v3_3Inst_0_U4  ( .A(\MCInst_MC0_v3_3Inst_0_n2 ), .B(
        \Red_MCInst_MC0_v3_3 [2]), .ZN(\MCInst_MC0_v3_3 [0]) );
  XNOR2_X1 \MCInst_MC0_v3_3Inst_0_U3  ( .A(\Red_MCInst_MC0_v3_1 [2]), .B(
        \MCInst_MC0_v3_2 [3]), .ZN(\MCInst_MC0_v3_3Inst_0_n2 ) );
  XOR2_X1 \MCInst_MC0_v0_0Inst_1_U3  ( .A(\MCInst_MC0_v0_3 [3]), .B(
        \Red_MCInst_MC0_v0_1 [0]), .Z(\MCInst_MC0_v0_0 [1]) );
  XOR2_X1 \MCInst_MC0_v0_1Inst_1_U3  ( .A(\Red_MCInst_MC0_v0_2 [2]), .B(
        \MCInst_MC0_v0_3 [3]), .Z(\MCInst_MC0_v0_1 [1]) );
  XNOR2_X1 \MCInst_MC0_v0_2Inst_1_U4  ( .A(\MCInst_MC0_v0_2Inst_1_n2 ), .B(
        \MCInst_MC0_v0_3 [3]), .ZN(\MCInst_MC0_v0_2 [1]) );
  XNOR2_X1 \MCInst_MC0_v0_2Inst_1_U3  ( .A(\Red_MCInst_MC0_v0_1 [0]), .B(
        \Red_MCInst_MC0_v0_0 [0]), .ZN(\MCInst_MC0_v0_2Inst_1_n2 ) );
  XOR2_X1 \MCInst_MC0_v0_3Inst_1_U3  ( .A(\Red_MCInst_MC0_v0_0 [0]), .B(
        \Red_MCInst_MC0_v0_1 [0]), .Z(\MCInst_MC0_v0_3 [1]) );
  XOR2_X1 \MCInst_MC0_v1_1Inst_1_U3  ( .A(\MCInst_MC0_v1_0 [0]), .B(
        \MCInst_MC0_v1_3 [3]), .Z(\MCInst_MC0_v1_1 [1]) );
  XOR2_X1 \MCInst_MC0_v1_2Inst_1_U3  ( .A(\MCInst_MC0_v1_0 [0]), .B(
        \Red_MCInst_MC0_v1_2 [1]), .Z(\MCInst_MC0_v1_2 [1]) );
  XOR2_X1 \MCInst_MC0_v1_3Inst_1_U3  ( .A(\MCInst_MC0_v1_0 [0]), .B(
        \Red_MCInst_MC0_v1_1 [2]), .Z(\MCInst_MC0_v1_3 [1]) );
  XOR2_X1 \MCInst_MC0_v2_0Inst_1_U3  ( .A(\Red_MCInst_MC0_v2_1 [1]), .B(
        \Red_MCInst_MC0_v2_2 [1]), .Z(\MCInst_MC0_v2_0 [1]) );
  XNOR2_X1 \MCInst_MC0_v2_1Inst_1_U4  ( .A(\MCInst_MC0_v2_1Inst_1_n2 ), .B(
        \MCInst_MC0_v2_0 [3]), .ZN(\MCInst_MC0_v2_1 [1]) );
  XNOR2_X1 \MCInst_MC0_v2_1Inst_1_U3  ( .A(\Red_MCInst_MC0_v2_2 [1]), .B(
        \MCInst_MC0_v2_0 [2]), .ZN(\MCInst_MC0_v2_1Inst_1_n2 ) );
  XNOR2_X1 \MCInst_MC0_v2_2Inst_1_U5  ( .A(\MCInst_MC0_v2_2Inst_1_n4 ), .B(
        \MCInst_MC0_v2_2Inst_1_n3 ), .ZN(\MCInst_MC0_v2_2 [1]) );
  XNOR2_X1 \MCInst_MC0_v2_2Inst_1_U4  ( .A(\MCInst_MC0_v2_0 [2]), .B(
        \Red_MCInst_MC0_v2_1 [1]), .ZN(\MCInst_MC0_v2_2Inst_1_n3 ) );
  XOR2_X1 \MCInst_MC0_v2_2Inst_1_U3  ( .A(\MCInst_MC0_v2_0 [3]), .B(
        \Red_MCInst_MC0_v2_2 [1]), .Z(\MCInst_MC0_v2_2Inst_1_n4 ) );
  XOR2_X1 \MCInst_MC0_v3_0Inst_1_U3  ( .A(\MCInst_MC0_v3_2 [3]), .B(
        \Red_MCInst_MC0_v3_1 [2]), .Z(\MCInst_MC0_v3_0 [1]) );
  XOR2_X1 \MCInst_MC0_v3_1Inst_1_U3  ( .A(\MCInst_MC0_v3_2 [3]), .B(
        \MCInst_MC0_v3_0 [3]), .Z(\MCInst_MC0_v3_1 [1]) );
  XNOR2_X1 \MCInst_MC0_v3_3Inst_1_U4  ( .A(\MCInst_MC0_v3_3Inst_1_n2 ), .B(
        \MCInst_MC0_v3_0 [3]), .ZN(\MCInst_MC0_v3_3 [1]) );
  XNOR2_X1 \MCInst_MC0_v3_3Inst_1_U3  ( .A(\Red_MCInst_MC0_v3_1 [2]), .B(
        \MCInst_MC0_v3_2 [3]), .ZN(\MCInst_MC0_v3_3Inst_1_n2 ) );
  XOR2_X1 \MCInst_MC0_v0_0Inst_2_U3  ( .A(\Red_MCInst_MC0_v0_0 [0]), .B(
        \Red_MCInst_MC0_v0_1 [0]), .Z(\MCInst_MC0_v0_0 [2]) );
  XOR2_X1 \MCInst_MC0_v0_1Inst_2_U3  ( .A(\MCInst_MC0_v0_3 [3]), .B(
        \Red_MCInst_MC0_v0_1 [0]), .Z(\MCInst_MC0_v0_1 [2]) );
  XOR2_X1 \MCInst_MC0_v0_2Inst_2_U3  ( .A(\Red_MCInst_MC0_v0_2 [2]), .B(
        \Red_MCInst_MC0_v0_1 [0]), .Z(\MCInst_MC0_v0_2 [2]) );
  XNOR2_X1 \MCInst_MC0_v1_1Inst_2_U4  ( .A(\MCInst_MC0_v1_1Inst_2_n2 ), .B(
        \Red_MCInst_MC0_v1_2 [1]), .ZN(\MCInst_MC0_v1_1 [2]) );
  XNOR2_X1 \MCInst_MC0_v1_1Inst_2_U3  ( .A(\Red_MCInst_MC0_v1_1 [2]), .B(
        \MCInst_MC0_v1_0 [0]), .ZN(\MCInst_MC0_v1_1Inst_2_n2 ) );
  XNOR2_X1 \MCInst_MC0_v1_2Inst_2_U4  ( .A(\MCInst_MC0_v1_2Inst_2_n2 ), .B(
        \Red_MCInst_MC0_v1_2 [1]), .ZN(\MCInst_MC0_v1_2 [2]) );
  XNOR2_X1 \MCInst_MC0_v1_2Inst_2_U3  ( .A(\MCInst_MC0_v1_3 [3]), .B(
        \MCInst_MC0_v1_0 [0]), .ZN(\MCInst_MC0_v1_2Inst_2_n2 ) );
  XNOR2_X1 \MCInst_MC0_v2_1Inst_2_U4  ( .A(\MCInst_MC0_v2_1Inst_2_n2 ), .B(
        \MCInst_MC0_v2_0 [3]), .ZN(\MCInst_MC0_v2_1 [2]) );
  XNOR2_X1 \MCInst_MC0_v2_1Inst_2_U3  ( .A(\Red_MCInst_MC0_v2_2 [1]), .B(
        \Red_MCInst_MC0_v2_1 [1]), .ZN(\MCInst_MC0_v2_1Inst_2_n2 ) );
  XNOR2_X1 \MCInst_MC0_v2_2Inst_2_U4  ( .A(\MCInst_MC0_v2_2Inst_2_n2 ), .B(
        \MCInst_MC0_v2_0 [3]), .ZN(\MCInst_MC0_v2_2 [2]) );
  XNOR2_X1 \MCInst_MC0_v2_2Inst_2_U3  ( .A(\Red_MCInst_MC0_v2_2 [1]), .B(
        \MCInst_MC0_v2_0 [2]), .ZN(\MCInst_MC0_v2_2Inst_2_n2 ) );
  XOR2_X1 \MCInst_MC0_v2_3Inst_2_U3  ( .A(\Red_MCInst_MC0_v2_1 [1]), .B(
        \MCInst_MC0_v2_0 [2]), .Z(\MCInst_MC0_v2_3 [2]) );
  XNOR2_X1 \MCInst_MC0_v3_1Inst_2_U4  ( .A(\MCInst_MC0_v3_1Inst_2_n2 ), .B(
        \Red_MCInst_MC0_v3_3 [2]), .ZN(\MCInst_MC0_v3_1 [2]) );
  XNOR2_X1 \MCInst_MC0_v3_1Inst_2_U3  ( .A(\Red_MCInst_MC0_v3_1 [2]), .B(
        \MCInst_MC0_v3_2 [3]), .ZN(\MCInst_MC0_v3_1Inst_2_n2 ) );
  XOR2_X1 \MCInst_MC0_v3_3Inst_2_U3  ( .A(\Red_MCInst_MC0_v3_3 [2]), .B(
        \Red_MCInst_MC0_v3_1 [2]), .Z(\MCInst_MC0_v3_3 [2]) );
  XOR2_X1 \MCInst_MC0_v0_1Inst_3_U3  ( .A(\Red_MCInst_MC0_v0_0 [0]), .B(
        \Red_MCInst_MC0_v0_1 [0]), .Z(\MCInst_MC0_v0_1 [3]) );
  XOR2_X1 \MCInst_MC0_v0_2Inst_3_U3  ( .A(\Red_MCInst_MC0_v0_0 [0]), .B(
        \MCInst_MC0_v0_3 [3]), .Z(\MCInst_MC0_v0_2 [3]) );
  XOR2_X1 \MCInst_MC0_v1_1Inst_3_U3  ( .A(\Red_MCInst_MC0_v1_2 [1]), .B(
        \MCInst_MC0_v1_3 [3]), .Z(\MCInst_MC0_v1_1 [3]) );
  XNOR2_X1 \MCInst_MC0_v1_2Inst_3_U5  ( .A(\MCInst_MC0_v1_2Inst_3_n4 ), .B(
        \MCInst_MC0_v1_2Inst_3_n3 ), .ZN(\MCInst_MC0_v1_2 [3]) );
  XNOR2_X1 \MCInst_MC0_v1_2Inst_3_U4  ( .A(\Red_MCInst_MC0_v1_2 [1]), .B(
        \MCInst_MC0_v1_0 [0]), .ZN(\MCInst_MC0_v1_2Inst_3_n3 ) );
  XOR2_X1 \MCInst_MC0_v1_2Inst_3_U3  ( .A(\MCInst_MC0_v1_3 [3]), .B(
        \Red_MCInst_MC0_v1_1 [2]), .Z(\MCInst_MC0_v1_2Inst_3_n4 ) );
  XOR2_X1 \MCInst_MC0_v2_1Inst_3_U3  ( .A(\MCInst_MC0_v2_0 [2]), .B(
        \Red_MCInst_MC0_v2_2 [1]), .Z(\MCInst_MC0_v2_1 [3]) );
  XNOR2_X1 \MCInst_MC0_v2_2Inst_3_U4  ( .A(\MCInst_MC0_v2_2Inst_3_n2 ), .B(
        \MCInst_MC0_v2_0 [3]), .ZN(\MCInst_MC0_v2_2 [3]) );
  XNOR2_X1 \MCInst_MC0_v2_2Inst_3_U3  ( .A(\Red_MCInst_MC0_v2_2 [1]), .B(
        \Red_MCInst_MC0_v2_1 [1]), .ZN(\MCInst_MC0_v2_2Inst_3_n2 ) );
  XNOR2_X1 \MCInst_MC0_v2_3Inst_3_U4  ( .A(\MCInst_MC0_v2_3Inst_3_n2 ), .B(
        \MCInst_MC0_v2_0 [2]), .ZN(\MCInst_MC0_v2_3 [3]) );
  XNOR2_X1 \MCInst_MC0_v2_3Inst_3_U3  ( .A(\MCInst_MC0_v2_0 [3]), .B(
        \Red_MCInst_MC0_v2_1 [1]), .ZN(\MCInst_MC0_v2_3Inst_3_n2 ) );
  XOR2_X1 \MCInst_MC0_v3_1Inst_3_U3  ( .A(\Red_MCInst_MC0_v3_3 [2]), .B(
        \MCInst_MC0_v3_0 [3]), .Z(\MCInst_MC0_v3_1 [3]) );
  XOR2_X1 \MCInst_MC0_v3_3Inst_3_U3  ( .A(\MCInst_MC0_v3_2 [3]), .B(
        \MCInst_MC0_v3_0 [3]), .Z(\MCInst_MC0_v3_3 [3]) );
  XNOR2_X1 \MCInst_MC0_r0Inst_XORInst_0_0_U3  ( .A(
        \MCInst_MC0_r0Inst_XORInst_0_0_n5 ), .B(
        \MCInst_MC0_r0Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[60]) );
  XNOR2_X1 \MCInst_MC0_r0Inst_XORInst_0_0_U2  ( .A(\Red_MCInst_MC0_v3_1 [2]), 
        .B(\Red_MCInst_MC0_v2_2 [1]), .ZN(\MCInst_MC0_r0Inst_XORInst_0_0_n4 )
         );
  XOR2_X1 \MCInst_MC0_r0Inst_XORInst_0_0_U1  ( .A(\MCInst_MC0_v0_3 [3]), .B(
        \MCInst_MC0_v1_0 [0]), .Z(\MCInst_MC0_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \MCInst_MC0_r0Inst_XORInst_0_1_U3  ( .A(
        \MCInst_MC0_r0Inst_XORInst_0_1_n5 ), .B(
        \MCInst_MC0_r0Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[61]) );
  XNOR2_X1 \MCInst_MC0_r0Inst_XORInst_0_1_U2  ( .A(\MCInst_MC0_v3_0 [1]), .B(
        \MCInst_MC0_v2_0 [1]), .ZN(\MCInst_MC0_r0Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \MCInst_MC0_r0Inst_XORInst_0_1_U1  ( .A(\MCInst_MC0_v0_0 [1]), .B(
        \Red_MCInst_MC0_v1_2 [1]), .Z(\MCInst_MC0_r0Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \MCInst_MC0_r0Inst_XORInst_0_2_U3  ( .A(
        \MCInst_MC0_r0Inst_XORInst_0_2_n5 ), .B(
        \MCInst_MC0_r0Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[62]) );
  XNOR2_X1 \MCInst_MC0_r0Inst_XORInst_0_2_U2  ( .A(\Red_MCInst_MC0_v3_3 [2]), 
        .B(\MCInst_MC0_v2_0 [2]), .ZN(\MCInst_MC0_r0Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \MCInst_MC0_r0Inst_XORInst_0_2_U1  ( .A(\MCInst_MC0_v0_0 [2]), .B(
        \MCInst_MC0_v1_3 [3]), .Z(\MCInst_MC0_r0Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \MCInst_MC0_r0Inst_XORInst_0_3_U3  ( .A(
        \MCInst_MC0_r0Inst_XORInst_0_3_n5 ), .B(
        \MCInst_MC0_r0Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[63]) );
  XNOR2_X1 \MCInst_MC0_r0Inst_XORInst_0_3_U2  ( .A(\MCInst_MC0_v3_0 [3]), .B(
        \MCInst_MC0_v2_0 [3]), .ZN(\MCInst_MC0_r0Inst_XORInst_0_3_n4 ) );
  XOR2_X1 \MCInst_MC0_r0Inst_XORInst_0_3_U1  ( .A(\Red_MCInst_MC0_v0_2 [2]), 
        .B(\Red_MCInst_MC0_v1_1 [2]), .Z(\MCInst_MC0_r0Inst_XORInst_0_3_n5 )
         );
  XNOR2_X1 \MCInst_MC0_r1Inst_XORInst_0_0_U3  ( .A(
        \MCInst_MC0_r1Inst_XORInst_0_0_n5 ), .B(
        \MCInst_MC0_r1Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[44]) );
  XNOR2_X1 \MCInst_MC0_r1Inst_XORInst_0_0_U2  ( .A(\MCInst_MC0_v3_1 [0]), .B(
        \MCInst_MC0_v2_1 [0]), .ZN(\MCInst_MC0_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \MCInst_MC0_r1Inst_XORInst_0_0_U1  ( .A(\Red_MCInst_MC0_v0_2 [2]), 
        .B(\MCInst_MC0_v1_1 [0]), .Z(\MCInst_MC0_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \MCInst_MC0_r1Inst_XORInst_0_1_U3  ( .A(
        \MCInst_MC0_r1Inst_XORInst_0_1_n5 ), .B(
        \MCInst_MC0_r1Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[45]) );
  XNOR2_X1 \MCInst_MC0_r1Inst_XORInst_0_1_U2  ( .A(\MCInst_MC0_v3_1 [1]), .B(
        \MCInst_MC0_v2_1 [1]), .ZN(\MCInst_MC0_r1Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \MCInst_MC0_r1Inst_XORInst_0_1_U1  ( .A(\MCInst_MC0_v0_1 [1]), .B(
        \MCInst_MC0_v1_1 [1]), .Z(\MCInst_MC0_r1Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \MCInst_MC0_r1Inst_XORInst_0_2_U3  ( .A(
        \MCInst_MC0_r1Inst_XORInst_0_2_n5 ), .B(
        \MCInst_MC0_r1Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[46]) );
  XNOR2_X1 \MCInst_MC0_r1Inst_XORInst_0_2_U2  ( .A(\MCInst_MC0_v3_1 [2]), .B(
        \MCInst_MC0_v2_1 [2]), .ZN(\MCInst_MC0_r1Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \MCInst_MC0_r1Inst_XORInst_0_2_U1  ( .A(\MCInst_MC0_v0_1 [2]), .B(
        \MCInst_MC0_v1_1 [2]), .Z(\MCInst_MC0_r1Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \MCInst_MC0_r1Inst_XORInst_0_3_U3  ( .A(
        \MCInst_MC0_r1Inst_XORInst_0_3_n5 ), .B(
        \MCInst_MC0_r1Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[47]) );
  XNOR2_X1 \MCInst_MC0_r1Inst_XORInst_0_3_U2  ( .A(\MCInst_MC0_v3_1 [3]), .B(
        \MCInst_MC0_v2_1 [3]), .ZN(\MCInst_MC0_r1Inst_XORInst_0_3_n4 ) );
  XOR2_X1 \MCInst_MC0_r1Inst_XORInst_0_3_U1  ( .A(\MCInst_MC0_v0_1 [3]), .B(
        \MCInst_MC0_v1_1 [3]), .Z(\MCInst_MC0_r1Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 \MCInst_MC0_r2Inst_XORInst_0_0_U3  ( .A(
        \MCInst_MC0_r2Inst_XORInst_0_0_n5 ), .B(
        \MCInst_MC0_r2Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[28]) );
  XNOR2_X1 \MCInst_MC0_r2Inst_XORInst_0_0_U2  ( .A(\MCInst_MC0_v3_2 [0]), .B(
        \MCInst_MC0_v2_2 [0]), .ZN(\MCInst_MC0_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \MCInst_MC0_r2Inst_XORInst_0_0_U1  ( .A(\MCInst_MC0_v0_2 [0]), .B(
        \MCInst_MC0_v1_2 [0]), .Z(\MCInst_MC0_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \MCInst_MC0_r2Inst_XORInst_0_1_U3  ( .A(
        \MCInst_MC0_r2Inst_XORInst_0_1_n5 ), .B(
        \MCInst_MC0_r2Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[29]) );
  XNOR2_X1 \MCInst_MC0_r2Inst_XORInst_0_1_U2  ( .A(\MCInst_MC0_v3_0 [3]), .B(
        \MCInst_MC0_v2_2 [1]), .ZN(\MCInst_MC0_r2Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \MCInst_MC0_r2Inst_XORInst_0_1_U1  ( .A(\MCInst_MC0_v0_2 [1]), .B(
        \MCInst_MC0_v1_2 [1]), .Z(\MCInst_MC0_r2Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \MCInst_MC0_r2Inst_XORInst_0_2_U3  ( .A(
        \MCInst_MC0_r2Inst_XORInst_0_2_n5 ), .B(
        \MCInst_MC0_r2Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[30]) );
  XNOR2_X1 \MCInst_MC0_r2Inst_XORInst_0_2_U2  ( .A(\Red_MCInst_MC0_v3_1 [2]), 
        .B(\MCInst_MC0_v2_2 [2]), .ZN(\MCInst_MC0_r2Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \MCInst_MC0_r2Inst_XORInst_0_2_U1  ( .A(\MCInst_MC0_v0_2 [2]), .B(
        \MCInst_MC0_v1_2 [2]), .Z(\MCInst_MC0_r2Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \MCInst_MC0_r2Inst_XORInst_0_3_U3  ( .A(
        \MCInst_MC0_r2Inst_XORInst_0_3_n5 ), .B(
        \MCInst_MC0_r2Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[31]) );
  XNOR2_X1 \MCInst_MC0_r2Inst_XORInst_0_3_U2  ( .A(\MCInst_MC0_v3_2 [3]), .B(
        \MCInst_MC0_v2_2 [3]), .ZN(\MCInst_MC0_r2Inst_XORInst_0_3_n4 ) );
  XOR2_X1 \MCInst_MC0_r2Inst_XORInst_0_3_U1  ( .A(\MCInst_MC0_v0_2 [3]), .B(
        \MCInst_MC0_v1_2 [3]), .Z(\MCInst_MC0_r2Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 \MCInst_MC0_r3Inst_XORInst_0_0_U3  ( .A(
        \MCInst_MC0_r3Inst_XORInst_0_0_n5 ), .B(
        \MCInst_MC0_r3Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[12]) );
  XNOR2_X1 \MCInst_MC0_r3Inst_XORInst_0_0_U2  ( .A(\MCInst_MC0_v3_3 [0]), .B(
        \MCInst_MC0_v2_3 [0]), .ZN(\MCInst_MC0_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \MCInst_MC0_r3Inst_XORInst_0_0_U1  ( .A(\Red_MCInst_MC0_v0_1 [0]), 
        .B(\Red_MCInst_MC0_v1_1 [2]), .Z(\MCInst_MC0_r3Inst_XORInst_0_0_n5 )
         );
  XNOR2_X1 \MCInst_MC0_r3Inst_XORInst_0_1_U3  ( .A(
        \MCInst_MC0_r3Inst_XORInst_0_1_n5 ), .B(
        \MCInst_MC0_r3Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[13]) );
  XNOR2_X1 \MCInst_MC0_r3Inst_XORInst_0_1_U2  ( .A(\MCInst_MC0_v3_3 [1]), .B(
        \Red_MCInst_MC0_v2_1 [1]), .ZN(\MCInst_MC0_r3Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \MCInst_MC0_r3Inst_XORInst_0_1_U1  ( .A(\MCInst_MC0_v0_3 [1]), .B(
        \MCInst_MC0_v1_3 [1]), .Z(\MCInst_MC0_r3Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \MCInst_MC0_r3Inst_XORInst_0_2_U3  ( .A(
        \MCInst_MC0_r3Inst_XORInst_0_2_n5 ), .B(
        \MCInst_MC0_r3Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[14]) );
  XNOR2_X1 \MCInst_MC0_r3Inst_XORInst_0_2_U2  ( .A(\MCInst_MC0_v3_3 [2]), .B(
        \MCInst_MC0_v2_3 [2]), .ZN(\MCInst_MC0_r3Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \MCInst_MC0_r3Inst_XORInst_0_2_U1  ( .A(\Red_MCInst_MC0_v0_2 [2]), 
        .B(\Red_MCInst_MC0_v1_2 [1]), .Z(\MCInst_MC0_r3Inst_XORInst_0_2_n5 )
         );
  XNOR2_X1 \MCInst_MC0_r3Inst_XORInst_0_3_U3  ( .A(
        \MCInst_MC0_r3Inst_XORInst_0_3_n5 ), .B(
        \MCInst_MC0_r3Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[15]) );
  XNOR2_X1 \MCInst_MC0_r3Inst_XORInst_0_3_U2  ( .A(\MCInst_MC0_v3_3 [3]), .B(
        \MCInst_MC0_v2_3 [3]), .ZN(\MCInst_MC0_r3Inst_XORInst_0_3_n4 ) );
  XOR2_X1 \MCInst_MC0_r3Inst_XORInst_0_3_U1  ( .A(\MCInst_MC0_v0_3 [3]), .B(
        \MCInst_MC0_v1_3 [3]), .Z(\MCInst_MC0_r3Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 \MCInst_MC1_v0_2Inst_0_U4  ( .A(\MCInst_MC1_v0_2Inst_0_n2 ), .B(
        \Red_MCInst_MC1_v0_2 [2]), .ZN(\MCInst_MC1_v0_2 [0]) );
  XNOR2_X1 \MCInst_MC1_v0_2Inst_0_U3  ( .A(\Red_MCInst_MC1_v0_1 [0]), .B(
        \Red_MCInst_MC1_v0_0 [0]), .ZN(\MCInst_MC1_v0_2Inst_0_n2 ) );
  XOR2_X1 \MCInst_MC1_v1_1Inst_0_U3  ( .A(\MCInst_MC1_v1_3 [3]), .B(
        \Red_MCInst_MC1_v1_1 [2]), .Z(\MCInst_MC1_v1_1 [0]) );
  XNOR2_X1 \MCInst_MC1_v1_2Inst_0_U4  ( .A(\MCInst_MC1_v1_2Inst_0_n2 ), .B(
        \MCInst_MC1_v1_3 [3]), .ZN(\MCInst_MC1_v1_2 [0]) );
  XNOR2_X1 \MCInst_MC1_v1_2Inst_0_U3  ( .A(\Red_MCInst_MC1_v1_1 [2]), .B(
        \Red_MCInst_MC1_v1_2 [1]), .ZN(\MCInst_MC1_v1_2Inst_0_n2 ) );
  XOR2_X1 \MCInst_MC1_v2_1Inst_0_U3  ( .A(\Red_MCInst_MC1_v2_1 [1]), .B(
        \MCInst_MC1_v2_0 [3]), .Z(\MCInst_MC1_v2_1 [0]) );
  XOR2_X1 \MCInst_MC1_v2_2Inst_0_U3  ( .A(\MCInst_MC1_v2_0 [2]), .B(
        \Red_MCInst_MC1_v2_2 [1]), .Z(\MCInst_MC1_v2_2 [0]) );
  XNOR2_X1 \MCInst_MC1_v2_3Inst_0_U5  ( .A(\MCInst_MC1_v2_3Inst_0_n4 ), .B(
        \MCInst_MC1_v2_3Inst_0_n3 ), .ZN(\MCInst_MC1_v2_3 [0]) );
  XNOR2_X1 \MCInst_MC1_v2_3Inst_0_U4  ( .A(\MCInst_MC1_v2_0 [2]), .B(
        \Red_MCInst_MC1_v2_1 [1]), .ZN(\MCInst_MC1_v2_3Inst_0_n3 ) );
  XOR2_X1 \MCInst_MC1_v2_3Inst_0_U3  ( .A(\MCInst_MC1_v2_0 [3]), .B(
        \Red_MCInst_MC1_v2_2 [1]), .Z(\MCInst_MC1_v2_3Inst_0_n4 ) );
  XOR2_X1 \MCInst_MC1_v3_1Inst_0_U3  ( .A(\MCInst_MC1_v3_0 [3]), .B(
        \Red_MCInst_MC1_v3_1 [2]), .Z(\MCInst_MC1_v3_1 [0]) );
  XOR2_X1 \MCInst_MC1_v3_2Inst_0_U3  ( .A(\MCInst_MC1_v3_2 [3]), .B(
        \Red_MCInst_MC1_v3_3 [2]), .Z(\MCInst_MC1_v3_2 [0]) );
  XNOR2_X1 \MCInst_MC1_v3_3Inst_0_U4  ( .A(\MCInst_MC1_v3_3Inst_0_n2 ), .B(
        \Red_MCInst_MC1_v3_3 [2]), .ZN(\MCInst_MC1_v3_3 [0]) );
  XNOR2_X1 \MCInst_MC1_v3_3Inst_0_U3  ( .A(\Red_MCInst_MC1_v3_1 [2]), .B(
        \MCInst_MC1_v3_2 [3]), .ZN(\MCInst_MC1_v3_3Inst_0_n2 ) );
  XOR2_X1 \MCInst_MC1_v0_0Inst_1_U3  ( .A(\MCInst_MC1_v0_3 [3]), .B(
        \Red_MCInst_MC1_v0_1 [0]), .Z(\MCInst_MC1_v0_0 [1]) );
  XOR2_X1 \MCInst_MC1_v0_1Inst_1_U3  ( .A(\Red_MCInst_MC1_v0_2 [2]), .B(
        \MCInst_MC1_v0_3 [3]), .Z(\MCInst_MC1_v0_1 [1]) );
  XNOR2_X1 \MCInst_MC1_v0_2Inst_1_U4  ( .A(\MCInst_MC1_v0_2Inst_1_n2 ), .B(
        \MCInst_MC1_v0_3 [3]), .ZN(\MCInst_MC1_v0_2 [1]) );
  XNOR2_X1 \MCInst_MC1_v0_2Inst_1_U3  ( .A(\Red_MCInst_MC1_v0_1 [0]), .B(
        \Red_MCInst_MC1_v0_0 [0]), .ZN(\MCInst_MC1_v0_2Inst_1_n2 ) );
  XOR2_X1 \MCInst_MC1_v0_3Inst_1_U3  ( .A(\Red_MCInst_MC1_v0_0 [0]), .B(
        \Red_MCInst_MC1_v0_1 [0]), .Z(\MCInst_MC1_v0_3 [1]) );
  XOR2_X1 \MCInst_MC1_v1_1Inst_1_U3  ( .A(\MCInst_MC1_v1_0 [0]), .B(
        \MCInst_MC1_v1_3 [3]), .Z(\MCInst_MC1_v1_1 [1]) );
  XOR2_X1 \MCInst_MC1_v1_2Inst_1_U3  ( .A(\MCInst_MC1_v1_0 [0]), .B(
        \Red_MCInst_MC1_v1_2 [1]), .Z(\MCInst_MC1_v1_2 [1]) );
  XOR2_X1 \MCInst_MC1_v1_3Inst_1_U3  ( .A(\MCInst_MC1_v1_0 [0]), .B(
        \Red_MCInst_MC1_v1_1 [2]), .Z(\MCInst_MC1_v1_3 [1]) );
  XOR2_X1 \MCInst_MC1_v2_0Inst_1_U3  ( .A(\Red_MCInst_MC1_v2_1 [1]), .B(
        \Red_MCInst_MC1_v2_2 [1]), .Z(\MCInst_MC1_v2_0 [1]) );
  XNOR2_X1 \MCInst_MC1_v2_1Inst_1_U4  ( .A(\MCInst_MC1_v2_1Inst_1_n2 ), .B(
        \MCInst_MC1_v2_0 [3]), .ZN(\MCInst_MC1_v2_1 [1]) );
  XNOR2_X1 \MCInst_MC1_v2_1Inst_1_U3  ( .A(\Red_MCInst_MC1_v2_2 [1]), .B(
        \MCInst_MC1_v2_0 [2]), .ZN(\MCInst_MC1_v2_1Inst_1_n2 ) );
  XNOR2_X1 \MCInst_MC1_v2_2Inst_1_U5  ( .A(\MCInst_MC1_v2_2Inst_1_n4 ), .B(
        \MCInst_MC1_v2_2Inst_1_n3 ), .ZN(\MCInst_MC1_v2_2 [1]) );
  XNOR2_X1 \MCInst_MC1_v2_2Inst_1_U4  ( .A(\MCInst_MC1_v2_0 [2]), .B(
        \Red_MCInst_MC1_v2_1 [1]), .ZN(\MCInst_MC1_v2_2Inst_1_n3 ) );
  XOR2_X1 \MCInst_MC1_v2_2Inst_1_U3  ( .A(\MCInst_MC1_v2_0 [3]), .B(
        \Red_MCInst_MC1_v2_2 [1]), .Z(\MCInst_MC1_v2_2Inst_1_n4 ) );
  XOR2_X1 \MCInst_MC1_v3_0Inst_1_U3  ( .A(\MCInst_MC1_v3_2 [3]), .B(
        \Red_MCInst_MC1_v3_1 [2]), .Z(\MCInst_MC1_v3_0 [1]) );
  XOR2_X1 \MCInst_MC1_v3_1Inst_1_U3  ( .A(\MCInst_MC1_v3_2 [3]), .B(
        \MCInst_MC1_v3_0 [3]), .Z(\MCInst_MC1_v3_1 [1]) );
  XNOR2_X1 \MCInst_MC1_v3_3Inst_1_U4  ( .A(\MCInst_MC1_v3_3Inst_1_n2 ), .B(
        \MCInst_MC1_v3_0 [3]), .ZN(\MCInst_MC1_v3_3 [1]) );
  XNOR2_X1 \MCInst_MC1_v3_3Inst_1_U3  ( .A(\Red_MCInst_MC1_v3_1 [2]), .B(
        \MCInst_MC1_v3_2 [3]), .ZN(\MCInst_MC1_v3_3Inst_1_n2 ) );
  XOR2_X1 \MCInst_MC1_v0_0Inst_2_U3  ( .A(\Red_MCInst_MC1_v0_0 [0]), .B(
        \Red_MCInst_MC1_v0_1 [0]), .Z(\MCInst_MC1_v0_0 [2]) );
  XOR2_X1 \MCInst_MC1_v0_1Inst_2_U3  ( .A(\MCInst_MC1_v0_3 [3]), .B(
        \Red_MCInst_MC1_v0_1 [0]), .Z(\MCInst_MC1_v0_1 [2]) );
  XOR2_X1 \MCInst_MC1_v0_2Inst_2_U3  ( .A(\Red_MCInst_MC1_v0_2 [2]), .B(
        \Red_MCInst_MC1_v0_1 [0]), .Z(\MCInst_MC1_v0_2 [2]) );
  XNOR2_X1 \MCInst_MC1_v1_1Inst_2_U4  ( .A(\MCInst_MC1_v1_1Inst_2_n2 ), .B(
        \Red_MCInst_MC1_v1_2 [1]), .ZN(\MCInst_MC1_v1_1 [2]) );
  XNOR2_X1 \MCInst_MC1_v1_1Inst_2_U3  ( .A(\Red_MCInst_MC1_v1_1 [2]), .B(
        \MCInst_MC1_v1_0 [0]), .ZN(\MCInst_MC1_v1_1Inst_2_n2 ) );
  XNOR2_X1 \MCInst_MC1_v1_2Inst_2_U4  ( .A(\MCInst_MC1_v1_2Inst_2_n2 ), .B(
        \Red_MCInst_MC1_v1_2 [1]), .ZN(\MCInst_MC1_v1_2 [2]) );
  XNOR2_X1 \MCInst_MC1_v1_2Inst_2_U3  ( .A(\MCInst_MC1_v1_3 [3]), .B(
        \MCInst_MC1_v1_0 [0]), .ZN(\MCInst_MC1_v1_2Inst_2_n2 ) );
  XNOR2_X1 \MCInst_MC1_v2_1Inst_2_U4  ( .A(\MCInst_MC1_v2_1Inst_2_n2 ), .B(
        \MCInst_MC1_v2_0 [3]), .ZN(\MCInst_MC1_v2_1 [2]) );
  XNOR2_X1 \MCInst_MC1_v2_1Inst_2_U3  ( .A(\Red_MCInst_MC1_v2_2 [1]), .B(
        \Red_MCInst_MC1_v2_1 [1]), .ZN(\MCInst_MC1_v2_1Inst_2_n2 ) );
  XNOR2_X1 \MCInst_MC1_v2_2Inst_2_U4  ( .A(\MCInst_MC1_v2_2Inst_2_n2 ), .B(
        \MCInst_MC1_v2_0 [3]), .ZN(\MCInst_MC1_v2_2 [2]) );
  XNOR2_X1 \MCInst_MC1_v2_2Inst_2_U3  ( .A(\Red_MCInst_MC1_v2_2 [1]), .B(
        \MCInst_MC1_v2_0 [2]), .ZN(\MCInst_MC1_v2_2Inst_2_n2 ) );
  XOR2_X1 \MCInst_MC1_v2_3Inst_2_U3  ( .A(\Red_MCInst_MC1_v2_1 [1]), .B(
        \MCInst_MC1_v2_0 [2]), .Z(\MCInst_MC1_v2_3 [2]) );
  XNOR2_X1 \MCInst_MC1_v3_1Inst_2_U4  ( .A(\MCInst_MC1_v3_1Inst_2_n2 ), .B(
        \Red_MCInst_MC1_v3_3 [2]), .ZN(\MCInst_MC1_v3_1 [2]) );
  XNOR2_X1 \MCInst_MC1_v3_1Inst_2_U3  ( .A(\Red_MCInst_MC1_v3_1 [2]), .B(
        \MCInst_MC1_v3_2 [3]), .ZN(\MCInst_MC1_v3_1Inst_2_n2 ) );
  XOR2_X1 \MCInst_MC1_v3_3Inst_2_U3  ( .A(\Red_MCInst_MC1_v3_3 [2]), .B(
        \Red_MCInst_MC1_v3_1 [2]), .Z(\MCInst_MC1_v3_3 [2]) );
  XOR2_X1 \MCInst_MC1_v0_1Inst_3_U3  ( .A(\Red_MCInst_MC1_v0_0 [0]), .B(
        \Red_MCInst_MC1_v0_1 [0]), .Z(\MCInst_MC1_v0_1 [3]) );
  XOR2_X1 \MCInst_MC1_v0_2Inst_3_U3  ( .A(\Red_MCInst_MC1_v0_0 [0]), .B(
        \MCInst_MC1_v0_3 [3]), .Z(\MCInst_MC1_v0_2 [3]) );
  XOR2_X1 \MCInst_MC1_v1_1Inst_3_U3  ( .A(\Red_MCInst_MC1_v1_2 [1]), .B(
        \MCInst_MC1_v1_3 [3]), .Z(\MCInst_MC1_v1_1 [3]) );
  XNOR2_X1 \MCInst_MC1_v1_2Inst_3_U5  ( .A(\MCInst_MC1_v1_2Inst_3_n4 ), .B(
        \MCInst_MC1_v1_2Inst_3_n3 ), .ZN(\MCInst_MC1_v1_2 [3]) );
  XNOR2_X1 \MCInst_MC1_v1_2Inst_3_U4  ( .A(\Red_MCInst_MC1_v1_2 [1]), .B(
        \MCInst_MC1_v1_0 [0]), .ZN(\MCInst_MC1_v1_2Inst_3_n3 ) );
  XOR2_X1 \MCInst_MC1_v1_2Inst_3_U3  ( .A(\MCInst_MC1_v1_3 [3]), .B(
        \Red_MCInst_MC1_v1_1 [2]), .Z(\MCInst_MC1_v1_2Inst_3_n4 ) );
  XOR2_X1 \MCInst_MC1_v2_1Inst_3_U3  ( .A(\MCInst_MC1_v2_0 [2]), .B(
        \Red_MCInst_MC1_v2_2 [1]), .Z(\MCInst_MC1_v2_1 [3]) );
  XNOR2_X1 \MCInst_MC1_v2_2Inst_3_U4  ( .A(\MCInst_MC1_v2_2Inst_3_n2 ), .B(
        \MCInst_MC1_v2_0 [3]), .ZN(\MCInst_MC1_v2_2 [3]) );
  XNOR2_X1 \MCInst_MC1_v2_2Inst_3_U3  ( .A(\Red_MCInst_MC1_v2_2 [1]), .B(
        \Red_MCInst_MC1_v2_1 [1]), .ZN(\MCInst_MC1_v2_2Inst_3_n2 ) );
  XNOR2_X1 \MCInst_MC1_v2_3Inst_3_U4  ( .A(\MCInst_MC1_v2_3Inst_3_n2 ), .B(
        \MCInst_MC1_v2_0 [2]), .ZN(\MCInst_MC1_v2_3 [3]) );
  XNOR2_X1 \MCInst_MC1_v2_3Inst_3_U3  ( .A(\MCInst_MC1_v2_0 [3]), .B(
        \Red_MCInst_MC1_v2_1 [1]), .ZN(\MCInst_MC1_v2_3Inst_3_n2 ) );
  XOR2_X1 \MCInst_MC1_v3_1Inst_3_U3  ( .A(\Red_MCInst_MC1_v3_3 [2]), .B(
        \MCInst_MC1_v3_0 [3]), .Z(\MCInst_MC1_v3_1 [3]) );
  XOR2_X1 \MCInst_MC1_v3_3Inst_3_U3  ( .A(\MCInst_MC1_v3_2 [3]), .B(
        \MCInst_MC1_v3_0 [3]), .Z(\MCInst_MC1_v3_3 [3]) );
  XNOR2_X1 \MCInst_MC1_r0Inst_XORInst_0_0_U3  ( .A(
        \MCInst_MC1_r0Inst_XORInst_0_0_n5 ), .B(
        \MCInst_MC1_r0Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[56]) );
  XNOR2_X1 \MCInst_MC1_r0Inst_XORInst_0_0_U2  ( .A(\Red_MCInst_MC1_v3_1 [2]), 
        .B(\Red_MCInst_MC1_v2_2 [1]), .ZN(\MCInst_MC1_r0Inst_XORInst_0_0_n4 )
         );
  XOR2_X1 \MCInst_MC1_r0Inst_XORInst_0_0_U1  ( .A(\MCInst_MC1_v0_3 [3]), .B(
        \MCInst_MC1_v1_0 [0]), .Z(\MCInst_MC1_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \MCInst_MC1_r0Inst_XORInst_0_1_U3  ( .A(
        \MCInst_MC1_r0Inst_XORInst_0_1_n5 ), .B(
        \MCInst_MC1_r0Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[57]) );
  XNOR2_X1 \MCInst_MC1_r0Inst_XORInst_0_1_U2  ( .A(\MCInst_MC1_v3_0 [1]), .B(
        \MCInst_MC1_v2_0 [1]), .ZN(\MCInst_MC1_r0Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \MCInst_MC1_r0Inst_XORInst_0_1_U1  ( .A(\MCInst_MC1_v0_0 [1]), .B(
        \Red_MCInst_MC1_v1_2 [1]), .Z(\MCInst_MC1_r0Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \MCInst_MC1_r0Inst_XORInst_0_2_U3  ( .A(
        \MCInst_MC1_r0Inst_XORInst_0_2_n5 ), .B(
        \MCInst_MC1_r0Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[58]) );
  XNOR2_X1 \MCInst_MC1_r0Inst_XORInst_0_2_U2  ( .A(\Red_MCInst_MC1_v3_3 [2]), 
        .B(\MCInst_MC1_v2_0 [2]), .ZN(\MCInst_MC1_r0Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \MCInst_MC1_r0Inst_XORInst_0_2_U1  ( .A(\MCInst_MC1_v0_0 [2]), .B(
        \MCInst_MC1_v1_3 [3]), .Z(\MCInst_MC1_r0Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \MCInst_MC1_r0Inst_XORInst_0_3_U3  ( .A(
        \MCInst_MC1_r0Inst_XORInst_0_3_n5 ), .B(
        \MCInst_MC1_r0Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[59]) );
  XNOR2_X1 \MCInst_MC1_r0Inst_XORInst_0_3_U2  ( .A(\MCInst_MC1_v3_0 [3]), .B(
        \MCInst_MC1_v2_0 [3]), .ZN(\MCInst_MC1_r0Inst_XORInst_0_3_n4 ) );
  XOR2_X1 \MCInst_MC1_r0Inst_XORInst_0_3_U1  ( .A(\Red_MCInst_MC1_v0_2 [2]), 
        .B(\Red_MCInst_MC1_v1_1 [2]), .Z(\MCInst_MC1_r0Inst_XORInst_0_3_n5 )
         );
  XNOR2_X1 \MCInst_MC1_r1Inst_XORInst_0_0_U3  ( .A(
        \MCInst_MC1_r1Inst_XORInst_0_0_n5 ), .B(
        \MCInst_MC1_r1Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[40]) );
  XNOR2_X1 \MCInst_MC1_r1Inst_XORInst_0_0_U2  ( .A(\MCInst_MC1_v3_1 [0]), .B(
        \MCInst_MC1_v2_1 [0]), .ZN(\MCInst_MC1_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \MCInst_MC1_r1Inst_XORInst_0_0_U1  ( .A(\Red_MCInst_MC1_v0_2 [2]), 
        .B(\MCInst_MC1_v1_1 [0]), .Z(\MCInst_MC1_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \MCInst_MC1_r1Inst_XORInst_0_1_U3  ( .A(
        \MCInst_MC1_r1Inst_XORInst_0_1_n5 ), .B(
        \MCInst_MC1_r1Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[41]) );
  XNOR2_X1 \MCInst_MC1_r1Inst_XORInst_0_1_U2  ( .A(\MCInst_MC1_v3_1 [1]), .B(
        \MCInst_MC1_v2_1 [1]), .ZN(\MCInst_MC1_r1Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \MCInst_MC1_r1Inst_XORInst_0_1_U1  ( .A(\MCInst_MC1_v0_1 [1]), .B(
        \MCInst_MC1_v1_1 [1]), .Z(\MCInst_MC1_r1Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \MCInst_MC1_r1Inst_XORInst_0_2_U3  ( .A(
        \MCInst_MC1_r1Inst_XORInst_0_2_n5 ), .B(
        \MCInst_MC1_r1Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[42]) );
  XNOR2_X1 \MCInst_MC1_r1Inst_XORInst_0_2_U2  ( .A(\MCInst_MC1_v3_1 [2]), .B(
        \MCInst_MC1_v2_1 [2]), .ZN(\MCInst_MC1_r1Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \MCInst_MC1_r1Inst_XORInst_0_2_U1  ( .A(\MCInst_MC1_v0_1 [2]), .B(
        \MCInst_MC1_v1_1 [2]), .Z(\MCInst_MC1_r1Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \MCInst_MC1_r1Inst_XORInst_0_3_U3  ( .A(
        \MCInst_MC1_r1Inst_XORInst_0_3_n5 ), .B(
        \MCInst_MC1_r1Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[43]) );
  XNOR2_X1 \MCInst_MC1_r1Inst_XORInst_0_3_U2  ( .A(\MCInst_MC1_v3_1 [3]), .B(
        \MCInst_MC1_v2_1 [3]), .ZN(\MCInst_MC1_r1Inst_XORInst_0_3_n4 ) );
  XOR2_X1 \MCInst_MC1_r1Inst_XORInst_0_3_U1  ( .A(\MCInst_MC1_v0_1 [3]), .B(
        \MCInst_MC1_v1_1 [3]), .Z(\MCInst_MC1_r1Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 \MCInst_MC1_r2Inst_XORInst_0_0_U3  ( .A(
        \MCInst_MC1_r2Inst_XORInst_0_0_n5 ), .B(
        \MCInst_MC1_r2Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[24]) );
  XNOR2_X1 \MCInst_MC1_r2Inst_XORInst_0_0_U2  ( .A(\MCInst_MC1_v3_2 [0]), .B(
        \MCInst_MC1_v2_2 [0]), .ZN(\MCInst_MC1_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \MCInst_MC1_r2Inst_XORInst_0_0_U1  ( .A(\MCInst_MC1_v0_2 [0]), .B(
        \MCInst_MC1_v1_2 [0]), .Z(\MCInst_MC1_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \MCInst_MC1_r2Inst_XORInst_0_1_U3  ( .A(
        \MCInst_MC1_r2Inst_XORInst_0_1_n5 ), .B(
        \MCInst_MC1_r2Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[25]) );
  XNOR2_X1 \MCInst_MC1_r2Inst_XORInst_0_1_U2  ( .A(\MCInst_MC1_v3_0 [3]), .B(
        \MCInst_MC1_v2_2 [1]), .ZN(\MCInst_MC1_r2Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \MCInst_MC1_r2Inst_XORInst_0_1_U1  ( .A(\MCInst_MC1_v0_2 [1]), .B(
        \MCInst_MC1_v1_2 [1]), .Z(\MCInst_MC1_r2Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \MCInst_MC1_r2Inst_XORInst_0_2_U3  ( .A(
        \MCInst_MC1_r2Inst_XORInst_0_2_n5 ), .B(
        \MCInst_MC1_r2Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[26]) );
  XNOR2_X1 \MCInst_MC1_r2Inst_XORInst_0_2_U2  ( .A(\Red_MCInst_MC1_v3_1 [2]), 
        .B(\MCInst_MC1_v2_2 [2]), .ZN(\MCInst_MC1_r2Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \MCInst_MC1_r2Inst_XORInst_0_2_U1  ( .A(\MCInst_MC1_v0_2 [2]), .B(
        \MCInst_MC1_v1_2 [2]), .Z(\MCInst_MC1_r2Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \MCInst_MC1_r2Inst_XORInst_0_3_U3  ( .A(
        \MCInst_MC1_r2Inst_XORInst_0_3_n5 ), .B(
        \MCInst_MC1_r2Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[27]) );
  XNOR2_X1 \MCInst_MC1_r2Inst_XORInst_0_3_U2  ( .A(\MCInst_MC1_v3_2 [3]), .B(
        \MCInst_MC1_v2_2 [3]), .ZN(\MCInst_MC1_r2Inst_XORInst_0_3_n4 ) );
  XOR2_X1 \MCInst_MC1_r2Inst_XORInst_0_3_U1  ( .A(\MCInst_MC1_v0_2 [3]), .B(
        \MCInst_MC1_v1_2 [3]), .Z(\MCInst_MC1_r2Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 \MCInst_MC1_r3Inst_XORInst_0_0_U3  ( .A(
        \MCInst_MC1_r3Inst_XORInst_0_0_n5 ), .B(
        \MCInst_MC1_r3Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[8]) );
  XNOR2_X1 \MCInst_MC1_r3Inst_XORInst_0_0_U2  ( .A(\MCInst_MC1_v3_3 [0]), .B(
        \MCInst_MC1_v2_3 [0]), .ZN(\MCInst_MC1_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \MCInst_MC1_r3Inst_XORInst_0_0_U1  ( .A(\Red_MCInst_MC1_v0_1 [0]), 
        .B(\Red_MCInst_MC1_v1_1 [2]), .Z(\MCInst_MC1_r3Inst_XORInst_0_0_n5 )
         );
  XNOR2_X1 \MCInst_MC1_r3Inst_XORInst_0_1_U3  ( .A(
        \MCInst_MC1_r3Inst_XORInst_0_1_n5 ), .B(
        \MCInst_MC1_r3Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[9]) );
  XNOR2_X1 \MCInst_MC1_r3Inst_XORInst_0_1_U2  ( .A(\MCInst_MC1_v3_3 [1]), .B(
        \Red_MCInst_MC1_v2_1 [1]), .ZN(\MCInst_MC1_r3Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \MCInst_MC1_r3Inst_XORInst_0_1_U1  ( .A(\MCInst_MC1_v0_3 [1]), .B(
        \MCInst_MC1_v1_3 [1]), .Z(\MCInst_MC1_r3Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \MCInst_MC1_r3Inst_XORInst_0_2_U3  ( .A(
        \MCInst_MC1_r3Inst_XORInst_0_2_n5 ), .B(
        \MCInst_MC1_r3Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[10]) );
  XNOR2_X1 \MCInst_MC1_r3Inst_XORInst_0_2_U2  ( .A(\MCInst_MC1_v3_3 [2]), .B(
        \MCInst_MC1_v2_3 [2]), .ZN(\MCInst_MC1_r3Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \MCInst_MC1_r3Inst_XORInst_0_2_U1  ( .A(\Red_MCInst_MC1_v0_2 [2]), 
        .B(\Red_MCInst_MC1_v1_2 [1]), .Z(\MCInst_MC1_r3Inst_XORInst_0_2_n5 )
         );
  XNOR2_X1 \MCInst_MC1_r3Inst_XORInst_0_3_U3  ( .A(
        \MCInst_MC1_r3Inst_XORInst_0_3_n5 ), .B(
        \MCInst_MC1_r3Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[11]) );
  XNOR2_X1 \MCInst_MC1_r3Inst_XORInst_0_3_U2  ( .A(\MCInst_MC1_v3_3 [3]), .B(
        \MCInst_MC1_v2_3 [3]), .ZN(\MCInst_MC1_r3Inst_XORInst_0_3_n4 ) );
  XOR2_X1 \MCInst_MC1_r3Inst_XORInst_0_3_U1  ( .A(\MCInst_MC1_v0_3 [3]), .B(
        \MCInst_MC1_v1_3 [3]), .Z(\MCInst_MC1_r3Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 \MCInst_MC2_v0_2Inst_0_U4  ( .A(\MCInst_MC2_v0_2Inst_0_n2 ), .B(
        \Red_MCInst_MC2_v0_2 [2]), .ZN(\MCInst_MC2_v0_2 [0]) );
  XNOR2_X1 \MCInst_MC2_v0_2Inst_0_U3  ( .A(\Red_MCInst_MC2_v0_1 [0]), .B(
        \Red_MCInst_MC2_v0_0 [0]), .ZN(\MCInst_MC2_v0_2Inst_0_n2 ) );
  XOR2_X1 \MCInst_MC2_v1_1Inst_0_U3  ( .A(\MCInst_MC2_v1_3 [3]), .B(
        \Red_MCInst_MC2_v1_1 [2]), .Z(\MCInst_MC2_v1_1 [0]) );
  XNOR2_X1 \MCInst_MC2_v1_2Inst_0_U4  ( .A(\MCInst_MC2_v1_2Inst_0_n2 ), .B(
        \MCInst_MC2_v1_3 [3]), .ZN(\MCInst_MC2_v1_2 [0]) );
  XNOR2_X1 \MCInst_MC2_v1_2Inst_0_U3  ( .A(\Red_MCInst_MC2_v1_1 [2]), .B(
        \Red_MCInst_MC2_v1_2 [1]), .ZN(\MCInst_MC2_v1_2Inst_0_n2 ) );
  XOR2_X1 \MCInst_MC2_v2_1Inst_0_U3  ( .A(\Red_MCInst_MC2_v2_1 [1]), .B(
        \MCInst_MC2_v2_0 [3]), .Z(\MCInst_MC2_v2_1 [0]) );
  XOR2_X1 \MCInst_MC2_v2_2Inst_0_U3  ( .A(\MCInst_MC2_v2_0 [2]), .B(
        \Red_MCInst_MC2_v2_2 [1]), .Z(\MCInst_MC2_v2_2 [0]) );
  XNOR2_X1 \MCInst_MC2_v2_3Inst_0_U5  ( .A(\MCInst_MC2_v2_3Inst_0_n4 ), .B(
        \MCInst_MC2_v2_3Inst_0_n3 ), .ZN(\MCInst_MC2_v2_3 [0]) );
  XNOR2_X1 \MCInst_MC2_v2_3Inst_0_U4  ( .A(\MCInst_MC2_v2_0 [2]), .B(
        \Red_MCInst_MC2_v2_1 [1]), .ZN(\MCInst_MC2_v2_3Inst_0_n3 ) );
  XOR2_X1 \MCInst_MC2_v2_3Inst_0_U3  ( .A(\MCInst_MC2_v2_0 [3]), .B(
        \Red_MCInst_MC2_v2_2 [1]), .Z(\MCInst_MC2_v2_3Inst_0_n4 ) );
  XOR2_X1 \MCInst_MC2_v3_1Inst_0_U3  ( .A(\MCInst_MC2_v3_0 [3]), .B(
        \Red_MCInst_MC2_v3_1 [2]), .Z(\MCInst_MC2_v3_1 [0]) );
  XOR2_X1 \MCInst_MC2_v3_2Inst_0_U3  ( .A(\MCInst_MC2_v3_2 [3]), .B(
        \Red_MCInst_MC2_v3_3 [2]), .Z(\MCInst_MC2_v3_2 [0]) );
  XNOR2_X1 \MCInst_MC2_v3_3Inst_0_U4  ( .A(\MCInst_MC2_v3_3Inst_0_n2 ), .B(
        \Red_MCInst_MC2_v3_3 [2]), .ZN(\MCInst_MC2_v3_3 [0]) );
  XNOR2_X1 \MCInst_MC2_v3_3Inst_0_U3  ( .A(\Red_MCInst_MC2_v3_1 [2]), .B(
        \MCInst_MC2_v3_2 [3]), .ZN(\MCInst_MC2_v3_3Inst_0_n2 ) );
  XOR2_X1 \MCInst_MC2_v0_0Inst_1_U3  ( .A(\MCInst_MC2_v0_3 [3]), .B(
        \Red_MCInst_MC2_v0_1 [0]), .Z(\MCInst_MC2_v0_0 [1]) );
  XOR2_X1 \MCInst_MC2_v0_1Inst_1_U3  ( .A(\Red_MCInst_MC2_v0_2 [2]), .B(
        \MCInst_MC2_v0_3 [3]), .Z(\MCInst_MC2_v0_1 [1]) );
  XNOR2_X1 \MCInst_MC2_v0_2Inst_1_U4  ( .A(\MCInst_MC2_v0_2Inst_1_n2 ), .B(
        \MCInst_MC2_v0_3 [3]), .ZN(\MCInst_MC2_v0_2 [1]) );
  XNOR2_X1 \MCInst_MC2_v0_2Inst_1_U3  ( .A(\Red_MCInst_MC2_v0_1 [0]), .B(
        \Red_MCInst_MC2_v0_0 [0]), .ZN(\MCInst_MC2_v0_2Inst_1_n2 ) );
  XOR2_X1 \MCInst_MC2_v0_3Inst_1_U3  ( .A(\Red_MCInst_MC2_v0_0 [0]), .B(
        \Red_MCInst_MC2_v0_1 [0]), .Z(\MCInst_MC2_v0_3 [1]) );
  XOR2_X1 \MCInst_MC2_v1_1Inst_1_U3  ( .A(\MCInst_MC2_v1_0 [0]), .B(
        \MCInst_MC2_v1_3 [3]), .Z(\MCInst_MC2_v1_1 [1]) );
  XOR2_X1 \MCInst_MC2_v1_2Inst_1_U3  ( .A(\MCInst_MC2_v1_0 [0]), .B(
        \Red_MCInst_MC2_v1_2 [1]), .Z(\MCInst_MC2_v1_2 [1]) );
  XOR2_X1 \MCInst_MC2_v1_3Inst_1_U3  ( .A(\MCInst_MC2_v1_0 [0]), .B(
        \Red_MCInst_MC2_v1_1 [2]), .Z(\MCInst_MC2_v1_3 [1]) );
  XOR2_X1 \MCInst_MC2_v2_0Inst_1_U3  ( .A(\Red_MCInst_MC2_v2_1 [1]), .B(
        \Red_MCInst_MC2_v2_2 [1]), .Z(\MCInst_MC2_v2_0 [1]) );
  XNOR2_X1 \MCInst_MC2_v2_1Inst_1_U4  ( .A(\MCInst_MC2_v2_1Inst_1_n2 ), .B(
        \MCInst_MC2_v2_0 [3]), .ZN(\MCInst_MC2_v2_1 [1]) );
  XNOR2_X1 \MCInst_MC2_v2_1Inst_1_U3  ( .A(\Red_MCInst_MC2_v2_2 [1]), .B(
        \MCInst_MC2_v2_0 [2]), .ZN(\MCInst_MC2_v2_1Inst_1_n2 ) );
  XNOR2_X1 \MCInst_MC2_v2_2Inst_1_U5  ( .A(\MCInst_MC2_v2_2Inst_1_n4 ), .B(
        \MCInst_MC2_v2_2Inst_1_n3 ), .ZN(\MCInst_MC2_v2_2 [1]) );
  XNOR2_X1 \MCInst_MC2_v2_2Inst_1_U4  ( .A(\MCInst_MC2_v2_0 [2]), .B(
        \Red_MCInst_MC2_v2_1 [1]), .ZN(\MCInst_MC2_v2_2Inst_1_n3 ) );
  XOR2_X1 \MCInst_MC2_v2_2Inst_1_U3  ( .A(\MCInst_MC2_v2_0 [3]), .B(
        \Red_MCInst_MC2_v2_2 [1]), .Z(\MCInst_MC2_v2_2Inst_1_n4 ) );
  XOR2_X1 \MCInst_MC2_v3_0Inst_1_U3  ( .A(\MCInst_MC2_v3_2 [3]), .B(
        \Red_MCInst_MC2_v3_1 [2]), .Z(\MCInst_MC2_v3_0 [1]) );
  XOR2_X1 \MCInst_MC2_v3_1Inst_1_U3  ( .A(\MCInst_MC2_v3_2 [3]), .B(
        \MCInst_MC2_v3_0 [3]), .Z(\MCInst_MC2_v3_1 [1]) );
  XNOR2_X1 \MCInst_MC2_v3_3Inst_1_U4  ( .A(\MCInst_MC2_v3_3Inst_1_n2 ), .B(
        \MCInst_MC2_v3_0 [3]), .ZN(\MCInst_MC2_v3_3 [1]) );
  XNOR2_X1 \MCInst_MC2_v3_3Inst_1_U3  ( .A(\Red_MCInst_MC2_v3_1 [2]), .B(
        \MCInst_MC2_v3_2 [3]), .ZN(\MCInst_MC2_v3_3Inst_1_n2 ) );
  XOR2_X1 \MCInst_MC2_v0_0Inst_2_U3  ( .A(\Red_MCInst_MC2_v0_0 [0]), .B(
        \Red_MCInst_MC2_v0_1 [0]), .Z(\MCInst_MC2_v0_0 [2]) );
  XOR2_X1 \MCInst_MC2_v0_1Inst_2_U3  ( .A(\MCInst_MC2_v0_3 [3]), .B(
        \Red_MCInst_MC2_v0_1 [0]), .Z(\MCInst_MC2_v0_1 [2]) );
  XOR2_X1 \MCInst_MC2_v0_2Inst_2_U3  ( .A(\Red_MCInst_MC2_v0_2 [2]), .B(
        \Red_MCInst_MC2_v0_1 [0]), .Z(\MCInst_MC2_v0_2 [2]) );
  XNOR2_X1 \MCInst_MC2_v1_1Inst_2_U4  ( .A(\MCInst_MC2_v1_1Inst_2_n2 ), .B(
        \Red_MCInst_MC2_v1_2 [1]), .ZN(\MCInst_MC2_v1_1 [2]) );
  XNOR2_X1 \MCInst_MC2_v1_1Inst_2_U3  ( .A(\Red_MCInst_MC2_v1_1 [2]), .B(
        \MCInst_MC2_v1_0 [0]), .ZN(\MCInst_MC2_v1_1Inst_2_n2 ) );
  XNOR2_X1 \MCInst_MC2_v1_2Inst_2_U4  ( .A(\MCInst_MC2_v1_2Inst_2_n2 ), .B(
        \Red_MCInst_MC2_v1_2 [1]), .ZN(\MCInst_MC2_v1_2 [2]) );
  XNOR2_X1 \MCInst_MC2_v1_2Inst_2_U3  ( .A(\MCInst_MC2_v1_3 [3]), .B(
        \MCInst_MC2_v1_0 [0]), .ZN(\MCInst_MC2_v1_2Inst_2_n2 ) );
  XNOR2_X1 \MCInst_MC2_v2_1Inst_2_U4  ( .A(\MCInst_MC2_v2_1Inst_2_n2 ), .B(
        \MCInst_MC2_v2_0 [3]), .ZN(\MCInst_MC2_v2_1 [2]) );
  XNOR2_X1 \MCInst_MC2_v2_1Inst_2_U3  ( .A(\Red_MCInst_MC2_v2_2 [1]), .B(
        \Red_MCInst_MC2_v2_1 [1]), .ZN(\MCInst_MC2_v2_1Inst_2_n2 ) );
  XNOR2_X1 \MCInst_MC2_v2_2Inst_2_U4  ( .A(\MCInst_MC2_v2_2Inst_2_n2 ), .B(
        \MCInst_MC2_v2_0 [3]), .ZN(\MCInst_MC2_v2_2 [2]) );
  XNOR2_X1 \MCInst_MC2_v2_2Inst_2_U3  ( .A(\Red_MCInst_MC2_v2_2 [1]), .B(
        \MCInst_MC2_v2_0 [2]), .ZN(\MCInst_MC2_v2_2Inst_2_n2 ) );
  XOR2_X1 \MCInst_MC2_v2_3Inst_2_U3  ( .A(\Red_MCInst_MC2_v2_1 [1]), .B(
        \MCInst_MC2_v2_0 [2]), .Z(\MCInst_MC2_v2_3 [2]) );
  XNOR2_X1 \MCInst_MC2_v3_1Inst_2_U4  ( .A(\MCInst_MC2_v3_1Inst_2_n2 ), .B(
        \Red_MCInst_MC2_v3_3 [2]), .ZN(\MCInst_MC2_v3_1 [2]) );
  XNOR2_X1 \MCInst_MC2_v3_1Inst_2_U3  ( .A(\Red_MCInst_MC2_v3_1 [2]), .B(
        \MCInst_MC2_v3_2 [3]), .ZN(\MCInst_MC2_v3_1Inst_2_n2 ) );
  XOR2_X1 \MCInst_MC2_v3_3Inst_2_U3  ( .A(\Red_MCInst_MC2_v3_3 [2]), .B(
        \Red_MCInst_MC2_v3_1 [2]), .Z(\MCInst_MC2_v3_3 [2]) );
  XOR2_X1 \MCInst_MC2_v0_1Inst_3_U3  ( .A(\Red_MCInst_MC2_v0_0 [0]), .B(
        \Red_MCInst_MC2_v0_1 [0]), .Z(\MCInst_MC2_v0_1 [3]) );
  XOR2_X1 \MCInst_MC2_v0_2Inst_3_U3  ( .A(\Red_MCInst_MC2_v0_0 [0]), .B(
        \MCInst_MC2_v0_3 [3]), .Z(\MCInst_MC2_v0_2 [3]) );
  XOR2_X1 \MCInst_MC2_v1_1Inst_3_U3  ( .A(\Red_MCInst_MC2_v1_2 [1]), .B(
        \MCInst_MC2_v1_3 [3]), .Z(\MCInst_MC2_v1_1 [3]) );
  XNOR2_X1 \MCInst_MC2_v1_2Inst_3_U5  ( .A(\MCInst_MC2_v1_2Inst_3_n4 ), .B(
        \MCInst_MC2_v1_2Inst_3_n3 ), .ZN(\MCInst_MC2_v1_2 [3]) );
  XNOR2_X1 \MCInst_MC2_v1_2Inst_3_U4  ( .A(\Red_MCInst_MC2_v1_2 [1]), .B(
        \MCInst_MC2_v1_0 [0]), .ZN(\MCInst_MC2_v1_2Inst_3_n3 ) );
  XOR2_X1 \MCInst_MC2_v1_2Inst_3_U3  ( .A(\MCInst_MC2_v1_3 [3]), .B(
        \Red_MCInst_MC2_v1_1 [2]), .Z(\MCInst_MC2_v1_2Inst_3_n4 ) );
  XOR2_X1 \MCInst_MC2_v2_1Inst_3_U3  ( .A(\MCInst_MC2_v2_0 [2]), .B(
        \Red_MCInst_MC2_v2_2 [1]), .Z(\MCInst_MC2_v2_1 [3]) );
  XNOR2_X1 \MCInst_MC2_v2_2Inst_3_U4  ( .A(\MCInst_MC2_v2_2Inst_3_n2 ), .B(
        \MCInst_MC2_v2_0 [3]), .ZN(\MCInst_MC2_v2_2 [3]) );
  XNOR2_X1 \MCInst_MC2_v2_2Inst_3_U3  ( .A(\Red_MCInst_MC2_v2_2 [1]), .B(
        \Red_MCInst_MC2_v2_1 [1]), .ZN(\MCInst_MC2_v2_2Inst_3_n2 ) );
  XNOR2_X1 \MCInst_MC2_v2_3Inst_3_U4  ( .A(\MCInst_MC2_v2_3Inst_3_n2 ), .B(
        \MCInst_MC2_v2_0 [2]), .ZN(\MCInst_MC2_v2_3 [3]) );
  XNOR2_X1 \MCInst_MC2_v2_3Inst_3_U3  ( .A(\MCInst_MC2_v2_0 [3]), .B(
        \Red_MCInst_MC2_v2_1 [1]), .ZN(\MCInst_MC2_v2_3Inst_3_n2 ) );
  XOR2_X1 \MCInst_MC2_v3_1Inst_3_U3  ( .A(\Red_MCInst_MC2_v3_3 [2]), .B(
        \MCInst_MC2_v3_0 [3]), .Z(\MCInst_MC2_v3_1 [3]) );
  XOR2_X1 \MCInst_MC2_v3_3Inst_3_U3  ( .A(\MCInst_MC2_v3_2 [3]), .B(
        \MCInst_MC2_v3_0 [3]), .Z(\MCInst_MC2_v3_3 [3]) );
  XNOR2_X1 \MCInst_MC2_r0Inst_XORInst_0_0_U3  ( .A(
        \MCInst_MC2_r0Inst_XORInst_0_0_n5 ), .B(
        \MCInst_MC2_r0Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[52]) );
  XNOR2_X1 \MCInst_MC2_r0Inst_XORInst_0_0_U2  ( .A(\Red_MCInst_MC2_v3_1 [2]), 
        .B(\Red_MCInst_MC2_v2_2 [1]), .ZN(\MCInst_MC2_r0Inst_XORInst_0_0_n4 )
         );
  XOR2_X1 \MCInst_MC2_r0Inst_XORInst_0_0_U1  ( .A(\MCInst_MC2_v0_3 [3]), .B(
        \MCInst_MC2_v1_0 [0]), .Z(\MCInst_MC2_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \MCInst_MC2_r0Inst_XORInst_0_1_U3  ( .A(
        \MCInst_MC2_r0Inst_XORInst_0_1_n5 ), .B(
        \MCInst_MC2_r0Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[53]) );
  XNOR2_X1 \MCInst_MC2_r0Inst_XORInst_0_1_U2  ( .A(\MCInst_MC2_v3_0 [1]), .B(
        \MCInst_MC2_v2_0 [1]), .ZN(\MCInst_MC2_r0Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \MCInst_MC2_r0Inst_XORInst_0_1_U1  ( .A(\MCInst_MC2_v0_0 [1]), .B(
        \Red_MCInst_MC2_v1_2 [1]), .Z(\MCInst_MC2_r0Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \MCInst_MC2_r0Inst_XORInst_0_2_U3  ( .A(
        \MCInst_MC2_r0Inst_XORInst_0_2_n5 ), .B(
        \MCInst_MC2_r0Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[54]) );
  XNOR2_X1 \MCInst_MC2_r0Inst_XORInst_0_2_U2  ( .A(\Red_MCInst_MC2_v3_3 [2]), 
        .B(\MCInst_MC2_v2_0 [2]), .ZN(\MCInst_MC2_r0Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \MCInst_MC2_r0Inst_XORInst_0_2_U1  ( .A(\MCInst_MC2_v0_0 [2]), .B(
        \MCInst_MC2_v1_3 [3]), .Z(\MCInst_MC2_r0Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \MCInst_MC2_r0Inst_XORInst_0_3_U3  ( .A(
        \MCInst_MC2_r0Inst_XORInst_0_3_n5 ), .B(
        \MCInst_MC2_r0Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[55]) );
  XNOR2_X1 \MCInst_MC2_r0Inst_XORInst_0_3_U2  ( .A(\MCInst_MC2_v3_0 [3]), .B(
        \MCInst_MC2_v2_0 [3]), .ZN(\MCInst_MC2_r0Inst_XORInst_0_3_n4 ) );
  XOR2_X1 \MCInst_MC2_r0Inst_XORInst_0_3_U1  ( .A(\Red_MCInst_MC2_v0_2 [2]), 
        .B(\Red_MCInst_MC2_v1_1 [2]), .Z(\MCInst_MC2_r0Inst_XORInst_0_3_n5 )
         );
  XNOR2_X1 \MCInst_MC2_r1Inst_XORInst_0_0_U3  ( .A(
        \MCInst_MC2_r1Inst_XORInst_0_0_n5 ), .B(
        \MCInst_MC2_r1Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[36]) );
  XNOR2_X1 \MCInst_MC2_r1Inst_XORInst_0_0_U2  ( .A(\MCInst_MC2_v3_1 [0]), .B(
        \MCInst_MC2_v2_1 [0]), .ZN(\MCInst_MC2_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \MCInst_MC2_r1Inst_XORInst_0_0_U1  ( .A(\Red_MCInst_MC2_v0_2 [2]), 
        .B(\MCInst_MC2_v1_1 [0]), .Z(\MCInst_MC2_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \MCInst_MC2_r1Inst_XORInst_0_1_U3  ( .A(
        \MCInst_MC2_r1Inst_XORInst_0_1_n5 ), .B(
        \MCInst_MC2_r1Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[37]) );
  XNOR2_X1 \MCInst_MC2_r1Inst_XORInst_0_1_U2  ( .A(\MCInst_MC2_v3_1 [1]), .B(
        \MCInst_MC2_v2_1 [1]), .ZN(\MCInst_MC2_r1Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \MCInst_MC2_r1Inst_XORInst_0_1_U1  ( .A(\MCInst_MC2_v0_1 [1]), .B(
        \MCInst_MC2_v1_1 [1]), .Z(\MCInst_MC2_r1Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \MCInst_MC2_r1Inst_XORInst_0_2_U3  ( .A(
        \MCInst_MC2_r1Inst_XORInst_0_2_n5 ), .B(
        \MCInst_MC2_r1Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[38]) );
  XNOR2_X1 \MCInst_MC2_r1Inst_XORInst_0_2_U2  ( .A(\MCInst_MC2_v3_1 [2]), .B(
        \MCInst_MC2_v2_1 [2]), .ZN(\MCInst_MC2_r1Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \MCInst_MC2_r1Inst_XORInst_0_2_U1  ( .A(\MCInst_MC2_v0_1 [2]), .B(
        \MCInst_MC2_v1_1 [2]), .Z(\MCInst_MC2_r1Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \MCInst_MC2_r1Inst_XORInst_0_3_U3  ( .A(
        \MCInst_MC2_r1Inst_XORInst_0_3_n5 ), .B(
        \MCInst_MC2_r1Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[39]) );
  XNOR2_X1 \MCInst_MC2_r1Inst_XORInst_0_3_U2  ( .A(\MCInst_MC2_v3_1 [3]), .B(
        \MCInst_MC2_v2_1 [3]), .ZN(\MCInst_MC2_r1Inst_XORInst_0_3_n4 ) );
  XOR2_X1 \MCInst_MC2_r1Inst_XORInst_0_3_U1  ( .A(\MCInst_MC2_v0_1 [3]), .B(
        \MCInst_MC2_v1_1 [3]), .Z(\MCInst_MC2_r1Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 \MCInst_MC2_r2Inst_XORInst_0_0_U3  ( .A(
        \MCInst_MC2_r2Inst_XORInst_0_0_n5 ), .B(
        \MCInst_MC2_r2Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[20]) );
  XNOR2_X1 \MCInst_MC2_r2Inst_XORInst_0_0_U2  ( .A(\MCInst_MC2_v3_2 [0]), .B(
        \MCInst_MC2_v2_2 [0]), .ZN(\MCInst_MC2_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \MCInst_MC2_r2Inst_XORInst_0_0_U1  ( .A(\MCInst_MC2_v0_2 [0]), .B(
        \MCInst_MC2_v1_2 [0]), .Z(\MCInst_MC2_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \MCInst_MC2_r2Inst_XORInst_0_1_U3  ( .A(
        \MCInst_MC2_r2Inst_XORInst_0_1_n5 ), .B(
        \MCInst_MC2_r2Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[21]) );
  XNOR2_X1 \MCInst_MC2_r2Inst_XORInst_0_1_U2  ( .A(\MCInst_MC2_v3_0 [3]), .B(
        \MCInst_MC2_v2_2 [1]), .ZN(\MCInst_MC2_r2Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \MCInst_MC2_r2Inst_XORInst_0_1_U1  ( .A(\MCInst_MC2_v0_2 [1]), .B(
        \MCInst_MC2_v1_2 [1]), .Z(\MCInst_MC2_r2Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \MCInst_MC2_r2Inst_XORInst_0_2_U3  ( .A(
        \MCInst_MC2_r2Inst_XORInst_0_2_n5 ), .B(
        \MCInst_MC2_r2Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[22]) );
  XNOR2_X1 \MCInst_MC2_r2Inst_XORInst_0_2_U2  ( .A(\Red_MCInst_MC2_v3_1 [2]), 
        .B(\MCInst_MC2_v2_2 [2]), .ZN(\MCInst_MC2_r2Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \MCInst_MC2_r2Inst_XORInst_0_2_U1  ( .A(\MCInst_MC2_v0_2 [2]), .B(
        \MCInst_MC2_v1_2 [2]), .Z(\MCInst_MC2_r2Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \MCInst_MC2_r2Inst_XORInst_0_3_U3  ( .A(
        \MCInst_MC2_r2Inst_XORInst_0_3_n5 ), .B(
        \MCInst_MC2_r2Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[23]) );
  XNOR2_X1 \MCInst_MC2_r2Inst_XORInst_0_3_U2  ( .A(\MCInst_MC2_v3_2 [3]), .B(
        \MCInst_MC2_v2_2 [3]), .ZN(\MCInst_MC2_r2Inst_XORInst_0_3_n4 ) );
  XOR2_X1 \MCInst_MC2_r2Inst_XORInst_0_3_U1  ( .A(\MCInst_MC2_v0_2 [3]), .B(
        \MCInst_MC2_v1_2 [3]), .Z(\MCInst_MC2_r2Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 \MCInst_MC2_r3Inst_XORInst_0_0_U3  ( .A(
        \MCInst_MC2_r3Inst_XORInst_0_0_n5 ), .B(
        \MCInst_MC2_r3Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[4]) );
  XNOR2_X1 \MCInst_MC2_r3Inst_XORInst_0_0_U2  ( .A(\MCInst_MC2_v3_3 [0]), .B(
        \MCInst_MC2_v2_3 [0]), .ZN(\MCInst_MC2_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \MCInst_MC2_r3Inst_XORInst_0_0_U1  ( .A(\Red_MCInst_MC2_v0_1 [0]), 
        .B(\Red_MCInst_MC2_v1_1 [2]), .Z(\MCInst_MC2_r3Inst_XORInst_0_0_n5 )
         );
  XNOR2_X1 \MCInst_MC2_r3Inst_XORInst_0_1_U3  ( .A(
        \MCInst_MC2_r3Inst_XORInst_0_1_n5 ), .B(
        \MCInst_MC2_r3Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[5]) );
  XNOR2_X1 \MCInst_MC2_r3Inst_XORInst_0_1_U2  ( .A(\MCInst_MC2_v3_3 [1]), .B(
        \Red_MCInst_MC2_v2_1 [1]), .ZN(\MCInst_MC2_r3Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \MCInst_MC2_r3Inst_XORInst_0_1_U1  ( .A(\MCInst_MC2_v0_3 [1]), .B(
        \MCInst_MC2_v1_3 [1]), .Z(\MCInst_MC2_r3Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \MCInst_MC2_r3Inst_XORInst_0_2_U3  ( .A(
        \MCInst_MC2_r3Inst_XORInst_0_2_n5 ), .B(
        \MCInst_MC2_r3Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[6]) );
  XNOR2_X1 \MCInst_MC2_r3Inst_XORInst_0_2_U2  ( .A(\MCInst_MC2_v3_3 [2]), .B(
        \MCInst_MC2_v2_3 [2]), .ZN(\MCInst_MC2_r3Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \MCInst_MC2_r3Inst_XORInst_0_2_U1  ( .A(\Red_MCInst_MC2_v0_2 [2]), 
        .B(\Red_MCInst_MC2_v1_2 [1]), .Z(\MCInst_MC2_r3Inst_XORInst_0_2_n5 )
         );
  XNOR2_X1 \MCInst_MC2_r3Inst_XORInst_0_3_U3  ( .A(
        \MCInst_MC2_r3Inst_XORInst_0_3_n5 ), .B(
        \MCInst_MC2_r3Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[7]) );
  XNOR2_X1 \MCInst_MC2_r3Inst_XORInst_0_3_U2  ( .A(\MCInst_MC2_v3_3 [3]), .B(
        \MCInst_MC2_v2_3 [3]), .ZN(\MCInst_MC2_r3Inst_XORInst_0_3_n4 ) );
  XOR2_X1 \MCInst_MC2_r3Inst_XORInst_0_3_U1  ( .A(\MCInst_MC2_v0_3 [3]), .B(
        \MCInst_MC2_v1_3 [3]), .Z(\MCInst_MC2_r3Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 \MCInst_MC3_v0_2Inst_0_U4  ( .A(\MCInst_MC3_v0_2Inst_0_n2 ), .B(
        \Red_MCInst_MC3_v0_2 [2]), .ZN(\MCInst_MC3_v0_2 [0]) );
  XNOR2_X1 \MCInst_MC3_v0_2Inst_0_U3  ( .A(\Red_MCInst_MC3_v0_1 [0]), .B(
        \Red_MCInst_MC3_v0_0 [0]), .ZN(\MCInst_MC3_v0_2Inst_0_n2 ) );
  XOR2_X1 \MCInst_MC3_v1_1Inst_0_U3  ( .A(\MCInst_MC3_v1_3 [3]), .B(
        \Red_MCInst_MC3_v1_1 [2]), .Z(\MCInst_MC3_v1_1 [0]) );
  XNOR2_X1 \MCInst_MC3_v1_2Inst_0_U4  ( .A(\MCInst_MC3_v1_2Inst_0_n2 ), .B(
        \MCInst_MC3_v1_3 [3]), .ZN(\MCInst_MC3_v1_2 [0]) );
  XNOR2_X1 \MCInst_MC3_v1_2Inst_0_U3  ( .A(\Red_MCInst_MC3_v1_1 [2]), .B(
        \Red_MCInst_MC3_v1_2 [1]), .ZN(\MCInst_MC3_v1_2Inst_0_n2 ) );
  XOR2_X1 \MCInst_MC3_v2_1Inst_0_U3  ( .A(\Red_MCInst_MC3_v2_1 [1]), .B(
        \MCInst_MC3_v2_0 [3]), .Z(\MCInst_MC3_v2_1 [0]) );
  XOR2_X1 \MCInst_MC3_v2_2Inst_0_U3  ( .A(\MCInst_MC3_v2_0 [2]), .B(
        \Red_MCInst_MC3_v2_2 [1]), .Z(\MCInst_MC3_v2_2 [0]) );
  XNOR2_X1 \MCInst_MC3_v2_3Inst_0_U5  ( .A(\MCInst_MC3_v2_3Inst_0_n4 ), .B(
        \MCInst_MC3_v2_3Inst_0_n3 ), .ZN(\MCInst_MC3_v2_3 [0]) );
  XNOR2_X1 \MCInst_MC3_v2_3Inst_0_U4  ( .A(\MCInst_MC3_v2_0 [2]), .B(
        \Red_MCInst_MC3_v2_1 [1]), .ZN(\MCInst_MC3_v2_3Inst_0_n3 ) );
  XOR2_X1 \MCInst_MC3_v2_3Inst_0_U3  ( .A(\MCInst_MC3_v2_0 [3]), .B(
        \Red_MCInst_MC3_v2_2 [1]), .Z(\MCInst_MC3_v2_3Inst_0_n4 ) );
  XOR2_X1 \MCInst_MC3_v3_1Inst_0_U3  ( .A(\MCInst_MC3_v3_0 [3]), .B(
        \Red_MCInst_MC3_v3_1 [2]), .Z(\MCInst_MC3_v3_1 [0]) );
  XOR2_X1 \MCInst_MC3_v3_2Inst_0_U3  ( .A(\MCInst_MC3_v3_2 [3]), .B(
        \Red_MCInst_MC3_v3_3 [2]), .Z(\MCInst_MC3_v3_2 [0]) );
  XNOR2_X1 \MCInst_MC3_v3_3Inst_0_U4  ( .A(\MCInst_MC3_v3_3Inst_0_n2 ), .B(
        \Red_MCInst_MC3_v3_3 [2]), .ZN(\MCInst_MC3_v3_3 [0]) );
  XNOR2_X1 \MCInst_MC3_v3_3Inst_0_U3  ( .A(\Red_MCInst_MC3_v3_1 [2]), .B(
        \MCInst_MC3_v3_2 [3]), .ZN(\MCInst_MC3_v3_3Inst_0_n2 ) );
  XOR2_X1 \MCInst_MC3_v0_0Inst_1_U3  ( .A(\MCInst_MC3_v0_3 [3]), .B(
        \Red_MCInst_MC3_v0_1 [0]), .Z(\MCInst_MC3_v0_0 [1]) );
  XOR2_X1 \MCInst_MC3_v0_1Inst_1_U3  ( .A(\Red_MCInst_MC3_v0_2 [2]), .B(
        \MCInst_MC3_v0_3 [3]), .Z(\MCInst_MC3_v0_1 [1]) );
  XNOR2_X1 \MCInst_MC3_v0_2Inst_1_U4  ( .A(\MCInst_MC3_v0_2Inst_1_n2 ), .B(
        \MCInst_MC3_v0_3 [3]), .ZN(\MCInst_MC3_v0_2 [1]) );
  XNOR2_X1 \MCInst_MC3_v0_2Inst_1_U3  ( .A(\Red_MCInst_MC3_v0_1 [0]), .B(
        \Red_MCInst_MC3_v0_0 [0]), .ZN(\MCInst_MC3_v0_2Inst_1_n2 ) );
  XOR2_X1 \MCInst_MC3_v0_3Inst_1_U3  ( .A(\Red_MCInst_MC3_v0_0 [0]), .B(
        \Red_MCInst_MC3_v0_1 [0]), .Z(\MCInst_MC3_v0_3 [1]) );
  XOR2_X1 \MCInst_MC3_v1_1Inst_1_U3  ( .A(\MCInst_MC3_v1_0 [0]), .B(
        \MCInst_MC3_v1_3 [3]), .Z(\MCInst_MC3_v1_1 [1]) );
  XOR2_X1 \MCInst_MC3_v1_2Inst_1_U3  ( .A(\MCInst_MC3_v1_0 [0]), .B(
        \Red_MCInst_MC3_v1_2 [1]), .Z(\MCInst_MC3_v1_2 [1]) );
  XOR2_X1 \MCInst_MC3_v1_3Inst_1_U3  ( .A(\MCInst_MC3_v1_0 [0]), .B(
        \Red_MCInst_MC3_v1_1 [2]), .Z(\MCInst_MC3_v1_3 [1]) );
  XOR2_X1 \MCInst_MC3_v2_0Inst_1_U3  ( .A(\Red_MCInst_MC3_v2_1 [1]), .B(
        \Red_MCInst_MC3_v2_2 [1]), .Z(\MCInst_MC3_v2_0 [1]) );
  XNOR2_X1 \MCInst_MC3_v2_1Inst_1_U4  ( .A(\MCInst_MC3_v2_1Inst_1_n2 ), .B(
        \MCInst_MC3_v2_0 [3]), .ZN(\MCInst_MC3_v2_1 [1]) );
  XNOR2_X1 \MCInst_MC3_v2_1Inst_1_U3  ( .A(\Red_MCInst_MC3_v2_2 [1]), .B(
        \MCInst_MC3_v2_0 [2]), .ZN(\MCInst_MC3_v2_1Inst_1_n2 ) );
  XNOR2_X1 \MCInst_MC3_v2_2Inst_1_U5  ( .A(\MCInst_MC3_v2_2Inst_1_n4 ), .B(
        \MCInst_MC3_v2_2Inst_1_n3 ), .ZN(\MCInst_MC3_v2_2 [1]) );
  XNOR2_X1 \MCInst_MC3_v2_2Inst_1_U4  ( .A(\MCInst_MC3_v2_0 [2]), .B(
        \Red_MCInst_MC3_v2_1 [1]), .ZN(\MCInst_MC3_v2_2Inst_1_n3 ) );
  XOR2_X1 \MCInst_MC3_v2_2Inst_1_U3  ( .A(\MCInst_MC3_v2_0 [3]), .B(
        \Red_MCInst_MC3_v2_2 [1]), .Z(\MCInst_MC3_v2_2Inst_1_n4 ) );
  XOR2_X1 \MCInst_MC3_v3_0Inst_1_U3  ( .A(\MCInst_MC3_v3_2 [3]), .B(
        \Red_MCInst_MC3_v3_1 [2]), .Z(\MCInst_MC3_v3_0 [1]) );
  XOR2_X1 \MCInst_MC3_v3_1Inst_1_U3  ( .A(\MCInst_MC3_v3_2 [3]), .B(
        \MCInst_MC3_v3_0 [3]), .Z(\MCInst_MC3_v3_1 [1]) );
  XNOR2_X1 \MCInst_MC3_v3_3Inst_1_U4  ( .A(\MCInst_MC3_v3_3Inst_1_n2 ), .B(
        \MCInst_MC3_v3_0 [3]), .ZN(\MCInst_MC3_v3_3 [1]) );
  XNOR2_X1 \MCInst_MC3_v3_3Inst_1_U3  ( .A(\Red_MCInst_MC3_v3_1 [2]), .B(
        \MCInst_MC3_v3_2 [3]), .ZN(\MCInst_MC3_v3_3Inst_1_n2 ) );
  XOR2_X1 \MCInst_MC3_v0_0Inst_2_U3  ( .A(\Red_MCInst_MC3_v0_0 [0]), .B(
        \Red_MCInst_MC3_v0_1 [0]), .Z(\MCInst_MC3_v0_0 [2]) );
  XOR2_X1 \MCInst_MC3_v0_1Inst_2_U3  ( .A(\MCInst_MC3_v0_3 [3]), .B(
        \Red_MCInst_MC3_v0_1 [0]), .Z(\MCInst_MC3_v0_1 [2]) );
  XOR2_X1 \MCInst_MC3_v0_2Inst_2_U3  ( .A(\Red_MCInst_MC3_v0_2 [2]), .B(
        \Red_MCInst_MC3_v0_1 [0]), .Z(\MCInst_MC3_v0_2 [2]) );
  XNOR2_X1 \MCInst_MC3_v1_1Inst_2_U4  ( .A(\MCInst_MC3_v1_1Inst_2_n2 ), .B(
        \Red_MCInst_MC3_v1_2 [1]), .ZN(\MCInst_MC3_v1_1 [2]) );
  XNOR2_X1 \MCInst_MC3_v1_1Inst_2_U3  ( .A(\Red_MCInst_MC3_v1_1 [2]), .B(
        \MCInst_MC3_v1_0 [0]), .ZN(\MCInst_MC3_v1_1Inst_2_n2 ) );
  XNOR2_X1 \MCInst_MC3_v1_2Inst_2_U4  ( .A(\MCInst_MC3_v1_2Inst_2_n2 ), .B(
        \Red_MCInst_MC3_v1_2 [1]), .ZN(\MCInst_MC3_v1_2 [2]) );
  XNOR2_X1 \MCInst_MC3_v1_2Inst_2_U3  ( .A(\MCInst_MC3_v1_3 [3]), .B(
        \MCInst_MC3_v1_0 [0]), .ZN(\MCInst_MC3_v1_2Inst_2_n2 ) );
  XNOR2_X1 \MCInst_MC3_v2_1Inst_2_U4  ( .A(\MCInst_MC3_v2_1Inst_2_n2 ), .B(
        \MCInst_MC3_v2_0 [3]), .ZN(\MCInst_MC3_v2_1 [2]) );
  XNOR2_X1 \MCInst_MC3_v2_1Inst_2_U3  ( .A(\Red_MCInst_MC3_v2_2 [1]), .B(
        \Red_MCInst_MC3_v2_1 [1]), .ZN(\MCInst_MC3_v2_1Inst_2_n2 ) );
  XNOR2_X1 \MCInst_MC3_v2_2Inst_2_U4  ( .A(\MCInst_MC3_v2_2Inst_2_n2 ), .B(
        \MCInst_MC3_v2_0 [3]), .ZN(\MCInst_MC3_v2_2 [2]) );
  XNOR2_X1 \MCInst_MC3_v2_2Inst_2_U3  ( .A(\Red_MCInst_MC3_v2_2 [1]), .B(
        \MCInst_MC3_v2_0 [2]), .ZN(\MCInst_MC3_v2_2Inst_2_n2 ) );
  XOR2_X1 \MCInst_MC3_v2_3Inst_2_U3  ( .A(\Red_MCInst_MC3_v2_1 [1]), .B(
        \MCInst_MC3_v2_0 [2]), .Z(\MCInst_MC3_v2_3 [2]) );
  XNOR2_X1 \MCInst_MC3_v3_1Inst_2_U4  ( .A(\MCInst_MC3_v3_1Inst_2_n2 ), .B(
        \Red_MCInst_MC3_v3_3 [2]), .ZN(\MCInst_MC3_v3_1 [2]) );
  XNOR2_X1 \MCInst_MC3_v3_1Inst_2_U3  ( .A(\Red_MCInst_MC3_v3_1 [2]), .B(
        \MCInst_MC3_v3_2 [3]), .ZN(\MCInst_MC3_v3_1Inst_2_n2 ) );
  XOR2_X1 \MCInst_MC3_v3_3Inst_2_U3  ( .A(\Red_MCInst_MC3_v3_3 [2]), .B(
        \Red_MCInst_MC3_v3_1 [2]), .Z(\MCInst_MC3_v3_3 [2]) );
  XOR2_X1 \MCInst_MC3_v0_1Inst_3_U3  ( .A(\Red_MCInst_MC3_v0_0 [0]), .B(
        \Red_MCInst_MC3_v0_1 [0]), .Z(\MCInst_MC3_v0_1 [3]) );
  XOR2_X1 \MCInst_MC3_v0_2Inst_3_U3  ( .A(\Red_MCInst_MC3_v0_0 [0]), .B(
        \MCInst_MC3_v0_3 [3]), .Z(\MCInst_MC3_v0_2 [3]) );
  XOR2_X1 \MCInst_MC3_v1_1Inst_3_U3  ( .A(\Red_MCInst_MC3_v1_2 [1]), .B(
        \MCInst_MC3_v1_3 [3]), .Z(\MCInst_MC3_v1_1 [3]) );
  XNOR2_X1 \MCInst_MC3_v1_2Inst_3_U5  ( .A(\MCInst_MC3_v1_2Inst_3_n4 ), .B(
        \MCInst_MC3_v1_2Inst_3_n3 ), .ZN(\MCInst_MC3_v1_2 [3]) );
  XNOR2_X1 \MCInst_MC3_v1_2Inst_3_U4  ( .A(\Red_MCInst_MC3_v1_2 [1]), .B(
        \MCInst_MC3_v1_0 [0]), .ZN(\MCInst_MC3_v1_2Inst_3_n3 ) );
  XOR2_X1 \MCInst_MC3_v1_2Inst_3_U3  ( .A(\MCInst_MC3_v1_3 [3]), .B(
        \Red_MCInst_MC3_v1_1 [2]), .Z(\MCInst_MC3_v1_2Inst_3_n4 ) );
  XOR2_X1 \MCInst_MC3_v2_1Inst_3_U3  ( .A(\MCInst_MC3_v2_0 [2]), .B(
        \Red_MCInst_MC3_v2_2 [1]), .Z(\MCInst_MC3_v2_1 [3]) );
  XNOR2_X1 \MCInst_MC3_v2_2Inst_3_U4  ( .A(\MCInst_MC3_v2_2Inst_3_n2 ), .B(
        \MCInst_MC3_v2_0 [3]), .ZN(\MCInst_MC3_v2_2 [3]) );
  XNOR2_X1 \MCInst_MC3_v2_2Inst_3_U3  ( .A(\Red_MCInst_MC3_v2_2 [1]), .B(
        \Red_MCInst_MC3_v2_1 [1]), .ZN(\MCInst_MC3_v2_2Inst_3_n2 ) );
  XNOR2_X1 \MCInst_MC3_v2_3Inst_3_U4  ( .A(\MCInst_MC3_v2_3Inst_3_n2 ), .B(
        \MCInst_MC3_v2_0 [2]), .ZN(\MCInst_MC3_v2_3 [3]) );
  XNOR2_X1 \MCInst_MC3_v2_3Inst_3_U3  ( .A(\MCInst_MC3_v2_0 [3]), .B(
        \Red_MCInst_MC3_v2_1 [1]), .ZN(\MCInst_MC3_v2_3Inst_3_n2 ) );
  XOR2_X1 \MCInst_MC3_v3_1Inst_3_U3  ( .A(\Red_MCInst_MC3_v3_3 [2]), .B(
        \MCInst_MC3_v3_0 [3]), .Z(\MCInst_MC3_v3_1 [3]) );
  XOR2_X1 \MCInst_MC3_v3_3Inst_3_U3  ( .A(\MCInst_MC3_v3_2 [3]), .B(
        \MCInst_MC3_v3_0 [3]), .Z(\MCInst_MC3_v3_3 [3]) );
  XNOR2_X1 \MCInst_MC3_r0Inst_XORInst_0_0_U3  ( .A(
        \MCInst_MC3_r0Inst_XORInst_0_0_n5 ), .B(
        \MCInst_MC3_r0Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[48]) );
  XNOR2_X1 \MCInst_MC3_r0Inst_XORInst_0_0_U2  ( .A(\Red_MCInst_MC3_v3_1 [2]), 
        .B(\Red_MCInst_MC3_v2_2 [1]), .ZN(\MCInst_MC3_r0Inst_XORInst_0_0_n4 )
         );
  XOR2_X1 \MCInst_MC3_r0Inst_XORInst_0_0_U1  ( .A(\MCInst_MC3_v0_3 [3]), .B(
        \MCInst_MC3_v1_0 [0]), .Z(\MCInst_MC3_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \MCInst_MC3_r0Inst_XORInst_0_1_U3  ( .A(
        \MCInst_MC3_r0Inst_XORInst_0_1_n5 ), .B(
        \MCInst_MC3_r0Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[49]) );
  XNOR2_X1 \MCInst_MC3_r0Inst_XORInst_0_1_U2  ( .A(\MCInst_MC3_v3_0 [1]), .B(
        \MCInst_MC3_v2_0 [1]), .ZN(\MCInst_MC3_r0Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \MCInst_MC3_r0Inst_XORInst_0_1_U1  ( .A(\MCInst_MC3_v0_0 [1]), .B(
        \Red_MCInst_MC3_v1_2 [1]), .Z(\MCInst_MC3_r0Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \MCInst_MC3_r0Inst_XORInst_0_2_U3  ( .A(
        \MCInst_MC3_r0Inst_XORInst_0_2_n5 ), .B(
        \MCInst_MC3_r0Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[50]) );
  XNOR2_X1 \MCInst_MC3_r0Inst_XORInst_0_2_U2  ( .A(\Red_MCInst_MC3_v3_3 [2]), 
        .B(\MCInst_MC3_v2_0 [2]), .ZN(\MCInst_MC3_r0Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \MCInst_MC3_r0Inst_XORInst_0_2_U1  ( .A(\MCInst_MC3_v0_0 [2]), .B(
        \MCInst_MC3_v1_3 [3]), .Z(\MCInst_MC3_r0Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \MCInst_MC3_r0Inst_XORInst_0_3_U3  ( .A(
        \MCInst_MC3_r0Inst_XORInst_0_3_n5 ), .B(
        \MCInst_MC3_r0Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[51]) );
  XNOR2_X1 \MCInst_MC3_r0Inst_XORInst_0_3_U2  ( .A(\MCInst_MC3_v3_0 [3]), .B(
        \MCInst_MC3_v2_0 [3]), .ZN(\MCInst_MC3_r0Inst_XORInst_0_3_n4 ) );
  XOR2_X1 \MCInst_MC3_r0Inst_XORInst_0_3_U1  ( .A(\Red_MCInst_MC3_v0_2 [2]), 
        .B(\Red_MCInst_MC3_v1_1 [2]), .Z(\MCInst_MC3_r0Inst_XORInst_0_3_n5 )
         );
  XNOR2_X1 \MCInst_MC3_r1Inst_XORInst_0_0_U3  ( .A(
        \MCInst_MC3_r1Inst_XORInst_0_0_n5 ), .B(
        \MCInst_MC3_r1Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[32]) );
  XNOR2_X1 \MCInst_MC3_r1Inst_XORInst_0_0_U2  ( .A(\MCInst_MC3_v3_1 [0]), .B(
        \MCInst_MC3_v2_1 [0]), .ZN(\MCInst_MC3_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \MCInst_MC3_r1Inst_XORInst_0_0_U1  ( .A(\Red_MCInst_MC3_v0_2 [2]), 
        .B(\MCInst_MC3_v1_1 [0]), .Z(\MCInst_MC3_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \MCInst_MC3_r1Inst_XORInst_0_1_U3  ( .A(
        \MCInst_MC3_r1Inst_XORInst_0_1_n5 ), .B(
        \MCInst_MC3_r1Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[33]) );
  XNOR2_X1 \MCInst_MC3_r1Inst_XORInst_0_1_U2  ( .A(\MCInst_MC3_v3_1 [1]), .B(
        \MCInst_MC3_v2_1 [1]), .ZN(\MCInst_MC3_r1Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \MCInst_MC3_r1Inst_XORInst_0_1_U1  ( .A(\MCInst_MC3_v0_1 [1]), .B(
        \MCInst_MC3_v1_1 [1]), .Z(\MCInst_MC3_r1Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \MCInst_MC3_r1Inst_XORInst_0_2_U3  ( .A(
        \MCInst_MC3_r1Inst_XORInst_0_2_n5 ), .B(
        \MCInst_MC3_r1Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[34]) );
  XNOR2_X1 \MCInst_MC3_r1Inst_XORInst_0_2_U2  ( .A(\MCInst_MC3_v3_1 [2]), .B(
        \MCInst_MC3_v2_1 [2]), .ZN(\MCInst_MC3_r1Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \MCInst_MC3_r1Inst_XORInst_0_2_U1  ( .A(\MCInst_MC3_v0_1 [2]), .B(
        \MCInst_MC3_v1_1 [2]), .Z(\MCInst_MC3_r1Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \MCInst_MC3_r1Inst_XORInst_0_3_U3  ( .A(
        \MCInst_MC3_r1Inst_XORInst_0_3_n5 ), .B(
        \MCInst_MC3_r1Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[35]) );
  XNOR2_X1 \MCInst_MC3_r1Inst_XORInst_0_3_U2  ( .A(\MCInst_MC3_v3_1 [3]), .B(
        \MCInst_MC3_v2_1 [3]), .ZN(\MCInst_MC3_r1Inst_XORInst_0_3_n4 ) );
  XOR2_X1 \MCInst_MC3_r1Inst_XORInst_0_3_U1  ( .A(\MCInst_MC3_v0_1 [3]), .B(
        \MCInst_MC3_v1_1 [3]), .Z(\MCInst_MC3_r1Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 \MCInst_MC3_r2Inst_XORInst_0_0_U3  ( .A(
        \MCInst_MC3_r2Inst_XORInst_0_0_n5 ), .B(
        \MCInst_MC3_r2Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[16]) );
  XNOR2_X1 \MCInst_MC3_r2Inst_XORInst_0_0_U2  ( .A(\MCInst_MC3_v3_2 [0]), .B(
        \MCInst_MC3_v2_2 [0]), .ZN(\MCInst_MC3_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \MCInst_MC3_r2Inst_XORInst_0_0_U1  ( .A(\MCInst_MC3_v0_2 [0]), .B(
        \MCInst_MC3_v1_2 [0]), .Z(\MCInst_MC3_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \MCInst_MC3_r2Inst_XORInst_0_1_U3  ( .A(
        \MCInst_MC3_r2Inst_XORInst_0_1_n5 ), .B(
        \MCInst_MC3_r2Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[17]) );
  XNOR2_X1 \MCInst_MC3_r2Inst_XORInst_0_1_U2  ( .A(\MCInst_MC3_v3_0 [3]), .B(
        \MCInst_MC3_v2_2 [1]), .ZN(\MCInst_MC3_r2Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \MCInst_MC3_r2Inst_XORInst_0_1_U1  ( .A(\MCInst_MC3_v0_2 [1]), .B(
        \MCInst_MC3_v1_2 [1]), .Z(\MCInst_MC3_r2Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \MCInst_MC3_r2Inst_XORInst_0_2_U3  ( .A(
        \MCInst_MC3_r2Inst_XORInst_0_2_n5 ), .B(
        \MCInst_MC3_r2Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[18]) );
  XNOR2_X1 \MCInst_MC3_r2Inst_XORInst_0_2_U2  ( .A(\Red_MCInst_MC3_v3_1 [2]), 
        .B(\MCInst_MC3_v2_2 [2]), .ZN(\MCInst_MC3_r2Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \MCInst_MC3_r2Inst_XORInst_0_2_U1  ( .A(\MCInst_MC3_v0_2 [2]), .B(
        \MCInst_MC3_v1_2 [2]), .Z(\MCInst_MC3_r2Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \MCInst_MC3_r2Inst_XORInst_0_3_U3  ( .A(
        \MCInst_MC3_r2Inst_XORInst_0_3_n5 ), .B(
        \MCInst_MC3_r2Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[19]) );
  XNOR2_X1 \MCInst_MC3_r2Inst_XORInst_0_3_U2  ( .A(\MCInst_MC3_v3_2 [3]), .B(
        \MCInst_MC3_v2_2 [3]), .ZN(\MCInst_MC3_r2Inst_XORInst_0_3_n4 ) );
  XOR2_X1 \MCInst_MC3_r2Inst_XORInst_0_3_U1  ( .A(\MCInst_MC3_v0_2 [3]), .B(
        \MCInst_MC3_v1_2 [3]), .Z(\MCInst_MC3_r2Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 \MCInst_MC3_r3Inst_XORInst_0_0_U3  ( .A(
        \MCInst_MC3_r3Inst_XORInst_0_0_n5 ), .B(
        \MCInst_MC3_r3Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[0]) );
  XNOR2_X1 \MCInst_MC3_r3Inst_XORInst_0_0_U2  ( .A(\MCInst_MC3_v3_3 [0]), .B(
        \MCInst_MC3_v2_3 [0]), .ZN(\MCInst_MC3_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \MCInst_MC3_r3Inst_XORInst_0_0_U1  ( .A(\Red_MCInst_MC3_v0_1 [0]), 
        .B(\Red_MCInst_MC3_v1_1 [2]), .Z(\MCInst_MC3_r3Inst_XORInst_0_0_n5 )
         );
  XNOR2_X1 \MCInst_MC3_r3Inst_XORInst_0_1_U3  ( .A(
        \MCInst_MC3_r3Inst_XORInst_0_1_n5 ), .B(
        \MCInst_MC3_r3Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[1]) );
  XNOR2_X1 \MCInst_MC3_r3Inst_XORInst_0_1_U2  ( .A(\MCInst_MC3_v3_3 [1]), .B(
        \Red_MCInst_MC3_v2_1 [1]), .ZN(\MCInst_MC3_r3Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \MCInst_MC3_r3Inst_XORInst_0_1_U1  ( .A(\MCInst_MC3_v0_3 [1]), .B(
        \MCInst_MC3_v1_3 [1]), .Z(\MCInst_MC3_r3Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \MCInst_MC3_r3Inst_XORInst_0_2_U3  ( .A(
        \MCInst_MC3_r3Inst_XORInst_0_2_n5 ), .B(
        \MCInst_MC3_r3Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[2]) );
  XNOR2_X1 \MCInst_MC3_r3Inst_XORInst_0_2_U2  ( .A(\MCInst_MC3_v3_3 [2]), .B(
        \MCInst_MC3_v2_3 [2]), .ZN(\MCInst_MC3_r3Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \MCInst_MC3_r3Inst_XORInst_0_2_U1  ( .A(\Red_MCInst_MC3_v0_2 [2]), 
        .B(\Red_MCInst_MC3_v1_2 [1]), .Z(\MCInst_MC3_r3Inst_XORInst_0_2_n5 )
         );
  XNOR2_X1 \MCInst_MC3_r3Inst_XORInst_0_3_U3  ( .A(
        \MCInst_MC3_r3Inst_XORInst_0_3_n5 ), .B(
        \MCInst_MC3_r3Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[3]) );
  XNOR2_X1 \MCInst_MC3_r3Inst_XORInst_0_3_U2  ( .A(\MCInst_MC3_v3_3 [3]), .B(
        \MCInst_MC3_v2_3 [3]), .ZN(\MCInst_MC3_r3Inst_XORInst_0_3_n4 ) );
  XOR2_X1 \MCInst_MC3_r3Inst_XORInst_0_3_U1  ( .A(\MCInst_MC3_v0_3 [3]), .B(
        \MCInst_MC3_v1_3 [3]), .Z(\MCInst_MC3_r3Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_0_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_0_LFInst_0_n2 ), .B(Plaintext[1]), .ZN(
        Red_Plaintext[0]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_0_LFInst_0_U3  ( .A(Plaintext[2]), .B(
        Plaintext[0]), .ZN(\Red_PlaintextInst_LFInst_0_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_0_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_0_LFInst_1_n2 ), .B(Plaintext[1]), .ZN(
        Red_Plaintext[1]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_0_LFInst_1_U3  ( .A(Plaintext[3]), .B(
        Plaintext[0]), .ZN(\Red_PlaintextInst_LFInst_0_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_0_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_0_LFInst_2_n2 ), .B(Plaintext[2]), .ZN(
        Red_Plaintext[2]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_0_LFInst_2_U3  ( .A(Plaintext[3]), .B(
        Plaintext[1]), .ZN(\Red_PlaintextInst_LFInst_0_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_1_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_1_LFInst_0_n2 ), .B(Plaintext[5]), .ZN(
        Red_Plaintext[3]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_1_LFInst_0_U3  ( .A(Plaintext[6]), .B(
        Plaintext[4]), .ZN(\Red_PlaintextInst_LFInst_1_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_1_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_1_LFInst_1_n2 ), .B(Plaintext[5]), .ZN(
        Red_Plaintext[4]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_1_LFInst_1_U3  ( .A(Plaintext[7]), .B(
        Plaintext[4]), .ZN(\Red_PlaintextInst_LFInst_1_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_1_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_1_LFInst_2_n2 ), .B(Plaintext[6]), .ZN(
        Red_Plaintext[5]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_1_LFInst_2_U3  ( .A(Plaintext[7]), .B(
        Plaintext[5]), .ZN(\Red_PlaintextInst_LFInst_1_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_2_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_2_LFInst_0_n2 ), .B(Plaintext[9]), .ZN(
        Red_Plaintext[6]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_2_LFInst_0_U3  ( .A(Plaintext[10]), .B(
        Plaintext[8]), .ZN(\Red_PlaintextInst_LFInst_2_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_2_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_2_LFInst_1_n2 ), .B(Plaintext[9]), .ZN(
        Red_Plaintext[7]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_2_LFInst_1_U3  ( .A(Plaintext[11]), .B(
        Plaintext[8]), .ZN(\Red_PlaintextInst_LFInst_2_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_2_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_2_LFInst_2_n2 ), .B(Plaintext[10]), .ZN(
        Red_Plaintext[8]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_2_LFInst_2_U3  ( .A(Plaintext[11]), .B(
        Plaintext[9]), .ZN(\Red_PlaintextInst_LFInst_2_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_3_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_3_LFInst_0_n2 ), .B(Plaintext[13]), .ZN(
        Red_Plaintext[9]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_3_LFInst_0_U3  ( .A(Plaintext[14]), .B(
        Plaintext[12]), .ZN(\Red_PlaintextInst_LFInst_3_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_3_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_3_LFInst_1_n2 ), .B(Plaintext[13]), .ZN(
        Red_Plaintext[10]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_3_LFInst_1_U3  ( .A(Plaintext[15]), .B(
        Plaintext[12]), .ZN(\Red_PlaintextInst_LFInst_3_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_3_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_3_LFInst_2_n2 ), .B(Plaintext[14]), .ZN(
        Red_Plaintext[11]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_3_LFInst_2_U3  ( .A(Plaintext[15]), .B(
        Plaintext[13]), .ZN(\Red_PlaintextInst_LFInst_3_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_4_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_4_LFInst_0_n2 ), .B(Plaintext[17]), .ZN(
        Red_Plaintext[12]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_4_LFInst_0_U3  ( .A(Plaintext[18]), .B(
        Plaintext[16]), .ZN(\Red_PlaintextInst_LFInst_4_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_4_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_4_LFInst_1_n2 ), .B(Plaintext[17]), .ZN(
        Red_Plaintext[13]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_4_LFInst_1_U3  ( .A(Plaintext[19]), .B(
        Plaintext[16]), .ZN(\Red_PlaintextInst_LFInst_4_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_4_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_4_LFInst_2_n2 ), .B(Plaintext[18]), .ZN(
        Red_Plaintext[14]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_4_LFInst_2_U3  ( .A(Plaintext[19]), .B(
        Plaintext[17]), .ZN(\Red_PlaintextInst_LFInst_4_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_5_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_5_LFInst_0_n2 ), .B(Plaintext[21]), .ZN(
        Red_Plaintext[15]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_5_LFInst_0_U3  ( .A(Plaintext[22]), .B(
        Plaintext[20]), .ZN(\Red_PlaintextInst_LFInst_5_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_5_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_5_LFInst_1_n2 ), .B(Plaintext[21]), .ZN(
        Red_Plaintext[16]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_5_LFInst_1_U3  ( .A(Plaintext[23]), .B(
        Plaintext[20]), .ZN(\Red_PlaintextInst_LFInst_5_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_5_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_5_LFInst_2_n2 ), .B(Plaintext[22]), .ZN(
        Red_Plaintext[17]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_5_LFInst_2_U3  ( .A(Plaintext[23]), .B(
        Plaintext[21]), .ZN(\Red_PlaintextInst_LFInst_5_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_6_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_6_LFInst_0_n2 ), .B(Plaintext[25]), .ZN(
        Red_Plaintext[18]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_6_LFInst_0_U3  ( .A(Plaintext[26]), .B(
        Plaintext[24]), .ZN(\Red_PlaintextInst_LFInst_6_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_6_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_6_LFInst_1_n2 ), .B(Plaintext[25]), .ZN(
        Red_Plaintext[19]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_6_LFInst_1_U3  ( .A(Plaintext[27]), .B(
        Plaintext[24]), .ZN(\Red_PlaintextInst_LFInst_6_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_6_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_6_LFInst_2_n2 ), .B(Plaintext[26]), .ZN(
        Red_Plaintext[20]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_6_LFInst_2_U3  ( .A(Plaintext[27]), .B(
        Plaintext[25]), .ZN(\Red_PlaintextInst_LFInst_6_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_7_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_7_LFInst_0_n2 ), .B(Plaintext[29]), .ZN(
        Red_Plaintext[21]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_7_LFInst_0_U3  ( .A(Plaintext[30]), .B(
        Plaintext[28]), .ZN(\Red_PlaintextInst_LFInst_7_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_7_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_7_LFInst_1_n2 ), .B(Plaintext[29]), .ZN(
        Red_Plaintext[22]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_7_LFInst_1_U3  ( .A(Plaintext[31]), .B(
        Plaintext[28]), .ZN(\Red_PlaintextInst_LFInst_7_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_7_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_7_LFInst_2_n2 ), .B(Plaintext[30]), .ZN(
        Red_Plaintext[23]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_7_LFInst_2_U3  ( .A(Plaintext[31]), .B(
        Plaintext[29]), .ZN(\Red_PlaintextInst_LFInst_7_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_8_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_8_LFInst_0_n2 ), .B(Plaintext[33]), .ZN(
        Red_Plaintext[24]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_8_LFInst_0_U3  ( .A(Plaintext[34]), .B(
        Plaintext[32]), .ZN(\Red_PlaintextInst_LFInst_8_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_8_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_8_LFInst_1_n2 ), .B(Plaintext[33]), .ZN(
        Red_Plaintext[25]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_8_LFInst_1_U3  ( .A(Plaintext[35]), .B(
        Plaintext[32]), .ZN(\Red_PlaintextInst_LFInst_8_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_8_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_8_LFInst_2_n2 ), .B(Plaintext[34]), .ZN(
        Red_Plaintext[26]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_8_LFInst_2_U3  ( .A(Plaintext[35]), .B(
        Plaintext[33]), .ZN(\Red_PlaintextInst_LFInst_8_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_9_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_9_LFInst_0_n2 ), .B(Plaintext[37]), .ZN(
        Red_Plaintext[27]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_9_LFInst_0_U3  ( .A(Plaintext[38]), .B(
        Plaintext[36]), .ZN(\Red_PlaintextInst_LFInst_9_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_9_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_9_LFInst_1_n2 ), .B(Plaintext[37]), .ZN(
        Red_Plaintext[28]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_9_LFInst_1_U3  ( .A(Plaintext[39]), .B(
        Plaintext[36]), .ZN(\Red_PlaintextInst_LFInst_9_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_9_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_9_LFInst_2_n2 ), .B(Plaintext[38]), .ZN(
        Red_Plaintext[29]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_9_LFInst_2_U3  ( .A(Plaintext[39]), .B(
        Plaintext[37]), .ZN(\Red_PlaintextInst_LFInst_9_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_10_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_10_LFInst_0_n2 ), .B(Plaintext[41]), .ZN(
        Red_Plaintext[30]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_10_LFInst_0_U3  ( .A(Plaintext[42]), .B(
        Plaintext[40]), .ZN(\Red_PlaintextInst_LFInst_10_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_10_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_10_LFInst_1_n2 ), .B(Plaintext[41]), .ZN(
        Red_Plaintext[31]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_10_LFInst_1_U3  ( .A(Plaintext[43]), .B(
        Plaintext[40]), .ZN(\Red_PlaintextInst_LFInst_10_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_10_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_10_LFInst_2_n2 ), .B(Plaintext[42]), .ZN(
        Red_Plaintext[32]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_10_LFInst_2_U3  ( .A(Plaintext[43]), .B(
        Plaintext[41]), .ZN(\Red_PlaintextInst_LFInst_10_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_11_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_11_LFInst_0_n2 ), .B(Plaintext[45]), .ZN(
        Red_Plaintext[33]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_11_LFInst_0_U3  ( .A(Plaintext[46]), .B(
        Plaintext[44]), .ZN(\Red_PlaintextInst_LFInst_11_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_11_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_11_LFInst_1_n2 ), .B(Plaintext[45]), .ZN(
        Red_Plaintext[34]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_11_LFInst_1_U3  ( .A(Plaintext[47]), .B(
        Plaintext[44]), .ZN(\Red_PlaintextInst_LFInst_11_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_11_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_11_LFInst_2_n2 ), .B(Plaintext[46]), .ZN(
        Red_Plaintext[35]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_11_LFInst_2_U3  ( .A(Plaintext[47]), .B(
        Plaintext[45]), .ZN(\Red_PlaintextInst_LFInst_11_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_12_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_12_LFInst_0_n2 ), .B(Plaintext[49]), .ZN(
        Red_Plaintext[36]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_12_LFInst_0_U3  ( .A(Plaintext[50]), .B(
        Plaintext[48]), .ZN(\Red_PlaintextInst_LFInst_12_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_12_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_12_LFInst_1_n2 ), .B(Plaintext[49]), .ZN(
        Red_Plaintext[37]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_12_LFInst_1_U3  ( .A(Plaintext[51]), .B(
        Plaintext[48]), .ZN(\Red_PlaintextInst_LFInst_12_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_12_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_12_LFInst_2_n2 ), .B(Plaintext[50]), .ZN(
        Red_Plaintext[38]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_12_LFInst_2_U3  ( .A(Plaintext[51]), .B(
        Plaintext[49]), .ZN(\Red_PlaintextInst_LFInst_12_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_13_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_13_LFInst_0_n2 ), .B(Plaintext[53]), .ZN(
        Red_Plaintext[39]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_13_LFInst_0_U3  ( .A(Plaintext[54]), .B(
        Plaintext[52]), .ZN(\Red_PlaintextInst_LFInst_13_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_13_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_13_LFInst_1_n2 ), .B(Plaintext[53]), .ZN(
        Red_Plaintext[40]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_13_LFInst_1_U3  ( .A(Plaintext[55]), .B(
        Plaintext[52]), .ZN(\Red_PlaintextInst_LFInst_13_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_13_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_13_LFInst_2_n2 ), .B(Plaintext[54]), .ZN(
        Red_Plaintext[41]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_13_LFInst_2_U3  ( .A(Plaintext[55]), .B(
        Plaintext[53]), .ZN(\Red_PlaintextInst_LFInst_13_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_14_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_14_LFInst_0_n2 ), .B(Plaintext[57]), .ZN(
        Red_Plaintext[42]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_14_LFInst_0_U3  ( .A(Plaintext[58]), .B(
        Plaintext[56]), .ZN(\Red_PlaintextInst_LFInst_14_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_14_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_14_LFInst_1_n2 ), .B(Plaintext[57]), .ZN(
        Red_Plaintext[43]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_14_LFInst_1_U3  ( .A(Plaintext[59]), .B(
        Plaintext[56]), .ZN(\Red_PlaintextInst_LFInst_14_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_14_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_14_LFInst_2_n2 ), .B(Plaintext[58]), .ZN(
        Red_Plaintext[44]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_14_LFInst_2_U3  ( .A(Plaintext[59]), .B(
        Plaintext[57]), .ZN(\Red_PlaintextInst_LFInst_14_LFInst_2_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_15_LFInst_0_U4  ( .A(
        \Red_PlaintextInst_LFInst_15_LFInst_0_n2 ), .B(Plaintext[61]), .ZN(
        Red_Plaintext[45]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_15_LFInst_0_U3  ( .A(Plaintext[62]), .B(
        Plaintext[60]), .ZN(\Red_PlaintextInst_LFInst_15_LFInst_0_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_15_LFInst_1_U4  ( .A(
        \Red_PlaintextInst_LFInst_15_LFInst_1_n2 ), .B(Plaintext[61]), .ZN(
        Red_Plaintext[46]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_15_LFInst_1_U3  ( .A(Plaintext[63]), .B(
        Plaintext[60]), .ZN(\Red_PlaintextInst_LFInst_15_LFInst_1_n2 ) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_15_LFInst_2_U4  ( .A(
        \Red_PlaintextInst_LFInst_15_LFInst_2_n2 ), .B(Plaintext[62]), .ZN(
        Red_Plaintext[47]) );
  XNOR2_X1 \Red_PlaintextInst_LFInst_15_LFInst_2_U3  ( .A(Plaintext[63]), .B(
        Plaintext[61]), .ZN(\Red_PlaintextInst_LFInst_15_LFInst_2_n2 ) );
  XOR2_X1 \RedAddKeyXOR_XORInst_0_0_U1  ( .A(Red_Plaintext[0]), .B(
        Red_RoundKey[0]), .Z(Red_AddRoundKeyOutput[0]) );
  XOR2_X1 \RedAddKeyXOR_XORInst_0_1_U1  ( .A(Red_Plaintext[1]), .B(
        Red_RoundKey[1]), .Z(Red_AddRoundKeyOutput[1]) );
  XOR2_X1 \RedAddKeyXOR_XORInst_0_2_U1  ( .A(Red_Plaintext[2]), .B(
        Red_RoundKey[2]), .Z(Red_AddRoundKeyOutput[2]) );
  XOR2_X1 \RedAddKeyXOR_XORInst_1_0_U1  ( .A(Red_Plaintext[3]), .B(
        Red_RoundKey[3]), .Z(Red_AddRoundKeyOutput[3]) );
  XOR2_X1 \RedAddKeyXOR_XORInst_1_1_U1  ( .A(Red_Plaintext[4]), .B(
        Red_RoundKey[4]), .Z(Red_AddRoundKeyOutput[4]) );
  XOR2_X1 \RedAddKeyXOR_XORInst_1_2_U1  ( .A(Red_Plaintext[5]), .B(
        Red_RoundKey[5]), .Z(Red_AddRoundKeyOutput[5]) );
  XOR2_X1 \RedAddKeyXOR_XORInst_2_0_U1  ( .A(Red_Plaintext[6]), .B(
        Red_RoundKey[6]), .Z(Red_AddRoundKeyOutput[6]) );
  XOR2_X1 \RedAddKeyXOR_XORInst_2_1_U1  ( .A(Red_Plaintext[7]), .B(
        Red_RoundKey[7]), .Z(Red_AddRoundKeyOutput[7]) );
  XOR2_X1 \RedAddKeyXOR_XORInst_2_2_U1  ( .A(Red_Plaintext[8]), .B(
        Red_RoundKey[8]), .Z(Red_AddRoundKeyOutput[8]) );
  XOR2_X1 \RedAddKeyXOR_XORInst_3_0_U1  ( .A(Red_Plaintext[9]), .B(
        Red_RoundKey[9]), .Z(Red_AddRoundKeyOutput[9]) );
  XOR2_X1 \RedAddKeyXOR_XORInst_3_1_U1  ( .A(Red_Plaintext[10]), .B(
        Red_RoundKey[10]), .Z(Red_AddRoundKeyOutput[10]) );
  XOR2_X1 \RedAddKeyXOR_XORInst_3_2_U1  ( .A(Red_Plaintext[11]), .B(
        Red_RoundKey[11]), .Z(Red_AddRoundKeyOutput[11]) );
  XOR2_X1 \RedAddKeyXOR_XORInst_4_0_U1  ( .A(Red_Plaintext[12]), .B(
        Red_RoundKey[12]), .Z(Red_AddRoundKeyOutput[12]) );
  XOR2_X1 \RedAddKeyXOR_XORInst_4_1_U1  ( .A(Red_Plaintext[13]), .B(
        Red_RoundKey[13]), .Z(Red_AddRoundKeyOutput[13]) );
  XOR2_X1 \RedAddKeyXOR_XORInst_4_2_U1  ( .A(Red_Plaintext[14]), .B(
        Red_RoundKey[14]), .Z(Red_AddRoundKeyOutput[14]) );
  XOR2_X1 \RedAddKeyXOR_XORInst_5_0_U1  ( .A(Red_Plaintext[15]), .B(
        Red_RoundKey[15]), .Z(Red_AddRoundKeyOutput[15]) );
  XOR2_X1 \RedAddKeyXOR_XORInst_5_1_U1  ( .A(Red_Plaintext[16]), .B(
        Red_RoundKey[16]), .Z(Red_AddRoundKeyOutput[16]) );
  XOR2_X1 \RedAddKeyXOR_XORInst_5_2_U1  ( .A(Red_Plaintext[17]), .B(
        Red_RoundKey[17]), .Z(Red_AddRoundKeyOutput[17]) );
  XOR2_X1 \RedAddKeyXOR_XORInst_6_0_U1  ( .A(Red_Plaintext[18]), .B(
        Red_RoundKey[18]), .Z(Red_AddRoundKeyOutput[18]) );
  XOR2_X1 \RedAddKeyXOR_XORInst_6_1_U1  ( .A(Red_Plaintext[19]), .B(
        Red_RoundKey[19]), .Z(Red_AddRoundKeyOutput[19]) );
  XOR2_X1 \RedAddKeyXOR_XORInst_6_2_U1  ( .A(Red_Plaintext[20]), .B(
        Red_RoundKey[20]), .Z(Red_AddRoundKeyOutput[20]) );
  XOR2_X1 \RedAddKeyXOR_XORInst_7_0_U1  ( .A(Red_Plaintext[21]), .B(
        Red_RoundKey[21]), .Z(Red_AddRoundKeyOutput[21]) );
  XOR2_X1 \RedAddKeyXOR_XORInst_7_1_U1  ( .A(Red_Plaintext[22]), .B(
        Red_RoundKey[22]), .Z(Red_AddRoundKeyOutput[22]) );
  XOR2_X1 \RedAddKeyXOR_XORInst_7_2_U1  ( .A(Red_Plaintext[23]), .B(
        Red_RoundKey[23]), .Z(Red_AddRoundKeyOutput[23]) );
  XOR2_X1 \RedAddKeyXOR_XORInst_8_0_U1  ( .A(Red_Plaintext[24]), .B(
        Red_RoundKey[24]), .Z(Red_AddRoundKeyOutput[24]) );
  XOR2_X1 \RedAddKeyXOR_XORInst_8_1_U1  ( .A(Red_Plaintext[25]), .B(
        Red_RoundKey[25]), .Z(Red_AddRoundKeyOutput[25]) );
  XOR2_X1 \RedAddKeyXOR_XORInst_8_2_U1  ( .A(Red_Plaintext[26]), .B(
        Red_RoundKey[26]), .Z(Red_AddRoundKeyOutput[26]) );
  XOR2_X1 \RedAddKeyXOR_XORInst_9_0_U1  ( .A(Red_Plaintext[27]), .B(
        Red_RoundKey[27]), .Z(Red_AddRoundKeyOutput[27]) );
  XOR2_X1 \RedAddKeyXOR_XORInst_9_1_U1  ( .A(Red_Plaintext[28]), .B(
        Red_RoundKey[28]), .Z(Red_AddRoundKeyOutput[28]) );
  XOR2_X1 \RedAddKeyXOR_XORInst_9_2_U1  ( .A(Red_Plaintext[29]), .B(
        Red_RoundKey[29]), .Z(Red_AddRoundKeyOutput[29]) );
  XOR2_X1 \RedAddKeyXOR_XORInst_10_0_U1  ( .A(Red_Plaintext[30]), .B(
        Red_RoundKey[30]), .Z(Red_AddRoundKeyOutput[30]) );
  XOR2_X1 \RedAddKeyXOR_XORInst_10_1_U1  ( .A(Red_Plaintext[31]), .B(
        Red_RoundKey[31]), .Z(Red_AddRoundKeyOutput[31]) );
  XOR2_X1 \RedAddKeyXOR_XORInst_10_2_U1  ( .A(Red_Plaintext[32]), .B(
        Red_RoundKey[32]), .Z(Red_AddRoundKeyOutput[32]) );
  XOR2_X1 \RedAddKeyXOR_XORInst_11_0_U1  ( .A(Red_Plaintext[33]), .B(
        Red_RoundKey[33]), .Z(Red_AddRoundKeyOutput[33]) );
  XOR2_X1 \RedAddKeyXOR_XORInst_11_1_U1  ( .A(Red_Plaintext[34]), .B(
        Red_RoundKey[34]), .Z(Red_AddRoundKeyOutput[34]) );
  XOR2_X1 \RedAddKeyXOR_XORInst_11_2_U1  ( .A(Red_Plaintext[35]), .B(
        Red_RoundKey[35]), .Z(Red_AddRoundKeyOutput[35]) );
  XOR2_X1 \RedAddKeyXOR_XORInst_12_0_U1  ( .A(Red_Plaintext[36]), .B(
        Red_RoundKey[36]), .Z(Red_AddRoundKeyOutput[36]) );
  XOR2_X1 \RedAddKeyXOR_XORInst_12_1_U1  ( .A(Red_Plaintext[37]), .B(
        Red_RoundKey[37]), .Z(Red_AddRoundKeyOutput[37]) );
  XOR2_X1 \RedAddKeyXOR_XORInst_12_2_U1  ( .A(Red_Plaintext[38]), .B(
        Red_RoundKey[38]), .Z(Red_AddRoundKeyOutput[38]) );
  XOR2_X1 \RedAddKeyXOR_XORInst_13_0_U1  ( .A(Red_Plaintext[39]), .B(
        Red_RoundKey[39]), .Z(Red_AddRoundKeyOutput[39]) );
  XOR2_X1 \RedAddKeyXOR_XORInst_13_1_U1  ( .A(Red_Plaintext[40]), .B(
        Red_RoundKey[40]), .Z(Red_AddRoundKeyOutput[40]) );
  XOR2_X1 \RedAddKeyXOR_XORInst_13_2_U1  ( .A(Red_Plaintext[41]), .B(
        Red_RoundKey[41]), .Z(Red_AddRoundKeyOutput[41]) );
  XOR2_X1 \RedAddKeyXOR_XORInst_14_0_U1  ( .A(Red_Plaintext[42]), .B(
        Red_RoundKey[42]), .Z(Red_AddRoundKeyOutput[42]) );
  XOR2_X1 \RedAddKeyXOR_XORInst_14_1_U1  ( .A(Red_Plaintext[43]), .B(
        Red_RoundKey[43]), .Z(Red_AddRoundKeyOutput[43]) );
  XOR2_X1 \RedAddKeyXOR_XORInst_14_2_U1  ( .A(Red_Plaintext[44]), .B(
        Red_RoundKey[44]), .Z(Red_AddRoundKeyOutput[44]) );
  XOR2_X1 \RedAddKeyXOR_XORInst_15_0_U1  ( .A(Red_Plaintext[45]), .B(
        Red_RoundKey[45]), .Z(Red_AddRoundKeyOutput[45]) );
  XOR2_X1 \RedAddKeyXOR_XORInst_15_1_U1  ( .A(Red_Plaintext[46]), .B(
        Red_RoundKey[46]), .Z(Red_AddRoundKeyOutput[46]) );
  XOR2_X1 \RedAddKeyXOR_XORInst_15_2_U1  ( .A(Red_Plaintext[47]), .B(
        Red_RoundKey[47]), .Z(Red_AddRoundKeyOutput[47]) );
  XOR2_X1 \Red_MCInst_MC0_v0_2Inst_0_U3  ( .A(\MCInst_MC0_v0_3 [3]), .B(
        \Red_MCInst_MC0_v0_1 [0]), .Z(\Red_MCInst_MC0_v0_2 [0]) );
  XOR2_X1 \Red_MCInst_MC0_v0_3Inst_0_U3  ( .A(\Red_MCInst_MC0_v0_0 [0]), .B(
        \Red_MCInst_MC0_v0_2 [2]), .Z(\Red_MCInst_MC0_v0_3 [0]) );
  XNOR2_X1 \Red_MCInst_MC0_v1_0Inst_0_U4  ( .A(\Red_MCInst_MC0_v1_0Inst_0_n2 ), 
        .B(\Red_MCInst_MC0_v1_2 [1]), .ZN(\Red_MCInst_MC0_v1_0 [0]) );
  XNOR2_X1 \Red_MCInst_MC0_v1_0Inst_0_U3  ( .A(\MCInst_MC0_v1_3 [3]), .B(
        \MCInst_MC0_v1_0 [0]), .ZN(\Red_MCInst_MC0_v1_0Inst_0_n2 ) );
  XOR2_X1 \Red_MCInst_MC0_v1_2Inst_0_U3  ( .A(\Red_MCInst_MC0_v1_2 [1]), .B(
        \Red_MCInst_MC0_v1_1 [2]), .Z(\Red_MCInst_MC0_v1_2 [0]) );
  XOR2_X1 \Red_MCInst_MC0_v1_3Inst_0_U3  ( .A(\MCInst_MC0_v1_0 [0]), .B(
        \Red_MCInst_MC0_v1_2 [1]), .Z(\Red_MCInst_MC0_v1_3 [0]) );
  XOR2_X1 \Red_MCInst_MC0_v2_0Inst_0_U3  ( .A(\Red_MCInst_MC0_v2_1 [1]), .B(
        \MCInst_MC0_v2_0 [2]), .Z(\Red_MCInst_MC0_v2_0 [0]) );
  XOR2_X1 \Red_MCInst_MC0_v2_1Inst_0_U3  ( .A(\MCInst_MC0_v2_0 [2]), .B(
        \MCInst_MC0_v2_0 [3]), .Z(\Red_MCInst_MC0_v2_1 [0]) );
  XNOR2_X1 \Red_MCInst_MC0_v2_2Inst_0_U4  ( .A(\Red_MCInst_MC0_v2_2Inst_0_n2 ), 
        .B(\MCInst_MC0_v2_0 [2]), .ZN(\Red_MCInst_MC0_v2_2 [0]) );
  XNOR2_X1 \Red_MCInst_MC0_v2_2Inst_0_U3  ( .A(\Red_MCInst_MC0_v2_2 [1]), .B(
        \Red_MCInst_MC0_v2_1 [1]), .ZN(\Red_MCInst_MC0_v2_2Inst_0_n2 ) );
  XNOR2_X1 \Red_MCInst_MC0_v2_3Inst_0_U4  ( .A(\Red_MCInst_MC0_v2_3Inst_0_n2 ), 
        .B(\MCInst_MC0_v2_0 [3]), .ZN(\Red_MCInst_MC0_v2_3 [0]) );
  XNOR2_X1 \Red_MCInst_MC0_v2_3Inst_0_U3  ( .A(\Red_MCInst_MC0_v2_2 [1]), .B(
        \Red_MCInst_MC0_v2_1 [1]), .ZN(\Red_MCInst_MC0_v2_3Inst_0_n2 ) );
  XOR2_X1 \Red_MCInst_MC0_v3_0Inst_0_U3  ( .A(\MCInst_MC0_v3_2 [3]), .B(
        \Red_MCInst_MC0_v3_3 [2]), .Z(\Red_MCInst_MC0_v3_0 [0]) );
  XNOR2_X1 \Red_MCInst_MC0_v3_2Inst_0_U5  ( .A(\Red_MCInst_MC0_v3_2Inst_0_n4 ), 
        .B(\Red_MCInst_MC0_v3_2Inst_0_n3 ), .ZN(\Red_MCInst_MC0_v3_2 [0]) );
  XNOR2_X1 \Red_MCInst_MC0_v3_2Inst_0_U4  ( .A(\Red_MCInst_MC0_v3_3 [2]), .B(
        \MCInst_MC0_v3_2 [3]), .ZN(\Red_MCInst_MC0_v3_2Inst_0_n3 ) );
  XOR2_X1 \Red_MCInst_MC0_v3_2Inst_0_U3  ( .A(\MCInst_MC0_v3_0 [3]), .B(
        \Red_MCInst_MC0_v3_1 [2]), .Z(\Red_MCInst_MC0_v3_2Inst_0_n4 ) );
  XOR2_X1 \Red_MCInst_MC0_v3_3Inst_0_U3  ( .A(\MCInst_MC0_v3_0 [3]), .B(
        \Red_MCInst_MC0_v3_1 [2]), .Z(\Red_MCInst_MC0_v3_3 [0]) );
  XOR2_X1 \Red_MCInst_MC0_v0_0Inst_1_U3  ( .A(\Red_MCInst_MC0_v0_2 [2]), .B(
        \Red_MCInst_MC0_v0_1 [0]), .Z(\Red_MCInst_MC0_v0_0 [1]) );
  XNOR2_X1 \Red_MCInst_MC0_v0_1Inst_1_U4  ( .A(\Red_MCInst_MC0_v0_1Inst_1_n2 ), 
        .B(\MCInst_MC0_v0_3 [3]), .ZN(\Red_MCInst_MC0_v0_1 [1]) );
  XNOR2_X1 \Red_MCInst_MC0_v0_1Inst_1_U3  ( .A(\Red_MCInst_MC0_v0_1 [0]), .B(
        \Red_MCInst_MC0_v0_0 [0]), .ZN(\Red_MCInst_MC0_v0_1Inst_1_n2 ) );
  XOR2_X1 \Red_MCInst_MC0_v0_2Inst_1_U3  ( .A(\Red_MCInst_MC0_v0_0 [0]), .B(
        \Red_MCInst_MC0_v0_2 [2]), .Z(\Red_MCInst_MC0_v0_2 [1]) );
  XOR2_X1 \Red_MCInst_MC0_v0_3Inst_1_U3  ( .A(\Red_MCInst_MC0_v0_0 [0]), .B(
        \MCInst_MC0_v0_3 [3]), .Z(\Red_MCInst_MC0_v0_3 [1]) );
  XNOR2_X1 \Red_MCInst_MC0_v1_0Inst_1_U4  ( .A(\Red_MCInst_MC0_v1_0Inst_1_n2 ), 
        .B(\Red_MCInst_MC0_v1_2 [1]), .ZN(\Red_MCInst_MC0_v1_0 [1]) );
  XNOR2_X1 \Red_MCInst_MC0_v1_0Inst_1_U3  ( .A(\Red_MCInst_MC0_v1_1 [2]), .B(
        \MCInst_MC0_v1_0 [0]), .ZN(\Red_MCInst_MC0_v1_0Inst_1_n2 ) );
  XNOR2_X1 \Red_MCInst_MC0_v1_1Inst_1_U5  ( .A(\Red_MCInst_MC0_v1_1Inst_1_n4 ), 
        .B(\Red_MCInst_MC0_v1_1Inst_1_n3 ), .ZN(\Red_MCInst_MC0_v1_1 [1]) );
  XNOR2_X1 \Red_MCInst_MC0_v1_1Inst_1_U4  ( .A(\Red_MCInst_MC0_v1_2 [1]), .B(
        \MCInst_MC0_v1_0 [0]), .ZN(\Red_MCInst_MC0_v1_1Inst_1_n3 ) );
  XOR2_X1 \Red_MCInst_MC0_v1_1Inst_1_U3  ( .A(\MCInst_MC0_v1_3 [3]), .B(
        \Red_MCInst_MC0_v1_1 [2]), .Z(\Red_MCInst_MC0_v1_1Inst_1_n4 ) );
  XOR2_X1 \Red_MCInst_MC0_v1_3Inst_1_U3  ( .A(\MCInst_MC0_v1_0 [0]), .B(
        \MCInst_MC0_v1_3 [3]), .Z(\Red_MCInst_MC0_v1_3 [1]) );
  XOR2_X1 \Red_MCInst_MC0_v2_0Inst_1_U3  ( .A(\Red_MCInst_MC0_v2_1 [1]), .B(
        \MCInst_MC0_v2_0 [3]), .Z(\Red_MCInst_MC0_v2_0 [1]) );
  XOR2_X1 \Red_MCInst_MC0_v2_3Inst_1_U3  ( .A(\Red_MCInst_MC0_v2_1 [1]), .B(
        \Red_MCInst_MC0_v2_2 [1]), .Z(\Red_MCInst_MC0_v2_3 [1]) );
  XOR2_X1 \Red_MCInst_MC0_v3_0Inst_1_U3  ( .A(\MCInst_MC0_v3_2 [3]), .B(
        \MCInst_MC0_v3_0 [3]), .Z(\Red_MCInst_MC0_v3_0 [1]) );
  XNOR2_X1 \Red_MCInst_MC0_v3_1Inst_1_U5  ( .A(\Red_MCInst_MC0_v3_1Inst_1_n4 ), 
        .B(\Red_MCInst_MC0_v3_1Inst_1_n3 ), .ZN(\Red_MCInst_MC0_v3_1 [1]) );
  XNOR2_X1 \Red_MCInst_MC0_v3_1Inst_1_U4  ( .A(\Red_MCInst_MC0_v3_3 [2]), .B(
        \MCInst_MC0_v3_2 [3]), .ZN(\Red_MCInst_MC0_v3_1Inst_1_n3 ) );
  XOR2_X1 \Red_MCInst_MC0_v3_1Inst_1_U3  ( .A(\MCInst_MC0_v3_0 [3]), .B(
        \Red_MCInst_MC0_v3_1 [2]), .Z(\Red_MCInst_MC0_v3_1Inst_1_n4 ) );
  XOR2_X1 \Red_MCInst_MC0_v3_2Inst_1_U3  ( .A(\Red_MCInst_MC0_v3_3 [2]), .B(
        \MCInst_MC0_v3_0 [3]), .Z(\Red_MCInst_MC0_v3_2 [1]) );
  XOR2_X1 \Red_MCInst_MC0_v3_3Inst_1_U3  ( .A(\MCInst_MC0_v3_2 [3]), .B(
        \Red_MCInst_MC0_v3_3 [2]), .Z(\Red_MCInst_MC0_v3_3 [1]) );
  XNOR2_X1 \Red_MCInst_MC0_v0_0Inst_2_U4  ( .A(\Red_MCInst_MC0_v0_0Inst_2_n2 ), 
        .B(\Red_MCInst_MC0_v0_2 [2]), .ZN(\Red_MCInst_MC0_v0_0 [2]) );
  XNOR2_X1 \Red_MCInst_MC0_v0_0Inst_2_U3  ( .A(\MCInst_MC0_v0_3 [3]), .B(
        \Red_MCInst_MC0_v0_0 [0]), .ZN(\Red_MCInst_MC0_v0_0Inst_2_n2 ) );
  XOR2_X1 \Red_MCInst_MC0_v0_1Inst_2_U3  ( .A(\Red_MCInst_MC0_v0_0 [0]), .B(
        \Red_MCInst_MC0_v0_2 [2]), .Z(\Red_MCInst_MC0_v0_1 [2]) );
  XNOR2_X1 \Red_MCInst_MC0_v0_3Inst_2_U5  ( .A(\Red_MCInst_MC0_v0_3Inst_2_n4 ), 
        .B(\Red_MCInst_MC0_v0_3Inst_2_n3 ), .ZN(\Red_MCInst_MC0_v0_3 [2]) );
  XNOR2_X1 \Red_MCInst_MC0_v0_3Inst_2_U4  ( .A(\Red_MCInst_MC0_v0_2 [2]), .B(
        \Red_MCInst_MC0_v0_0 [0]), .ZN(\Red_MCInst_MC0_v0_3Inst_2_n3 ) );
  XOR2_X1 \Red_MCInst_MC0_v0_3Inst_2_U3  ( .A(\MCInst_MC0_v0_3 [3]), .B(
        \Red_MCInst_MC0_v0_1 [0]), .Z(\Red_MCInst_MC0_v0_3Inst_2_n4 ) );
  XNOR2_X1 \Red_MCInst_MC0_v1_0Inst_2_U4  ( .A(\Red_MCInst_MC0_v1_0Inst_2_n2 ), 
        .B(\MCInst_MC0_v1_3 [3]), .ZN(\Red_MCInst_MC0_v1_0 [2]) );
  XNOR2_X1 \Red_MCInst_MC0_v1_0Inst_2_U3  ( .A(\Red_MCInst_MC0_v1_1 [2]), .B(
        \Red_MCInst_MC0_v1_2 [1]), .ZN(\Red_MCInst_MC0_v1_0Inst_2_n2 ) );
  XNOR2_X1 \Red_MCInst_MC0_v1_2Inst_2_U4  ( .A(\Red_MCInst_MC0_v1_2Inst_2_n2 ), 
        .B(\Red_MCInst_MC0_v1_2 [1]), .ZN(\Red_MCInst_MC0_v1_2 [2]) );
  XNOR2_X1 \Red_MCInst_MC0_v1_2Inst_2_U3  ( .A(\Red_MCInst_MC0_v1_1 [2]), .B(
        \MCInst_MC0_v1_0 [0]), .ZN(\Red_MCInst_MC0_v1_2Inst_2_n2 ) );
  XNOR2_X1 \Red_MCInst_MC0_v1_3Inst_2_U5  ( .A(\Red_MCInst_MC0_v1_3Inst_2_n4 ), 
        .B(\Red_MCInst_MC0_v1_3Inst_2_n3 ), .ZN(\Red_MCInst_MC0_v1_3 [2]) );
  XNOR2_X1 \Red_MCInst_MC0_v1_3Inst_2_U4  ( .A(\Red_MCInst_MC0_v1_2 [1]), .B(
        \MCInst_MC0_v1_0 [0]), .ZN(\Red_MCInst_MC0_v1_3Inst_2_n3 ) );
  XOR2_X1 \Red_MCInst_MC0_v1_3Inst_2_U3  ( .A(\MCInst_MC0_v1_3 [3]), .B(
        \Red_MCInst_MC0_v1_1 [2]), .Z(\Red_MCInst_MC0_v1_3Inst_2_n4 ) );
  XNOR2_X1 \Red_MCInst_MC0_v2_0Inst_2_U5  ( .A(\Red_MCInst_MC0_v2_0Inst_2_n4 ), 
        .B(\Red_MCInst_MC0_v2_0Inst_2_n3 ), .ZN(\Red_MCInst_MC0_v2_0 [2]) );
  XNOR2_X1 \Red_MCInst_MC0_v2_0Inst_2_U4  ( .A(\MCInst_MC0_v2_0 [2]), .B(
        \Red_MCInst_MC0_v2_1 [1]), .ZN(\Red_MCInst_MC0_v2_0Inst_2_n3 ) );
  XOR2_X1 \Red_MCInst_MC0_v2_0Inst_2_U3  ( .A(\MCInst_MC0_v2_0 [3]), .B(
        \Red_MCInst_MC0_v2_2 [1]), .Z(\Red_MCInst_MC0_v2_0Inst_2_n4 ) );
  XOR2_X1 \Red_MCInst_MC0_v2_1Inst_2_U3  ( .A(\Red_MCInst_MC0_v2_1 [1]), .B(
        \Red_MCInst_MC0_v2_2 [1]), .Z(\Red_MCInst_MC0_v2_1 [2]) );
  XOR2_X1 \Red_MCInst_MC0_v2_2Inst_2_U3  ( .A(\MCInst_MC0_v2_0 [3]), .B(
        \Red_MCInst_MC0_v2_2 [1]), .Z(\Red_MCInst_MC0_v2_2 [2]) );
  XOR2_X1 \Red_MCInst_MC0_v2_3Inst_2_U3  ( .A(\Red_MCInst_MC0_v2_1 [1]), .B(
        \MCInst_MC0_v2_0 [3]), .Z(\Red_MCInst_MC0_v2_3 [2]) );
  XNOR2_X1 \Red_MCInst_MC0_v3_0Inst_2_U5  ( .A(\Red_MCInst_MC0_v3_0Inst_2_n4 ), 
        .B(\Red_MCInst_MC0_v3_0Inst_2_n3 ), .ZN(\Red_MCInst_MC0_v3_0 [2]) );
  XNOR2_X1 \Red_MCInst_MC0_v3_0Inst_2_U4  ( .A(\Red_MCInst_MC0_v3_3 [2]), .B(
        \MCInst_MC0_v3_2 [3]), .ZN(\Red_MCInst_MC0_v3_0Inst_2_n3 ) );
  XOR2_X1 \Red_MCInst_MC0_v3_0Inst_2_U3  ( .A(\MCInst_MC0_v3_0 [3]), .B(
        \Red_MCInst_MC0_v3_1 [2]), .Z(\Red_MCInst_MC0_v3_0Inst_2_n4 ) );
  XNOR2_X1 \Red_MCInst_MC0_v3_2Inst_2_U4  ( .A(\Red_MCInst_MC0_v3_2Inst_2_n2 ), 
        .B(\MCInst_MC0_v3_0 [3]), .ZN(\Red_MCInst_MC0_v3_2 [2]) );
  XNOR2_X1 \Red_MCInst_MC0_v3_2Inst_2_U3  ( .A(\Red_MCInst_MC0_v3_1 [2]), .B(
        \MCInst_MC0_v3_2 [3]), .ZN(\Red_MCInst_MC0_v3_2Inst_2_n2 ) );
  XNOR2_X1 \Red_MCInst_MC0_r0Inst_XORInst_0_0_U3  ( .A(
        \Red_MCInst_MC0_r0Inst_XORInst_0_0_n5 ), .B(
        \Red_MCInst_MC0_r0Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback[45]) );
  XNOR2_X1 \Red_MCInst_MC0_r0Inst_XORInst_0_0_U2  ( .A(
        \Red_MCInst_MC0_v3_0 [0]), .B(\Red_MCInst_MC0_v2_0 [0]), .ZN(
        \Red_MCInst_MC0_r0Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \Red_MCInst_MC0_r0Inst_XORInst_0_0_U1  ( .A(\Red_MCInst_MC0_v0_0 [0]), .B(\Red_MCInst_MC0_v1_0 [0]), .Z(\Red_MCInst_MC0_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \Red_MCInst_MC0_r0Inst_XORInst_0_1_U3  ( .A(
        \Red_MCInst_MC0_r0Inst_XORInst_0_1_n5 ), .B(
        \Red_MCInst_MC0_r0Inst_XORInst_0_1_n4 ), .ZN(Red_Feedback[46]) );
  XNOR2_X1 \Red_MCInst_MC0_r0Inst_XORInst_0_1_U2  ( .A(
        \Red_MCInst_MC0_v3_0 [1]), .B(\Red_MCInst_MC0_v2_0 [1]), .ZN(
        \Red_MCInst_MC0_r0Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \Red_MCInst_MC0_r0Inst_XORInst_0_1_U1  ( .A(\Red_MCInst_MC0_v0_0 [1]), .B(\Red_MCInst_MC0_v1_0 [1]), .Z(\Red_MCInst_MC0_r0Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \Red_MCInst_MC0_r0Inst_XORInst_0_2_U3  ( .A(
        \Red_MCInst_MC0_r0Inst_XORInst_0_2_n5 ), .B(
        \Red_MCInst_MC0_r0Inst_XORInst_0_2_n4 ), .ZN(Red_Feedback[47]) );
  XNOR2_X1 \Red_MCInst_MC0_r0Inst_XORInst_0_2_U2  ( .A(
        \Red_MCInst_MC0_v3_0 [2]), .B(\Red_MCInst_MC0_v2_0 [2]), .ZN(
        \Red_MCInst_MC0_r0Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \Red_MCInst_MC0_r0Inst_XORInst_0_2_U1  ( .A(\Red_MCInst_MC0_v0_0 [2]), .B(\Red_MCInst_MC0_v1_0 [2]), .Z(\Red_MCInst_MC0_r0Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \Red_MCInst_MC0_r1Inst_XORInst_0_0_U3  ( .A(
        \Red_MCInst_MC0_r1Inst_XORInst_0_0_n5 ), .B(
        \Red_MCInst_MC0_r1Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback[33]) );
  XNOR2_X1 \Red_MCInst_MC0_r1Inst_XORInst_0_0_U2  ( .A(
        \Red_MCInst_MC0_v3_3 [2]), .B(\Red_MCInst_MC0_v2_1 [0]), .ZN(
        \Red_MCInst_MC0_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \Red_MCInst_MC0_r1Inst_XORInst_0_0_U1  ( .A(\Red_MCInst_MC0_v0_1 [0]), .B(\Red_MCInst_MC0_v1_2 [1]), .Z(\Red_MCInst_MC0_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \Red_MCInst_MC0_r1Inst_XORInst_0_1_U3  ( .A(
        \Red_MCInst_MC0_r1Inst_XORInst_0_1_n5 ), .B(
        \Red_MCInst_MC0_r1Inst_XORInst_0_1_n4 ), .ZN(Red_Feedback[34]) );
  XNOR2_X1 \Red_MCInst_MC0_r1Inst_XORInst_0_1_U2  ( .A(
        \Red_MCInst_MC0_v3_1 [1]), .B(\Red_MCInst_MC0_v2_1 [1]), .ZN(
        \Red_MCInst_MC0_r1Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \Red_MCInst_MC0_r1Inst_XORInst_0_1_U1  ( .A(\Red_MCInst_MC0_v0_1 [1]), .B(\Red_MCInst_MC0_v1_1 [1]), .Z(\Red_MCInst_MC0_r1Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \Red_MCInst_MC0_r1Inst_XORInst_0_2_U3  ( .A(
        \Red_MCInst_MC0_r1Inst_XORInst_0_2_n5 ), .B(
        \Red_MCInst_MC0_r1Inst_XORInst_0_2_n4 ), .ZN(Red_Feedback[35]) );
  XNOR2_X1 \Red_MCInst_MC0_r1Inst_XORInst_0_2_U2  ( .A(
        \Red_MCInst_MC0_v3_1 [2]), .B(\Red_MCInst_MC0_v2_1 [2]), .ZN(
        \Red_MCInst_MC0_r1Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \Red_MCInst_MC0_r1Inst_XORInst_0_2_U1  ( .A(\Red_MCInst_MC0_v0_1 [2]), .B(\Red_MCInst_MC0_v1_1 [2]), .Z(\Red_MCInst_MC0_r1Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \Red_MCInst_MC0_r2Inst_XORInst_0_0_U3  ( .A(
        \Red_MCInst_MC0_r2Inst_XORInst_0_0_n5 ), .B(
        \Red_MCInst_MC0_r2Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback[21]) );
  XNOR2_X1 \Red_MCInst_MC0_r2Inst_XORInst_0_0_U2  ( .A(
        \Red_MCInst_MC0_v3_2 [0]), .B(\Red_MCInst_MC0_v2_2 [0]), .ZN(
        \Red_MCInst_MC0_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \Red_MCInst_MC0_r2Inst_XORInst_0_0_U1  ( .A(\Red_MCInst_MC0_v0_2 [0]), .B(\Red_MCInst_MC0_v1_2 [0]), .Z(\Red_MCInst_MC0_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \Red_MCInst_MC0_r2Inst_XORInst_0_1_U3  ( .A(
        \Red_MCInst_MC0_r2Inst_XORInst_0_1_n5 ), .B(
        \Red_MCInst_MC0_r2Inst_XORInst_0_1_n4 ), .ZN(Red_Feedback[22]) );
  XNOR2_X1 \Red_MCInst_MC0_r2Inst_XORInst_0_1_U2  ( .A(
        \Red_MCInst_MC0_v3_2 [1]), .B(\Red_MCInst_MC0_v2_2 [1]), .ZN(
        \Red_MCInst_MC0_r2Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \Red_MCInst_MC0_r2Inst_XORInst_0_1_U1  ( .A(\Red_MCInst_MC0_v0_2 [1]), .B(\Red_MCInst_MC0_v1_2 [1]), .Z(\Red_MCInst_MC0_r2Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \Red_MCInst_MC0_r2Inst_XORInst_0_2_U3  ( .A(
        \Red_MCInst_MC0_r2Inst_XORInst_0_2_n5 ), .B(
        \Red_MCInst_MC0_r2Inst_XORInst_0_2_n4 ), .ZN(Red_Feedback[23]) );
  XNOR2_X1 \Red_MCInst_MC0_r2Inst_XORInst_0_2_U2  ( .A(
        \Red_MCInst_MC0_v3_2 [2]), .B(\Red_MCInst_MC0_v2_2 [2]), .ZN(
        \Red_MCInst_MC0_r2Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \Red_MCInst_MC0_r2Inst_XORInst_0_2_U1  ( .A(\Red_MCInst_MC0_v0_2 [2]), .B(\Red_MCInst_MC0_v1_2 [2]), .Z(\Red_MCInst_MC0_r2Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \Red_MCInst_MC0_r3Inst_XORInst_0_0_U3  ( .A(
        \Red_MCInst_MC0_r3Inst_XORInst_0_0_n5 ), .B(
        \Red_MCInst_MC0_r3Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback[9]) );
  XNOR2_X1 \Red_MCInst_MC0_r3Inst_XORInst_0_0_U2  ( .A(
        \Red_MCInst_MC0_v3_3 [0]), .B(\Red_MCInst_MC0_v2_3 [0]), .ZN(
        \Red_MCInst_MC0_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \Red_MCInst_MC0_r3Inst_XORInst_0_0_U1  ( .A(\Red_MCInst_MC0_v0_3 [0]), .B(\Red_MCInst_MC0_v1_3 [0]), .Z(\Red_MCInst_MC0_r3Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \Red_MCInst_MC0_r3Inst_XORInst_0_1_U3  ( .A(
        \Red_MCInst_MC0_r3Inst_XORInst_0_1_n5 ), .B(
        \Red_MCInst_MC0_r3Inst_XORInst_0_1_n4 ), .ZN(Red_Feedback[10]) );
  XNOR2_X1 \Red_MCInst_MC0_r3Inst_XORInst_0_1_U2  ( .A(
        \Red_MCInst_MC0_v3_3 [1]), .B(\Red_MCInst_MC0_v2_3 [1]), .ZN(
        \Red_MCInst_MC0_r3Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \Red_MCInst_MC0_r3Inst_XORInst_0_1_U1  ( .A(\Red_MCInst_MC0_v0_3 [1]), .B(\Red_MCInst_MC0_v1_3 [1]), .Z(\Red_MCInst_MC0_r3Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \Red_MCInst_MC0_r3Inst_XORInst_0_2_U3  ( .A(
        \Red_MCInst_MC0_r3Inst_XORInst_0_2_n5 ), .B(
        \Red_MCInst_MC0_r3Inst_XORInst_0_2_n4 ), .ZN(Red_Feedback[11]) );
  XNOR2_X1 \Red_MCInst_MC0_r3Inst_XORInst_0_2_U2  ( .A(
        \Red_MCInst_MC0_v3_3 [2]), .B(\Red_MCInst_MC0_v2_3 [2]), .ZN(
        \Red_MCInst_MC0_r3Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \Red_MCInst_MC0_r3Inst_XORInst_0_2_U1  ( .A(\Red_MCInst_MC0_v0_3 [2]), .B(\Red_MCInst_MC0_v1_3 [2]), .Z(\Red_MCInst_MC0_r3Inst_XORInst_0_2_n5 ) );
  XOR2_X1 \Red_MCInst_MC1_v0_2Inst_0_U3  ( .A(\MCInst_MC1_v0_3 [3]), .B(
        \Red_MCInst_MC1_v0_1 [0]), .Z(\Red_MCInst_MC1_v0_2 [0]) );
  XOR2_X1 \Red_MCInst_MC1_v0_3Inst_0_U3  ( .A(\Red_MCInst_MC1_v0_0 [0]), .B(
        \Red_MCInst_MC1_v0_2 [2]), .Z(\Red_MCInst_MC1_v0_3 [0]) );
  XNOR2_X1 \Red_MCInst_MC1_v1_0Inst_0_U4  ( .A(\Red_MCInst_MC1_v1_0Inst_0_n2 ), 
        .B(\Red_MCInst_MC1_v1_2 [1]), .ZN(\Red_MCInst_MC1_v1_0 [0]) );
  XNOR2_X1 \Red_MCInst_MC1_v1_0Inst_0_U3  ( .A(\MCInst_MC1_v1_3 [3]), .B(
        \MCInst_MC1_v1_0 [0]), .ZN(\Red_MCInst_MC1_v1_0Inst_0_n2 ) );
  XOR2_X1 \Red_MCInst_MC1_v1_2Inst_0_U3  ( .A(\Red_MCInst_MC1_v1_2 [1]), .B(
        \Red_MCInst_MC1_v1_1 [2]), .Z(\Red_MCInst_MC1_v1_2 [0]) );
  XOR2_X1 \Red_MCInst_MC1_v1_3Inst_0_U3  ( .A(\MCInst_MC1_v1_0 [0]), .B(
        \Red_MCInst_MC1_v1_2 [1]), .Z(\Red_MCInst_MC1_v1_3 [0]) );
  XOR2_X1 \Red_MCInst_MC1_v2_0Inst_0_U3  ( .A(\Red_MCInst_MC1_v2_1 [1]), .B(
        \MCInst_MC1_v2_0 [2]), .Z(\Red_MCInst_MC1_v2_0 [0]) );
  XOR2_X1 \Red_MCInst_MC1_v2_1Inst_0_U3  ( .A(\MCInst_MC1_v2_0 [2]), .B(
        \MCInst_MC1_v2_0 [3]), .Z(\Red_MCInst_MC1_v2_1 [0]) );
  XNOR2_X1 \Red_MCInst_MC1_v2_2Inst_0_U4  ( .A(\Red_MCInst_MC1_v2_2Inst_0_n2 ), 
        .B(\MCInst_MC1_v2_0 [2]), .ZN(\Red_MCInst_MC1_v2_2 [0]) );
  XNOR2_X1 \Red_MCInst_MC1_v2_2Inst_0_U3  ( .A(\Red_MCInst_MC1_v2_2 [1]), .B(
        \Red_MCInst_MC1_v2_1 [1]), .ZN(\Red_MCInst_MC1_v2_2Inst_0_n2 ) );
  XNOR2_X1 \Red_MCInst_MC1_v2_3Inst_0_U4  ( .A(\Red_MCInst_MC1_v2_3Inst_0_n2 ), 
        .B(\MCInst_MC1_v2_0 [3]), .ZN(\Red_MCInst_MC1_v2_3 [0]) );
  XNOR2_X1 \Red_MCInst_MC1_v2_3Inst_0_U3  ( .A(\Red_MCInst_MC1_v2_2 [1]), .B(
        \Red_MCInst_MC1_v2_1 [1]), .ZN(\Red_MCInst_MC1_v2_3Inst_0_n2 ) );
  XOR2_X1 \Red_MCInst_MC1_v3_0Inst_0_U3  ( .A(\MCInst_MC1_v3_2 [3]), .B(
        \Red_MCInst_MC1_v3_3 [2]), .Z(\Red_MCInst_MC1_v3_0 [0]) );
  XNOR2_X1 \Red_MCInst_MC1_v3_2Inst_0_U5  ( .A(\Red_MCInst_MC1_v3_2Inst_0_n4 ), 
        .B(\Red_MCInst_MC1_v3_2Inst_0_n3 ), .ZN(\Red_MCInst_MC1_v3_2 [0]) );
  XNOR2_X1 \Red_MCInst_MC1_v3_2Inst_0_U4  ( .A(\Red_MCInst_MC1_v3_3 [2]), .B(
        \MCInst_MC1_v3_2 [3]), .ZN(\Red_MCInst_MC1_v3_2Inst_0_n3 ) );
  XOR2_X1 \Red_MCInst_MC1_v3_2Inst_0_U3  ( .A(\MCInst_MC1_v3_0 [3]), .B(
        \Red_MCInst_MC1_v3_1 [2]), .Z(\Red_MCInst_MC1_v3_2Inst_0_n4 ) );
  XOR2_X1 \Red_MCInst_MC1_v3_3Inst_0_U3  ( .A(\MCInst_MC1_v3_0 [3]), .B(
        \Red_MCInst_MC1_v3_1 [2]), .Z(\Red_MCInst_MC1_v3_3 [0]) );
  XOR2_X1 \Red_MCInst_MC1_v0_0Inst_1_U3  ( .A(\Red_MCInst_MC1_v0_2 [2]), .B(
        \Red_MCInst_MC1_v0_1 [0]), .Z(\Red_MCInst_MC1_v0_0 [1]) );
  XNOR2_X1 \Red_MCInst_MC1_v0_1Inst_1_U4  ( .A(\Red_MCInst_MC1_v0_1Inst_1_n2 ), 
        .B(\MCInst_MC1_v0_3 [3]), .ZN(\Red_MCInst_MC1_v0_1 [1]) );
  XNOR2_X1 \Red_MCInst_MC1_v0_1Inst_1_U3  ( .A(\Red_MCInst_MC1_v0_1 [0]), .B(
        \Red_MCInst_MC1_v0_0 [0]), .ZN(\Red_MCInst_MC1_v0_1Inst_1_n2 ) );
  XOR2_X1 \Red_MCInst_MC1_v0_2Inst_1_U3  ( .A(\Red_MCInst_MC1_v0_0 [0]), .B(
        \Red_MCInst_MC1_v0_2 [2]), .Z(\Red_MCInst_MC1_v0_2 [1]) );
  XOR2_X1 \Red_MCInst_MC1_v0_3Inst_1_U3  ( .A(\Red_MCInst_MC1_v0_0 [0]), .B(
        \MCInst_MC1_v0_3 [3]), .Z(\Red_MCInst_MC1_v0_3 [1]) );
  XNOR2_X1 \Red_MCInst_MC1_v1_0Inst_1_U4  ( .A(\Red_MCInst_MC1_v1_0Inst_1_n2 ), 
        .B(\Red_MCInst_MC1_v1_2 [1]), .ZN(\Red_MCInst_MC1_v1_0 [1]) );
  XNOR2_X1 \Red_MCInst_MC1_v1_0Inst_1_U3  ( .A(\Red_MCInst_MC1_v1_1 [2]), .B(
        \MCInst_MC1_v1_0 [0]), .ZN(\Red_MCInst_MC1_v1_0Inst_1_n2 ) );
  XNOR2_X1 \Red_MCInst_MC1_v1_1Inst_1_U5  ( .A(\Red_MCInst_MC1_v1_1Inst_1_n4 ), 
        .B(\Red_MCInst_MC1_v1_1Inst_1_n3 ), .ZN(\Red_MCInst_MC1_v1_1 [1]) );
  XNOR2_X1 \Red_MCInst_MC1_v1_1Inst_1_U4  ( .A(\Red_MCInst_MC1_v1_2 [1]), .B(
        \MCInst_MC1_v1_0 [0]), .ZN(\Red_MCInst_MC1_v1_1Inst_1_n3 ) );
  XOR2_X1 \Red_MCInst_MC1_v1_1Inst_1_U3  ( .A(\MCInst_MC1_v1_3 [3]), .B(
        \Red_MCInst_MC1_v1_1 [2]), .Z(\Red_MCInst_MC1_v1_1Inst_1_n4 ) );
  XOR2_X1 \Red_MCInst_MC1_v1_3Inst_1_U3  ( .A(\MCInst_MC1_v1_0 [0]), .B(
        \MCInst_MC1_v1_3 [3]), .Z(\Red_MCInst_MC1_v1_3 [1]) );
  XOR2_X1 \Red_MCInst_MC1_v2_0Inst_1_U3  ( .A(\Red_MCInst_MC1_v2_1 [1]), .B(
        \MCInst_MC1_v2_0 [3]), .Z(\Red_MCInst_MC1_v2_0 [1]) );
  XOR2_X1 \Red_MCInst_MC1_v2_3Inst_1_U3  ( .A(\Red_MCInst_MC1_v2_1 [1]), .B(
        \Red_MCInst_MC1_v2_2 [1]), .Z(\Red_MCInst_MC1_v2_3 [1]) );
  XOR2_X1 \Red_MCInst_MC1_v3_0Inst_1_U3  ( .A(\MCInst_MC1_v3_2 [3]), .B(
        \MCInst_MC1_v3_0 [3]), .Z(\Red_MCInst_MC1_v3_0 [1]) );
  XNOR2_X1 \Red_MCInst_MC1_v3_1Inst_1_U5  ( .A(\Red_MCInst_MC1_v3_1Inst_1_n4 ), 
        .B(\Red_MCInst_MC1_v3_1Inst_1_n3 ), .ZN(\Red_MCInst_MC1_v3_1 [1]) );
  XNOR2_X1 \Red_MCInst_MC1_v3_1Inst_1_U4  ( .A(\Red_MCInst_MC1_v3_3 [2]), .B(
        \MCInst_MC1_v3_2 [3]), .ZN(\Red_MCInst_MC1_v3_1Inst_1_n3 ) );
  XOR2_X1 \Red_MCInst_MC1_v3_1Inst_1_U3  ( .A(\MCInst_MC1_v3_0 [3]), .B(
        \Red_MCInst_MC1_v3_1 [2]), .Z(\Red_MCInst_MC1_v3_1Inst_1_n4 ) );
  XOR2_X1 \Red_MCInst_MC1_v3_2Inst_1_U3  ( .A(\Red_MCInst_MC1_v3_3 [2]), .B(
        \MCInst_MC1_v3_0 [3]), .Z(\Red_MCInst_MC1_v3_2 [1]) );
  XOR2_X1 \Red_MCInst_MC1_v3_3Inst_1_U3  ( .A(\MCInst_MC1_v3_2 [3]), .B(
        \Red_MCInst_MC1_v3_3 [2]), .Z(\Red_MCInst_MC1_v3_3 [1]) );
  XNOR2_X1 \Red_MCInst_MC1_v0_0Inst_2_U4  ( .A(\Red_MCInst_MC1_v0_0Inst_2_n2 ), 
        .B(\Red_MCInst_MC1_v0_2 [2]), .ZN(\Red_MCInst_MC1_v0_0 [2]) );
  XNOR2_X1 \Red_MCInst_MC1_v0_0Inst_2_U3  ( .A(\MCInst_MC1_v0_3 [3]), .B(
        \Red_MCInst_MC1_v0_0 [0]), .ZN(\Red_MCInst_MC1_v0_0Inst_2_n2 ) );
  XOR2_X1 \Red_MCInst_MC1_v0_1Inst_2_U3  ( .A(\Red_MCInst_MC1_v0_0 [0]), .B(
        \Red_MCInst_MC1_v0_2 [2]), .Z(\Red_MCInst_MC1_v0_1 [2]) );
  XNOR2_X1 \Red_MCInst_MC1_v0_3Inst_2_U5  ( .A(\Red_MCInst_MC1_v0_3Inst_2_n4 ), 
        .B(\Red_MCInst_MC1_v0_3Inst_2_n3 ), .ZN(\Red_MCInst_MC1_v0_3 [2]) );
  XNOR2_X1 \Red_MCInst_MC1_v0_3Inst_2_U4  ( .A(\Red_MCInst_MC1_v0_2 [2]), .B(
        \Red_MCInst_MC1_v0_0 [0]), .ZN(\Red_MCInst_MC1_v0_3Inst_2_n3 ) );
  XOR2_X1 \Red_MCInst_MC1_v0_3Inst_2_U3  ( .A(\MCInst_MC1_v0_3 [3]), .B(
        \Red_MCInst_MC1_v0_1 [0]), .Z(\Red_MCInst_MC1_v0_3Inst_2_n4 ) );
  XNOR2_X1 \Red_MCInst_MC1_v1_0Inst_2_U4  ( .A(\Red_MCInst_MC1_v1_0Inst_2_n2 ), 
        .B(\MCInst_MC1_v1_3 [3]), .ZN(\Red_MCInst_MC1_v1_0 [2]) );
  XNOR2_X1 \Red_MCInst_MC1_v1_0Inst_2_U3  ( .A(\Red_MCInst_MC1_v1_1 [2]), .B(
        \Red_MCInst_MC1_v1_2 [1]), .ZN(\Red_MCInst_MC1_v1_0Inst_2_n2 ) );
  XNOR2_X1 \Red_MCInst_MC1_v1_2Inst_2_U4  ( .A(\Red_MCInst_MC1_v1_2Inst_2_n2 ), 
        .B(\Red_MCInst_MC1_v1_2 [1]), .ZN(\Red_MCInst_MC1_v1_2 [2]) );
  XNOR2_X1 \Red_MCInst_MC1_v1_2Inst_2_U3  ( .A(\Red_MCInst_MC1_v1_1 [2]), .B(
        \MCInst_MC1_v1_0 [0]), .ZN(\Red_MCInst_MC1_v1_2Inst_2_n2 ) );
  XNOR2_X1 \Red_MCInst_MC1_v1_3Inst_2_U5  ( .A(\Red_MCInst_MC1_v1_3Inst_2_n4 ), 
        .B(\Red_MCInst_MC1_v1_3Inst_2_n3 ), .ZN(\Red_MCInst_MC1_v1_3 [2]) );
  XNOR2_X1 \Red_MCInst_MC1_v1_3Inst_2_U4  ( .A(\Red_MCInst_MC1_v1_2 [1]), .B(
        \MCInst_MC1_v1_0 [0]), .ZN(\Red_MCInst_MC1_v1_3Inst_2_n3 ) );
  XOR2_X1 \Red_MCInst_MC1_v1_3Inst_2_U3  ( .A(\MCInst_MC1_v1_3 [3]), .B(
        \Red_MCInst_MC1_v1_1 [2]), .Z(\Red_MCInst_MC1_v1_3Inst_2_n4 ) );
  XNOR2_X1 \Red_MCInst_MC1_v2_0Inst_2_U5  ( .A(\Red_MCInst_MC1_v2_0Inst_2_n4 ), 
        .B(\Red_MCInst_MC1_v2_0Inst_2_n3 ), .ZN(\Red_MCInst_MC1_v2_0 [2]) );
  XNOR2_X1 \Red_MCInst_MC1_v2_0Inst_2_U4  ( .A(\MCInst_MC1_v2_0 [2]), .B(
        \Red_MCInst_MC1_v2_1 [1]), .ZN(\Red_MCInst_MC1_v2_0Inst_2_n3 ) );
  XOR2_X1 \Red_MCInst_MC1_v2_0Inst_2_U3  ( .A(\MCInst_MC1_v2_0 [3]), .B(
        \Red_MCInst_MC1_v2_2 [1]), .Z(\Red_MCInst_MC1_v2_0Inst_2_n4 ) );
  XOR2_X1 \Red_MCInst_MC1_v2_1Inst_2_U3  ( .A(\Red_MCInst_MC1_v2_1 [1]), .B(
        \Red_MCInst_MC1_v2_2 [1]), .Z(\Red_MCInst_MC1_v2_1 [2]) );
  XOR2_X1 \Red_MCInst_MC1_v2_2Inst_2_U3  ( .A(\MCInst_MC1_v2_0 [3]), .B(
        \Red_MCInst_MC1_v2_2 [1]), .Z(\Red_MCInst_MC1_v2_2 [2]) );
  XOR2_X1 \Red_MCInst_MC1_v2_3Inst_2_U3  ( .A(\Red_MCInst_MC1_v2_1 [1]), .B(
        \MCInst_MC1_v2_0 [3]), .Z(\Red_MCInst_MC1_v2_3 [2]) );
  XNOR2_X1 \Red_MCInst_MC1_v3_0Inst_2_U5  ( .A(\Red_MCInst_MC1_v3_0Inst_2_n4 ), 
        .B(\Red_MCInst_MC1_v3_0Inst_2_n3 ), .ZN(\Red_MCInst_MC1_v3_0 [2]) );
  XNOR2_X1 \Red_MCInst_MC1_v3_0Inst_2_U4  ( .A(\Red_MCInst_MC1_v3_3 [2]), .B(
        \MCInst_MC1_v3_2 [3]), .ZN(\Red_MCInst_MC1_v3_0Inst_2_n3 ) );
  XOR2_X1 \Red_MCInst_MC1_v3_0Inst_2_U3  ( .A(\MCInst_MC1_v3_0 [3]), .B(
        \Red_MCInst_MC1_v3_1 [2]), .Z(\Red_MCInst_MC1_v3_0Inst_2_n4 ) );
  XNOR2_X1 \Red_MCInst_MC1_v3_2Inst_2_U4  ( .A(\Red_MCInst_MC1_v3_2Inst_2_n2 ), 
        .B(\MCInst_MC1_v3_0 [3]), .ZN(\Red_MCInst_MC1_v3_2 [2]) );
  XNOR2_X1 \Red_MCInst_MC1_v3_2Inst_2_U3  ( .A(\Red_MCInst_MC1_v3_1 [2]), .B(
        \MCInst_MC1_v3_2 [3]), .ZN(\Red_MCInst_MC1_v3_2Inst_2_n2 ) );
  XNOR2_X1 \Red_MCInst_MC1_r0Inst_XORInst_0_0_U3  ( .A(
        \Red_MCInst_MC1_r0Inst_XORInst_0_0_n5 ), .B(
        \Red_MCInst_MC1_r0Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback[42]) );
  XNOR2_X1 \Red_MCInst_MC1_r0Inst_XORInst_0_0_U2  ( .A(
        \Red_MCInst_MC1_v3_0 [0]), .B(\Red_MCInst_MC1_v2_0 [0]), .ZN(
        \Red_MCInst_MC1_r0Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \Red_MCInst_MC1_r0Inst_XORInst_0_0_U1  ( .A(\Red_MCInst_MC1_v0_0 [0]), .B(\Red_MCInst_MC1_v1_0 [0]), .Z(\Red_MCInst_MC1_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \Red_MCInst_MC1_r0Inst_XORInst_0_1_U3  ( .A(
        \Red_MCInst_MC1_r0Inst_XORInst_0_1_n5 ), .B(
        \Red_MCInst_MC1_r0Inst_XORInst_0_1_n4 ), .ZN(Red_Feedback[43]) );
  XNOR2_X1 \Red_MCInst_MC1_r0Inst_XORInst_0_1_U2  ( .A(
        \Red_MCInst_MC1_v3_0 [1]), .B(\Red_MCInst_MC1_v2_0 [1]), .ZN(
        \Red_MCInst_MC1_r0Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \Red_MCInst_MC1_r0Inst_XORInst_0_1_U1  ( .A(\Red_MCInst_MC1_v0_0 [1]), .B(\Red_MCInst_MC1_v1_0 [1]), .Z(\Red_MCInst_MC1_r0Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \Red_MCInst_MC1_r0Inst_XORInst_0_2_U3  ( .A(
        \Red_MCInst_MC1_r0Inst_XORInst_0_2_n5 ), .B(
        \Red_MCInst_MC1_r0Inst_XORInst_0_2_n4 ), .ZN(Red_Feedback[44]) );
  XNOR2_X1 \Red_MCInst_MC1_r0Inst_XORInst_0_2_U2  ( .A(
        \Red_MCInst_MC1_v3_0 [2]), .B(\Red_MCInst_MC1_v2_0 [2]), .ZN(
        \Red_MCInst_MC1_r0Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \Red_MCInst_MC1_r0Inst_XORInst_0_2_U1  ( .A(\Red_MCInst_MC1_v0_0 [2]), .B(\Red_MCInst_MC1_v1_0 [2]), .Z(\Red_MCInst_MC1_r0Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \Red_MCInst_MC1_r1Inst_XORInst_0_0_U3  ( .A(
        \Red_MCInst_MC1_r1Inst_XORInst_0_0_n5 ), .B(
        \Red_MCInst_MC1_r1Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback[30]) );
  XNOR2_X1 \Red_MCInst_MC1_r1Inst_XORInst_0_0_U2  ( .A(
        \Red_MCInst_MC1_v3_3 [2]), .B(\Red_MCInst_MC1_v2_1 [0]), .ZN(
        \Red_MCInst_MC1_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \Red_MCInst_MC1_r1Inst_XORInst_0_0_U1  ( .A(\Red_MCInst_MC1_v0_1 [0]), .B(\Red_MCInst_MC1_v1_2 [1]), .Z(\Red_MCInst_MC1_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \Red_MCInst_MC1_r1Inst_XORInst_0_1_U3  ( .A(
        \Red_MCInst_MC1_r1Inst_XORInst_0_1_n5 ), .B(
        \Red_MCInst_MC1_r1Inst_XORInst_0_1_n4 ), .ZN(Red_Feedback[31]) );
  XNOR2_X1 \Red_MCInst_MC1_r1Inst_XORInst_0_1_U2  ( .A(
        \Red_MCInst_MC1_v3_1 [1]), .B(\Red_MCInst_MC1_v2_1 [1]), .ZN(
        \Red_MCInst_MC1_r1Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \Red_MCInst_MC1_r1Inst_XORInst_0_1_U1  ( .A(\Red_MCInst_MC1_v0_1 [1]), .B(\Red_MCInst_MC1_v1_1 [1]), .Z(\Red_MCInst_MC1_r1Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \Red_MCInst_MC1_r1Inst_XORInst_0_2_U3  ( .A(
        \Red_MCInst_MC1_r1Inst_XORInst_0_2_n5 ), .B(
        \Red_MCInst_MC1_r1Inst_XORInst_0_2_n4 ), .ZN(Red_Feedback[32]) );
  XNOR2_X1 \Red_MCInst_MC1_r1Inst_XORInst_0_2_U2  ( .A(
        \Red_MCInst_MC1_v3_1 [2]), .B(\Red_MCInst_MC1_v2_1 [2]), .ZN(
        \Red_MCInst_MC1_r1Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \Red_MCInst_MC1_r1Inst_XORInst_0_2_U1  ( .A(\Red_MCInst_MC1_v0_1 [2]), .B(\Red_MCInst_MC1_v1_1 [2]), .Z(\Red_MCInst_MC1_r1Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \Red_MCInst_MC1_r2Inst_XORInst_0_0_U3  ( .A(
        \Red_MCInst_MC1_r2Inst_XORInst_0_0_n5 ), .B(
        \Red_MCInst_MC1_r2Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback[18]) );
  XNOR2_X1 \Red_MCInst_MC1_r2Inst_XORInst_0_0_U2  ( .A(
        \Red_MCInst_MC1_v3_2 [0]), .B(\Red_MCInst_MC1_v2_2 [0]), .ZN(
        \Red_MCInst_MC1_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \Red_MCInst_MC1_r2Inst_XORInst_0_0_U1  ( .A(\Red_MCInst_MC1_v0_2 [0]), .B(\Red_MCInst_MC1_v1_2 [0]), .Z(\Red_MCInst_MC1_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \Red_MCInst_MC1_r2Inst_XORInst_0_1_U3  ( .A(
        \Red_MCInst_MC1_r2Inst_XORInst_0_1_n5 ), .B(
        \Red_MCInst_MC1_r2Inst_XORInst_0_1_n4 ), .ZN(Red_Feedback[19]) );
  XNOR2_X1 \Red_MCInst_MC1_r2Inst_XORInst_0_1_U2  ( .A(
        \Red_MCInst_MC1_v3_2 [1]), .B(\Red_MCInst_MC1_v2_2 [1]), .ZN(
        \Red_MCInst_MC1_r2Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \Red_MCInst_MC1_r2Inst_XORInst_0_1_U1  ( .A(\Red_MCInst_MC1_v0_2 [1]), .B(\Red_MCInst_MC1_v1_2 [1]), .Z(\Red_MCInst_MC1_r2Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \Red_MCInst_MC1_r2Inst_XORInst_0_2_U3  ( .A(
        \Red_MCInst_MC1_r2Inst_XORInst_0_2_n5 ), .B(
        \Red_MCInst_MC1_r2Inst_XORInst_0_2_n4 ), .ZN(Red_Feedback[20]) );
  XNOR2_X1 \Red_MCInst_MC1_r2Inst_XORInst_0_2_U2  ( .A(
        \Red_MCInst_MC1_v3_2 [2]), .B(\Red_MCInst_MC1_v2_2 [2]), .ZN(
        \Red_MCInst_MC1_r2Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \Red_MCInst_MC1_r2Inst_XORInst_0_2_U1  ( .A(\Red_MCInst_MC1_v0_2 [2]), .B(\Red_MCInst_MC1_v1_2 [2]), .Z(\Red_MCInst_MC1_r2Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \Red_MCInst_MC1_r3Inst_XORInst_0_0_U3  ( .A(
        \Red_MCInst_MC1_r3Inst_XORInst_0_0_n5 ), .B(
        \Red_MCInst_MC1_r3Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback[6]) );
  XNOR2_X1 \Red_MCInst_MC1_r3Inst_XORInst_0_0_U2  ( .A(
        \Red_MCInst_MC1_v3_3 [0]), .B(\Red_MCInst_MC1_v2_3 [0]), .ZN(
        \Red_MCInst_MC1_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \Red_MCInst_MC1_r3Inst_XORInst_0_0_U1  ( .A(\Red_MCInst_MC1_v0_3 [0]), .B(\Red_MCInst_MC1_v1_3 [0]), .Z(\Red_MCInst_MC1_r3Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \Red_MCInst_MC1_r3Inst_XORInst_0_1_U3  ( .A(
        \Red_MCInst_MC1_r3Inst_XORInst_0_1_n5 ), .B(
        \Red_MCInst_MC1_r3Inst_XORInst_0_1_n4 ), .ZN(Red_Feedback[7]) );
  XNOR2_X1 \Red_MCInst_MC1_r3Inst_XORInst_0_1_U2  ( .A(
        \Red_MCInst_MC1_v3_3 [1]), .B(\Red_MCInst_MC1_v2_3 [1]), .ZN(
        \Red_MCInst_MC1_r3Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \Red_MCInst_MC1_r3Inst_XORInst_0_1_U1  ( .A(\Red_MCInst_MC1_v0_3 [1]), .B(\Red_MCInst_MC1_v1_3 [1]), .Z(\Red_MCInst_MC1_r3Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \Red_MCInst_MC1_r3Inst_XORInst_0_2_U3  ( .A(
        \Red_MCInst_MC1_r3Inst_XORInst_0_2_n5 ), .B(
        \Red_MCInst_MC1_r3Inst_XORInst_0_2_n4 ), .ZN(Red_Feedback[8]) );
  XNOR2_X1 \Red_MCInst_MC1_r3Inst_XORInst_0_2_U2  ( .A(
        \Red_MCInst_MC1_v3_3 [2]), .B(\Red_MCInst_MC1_v2_3 [2]), .ZN(
        \Red_MCInst_MC1_r3Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \Red_MCInst_MC1_r3Inst_XORInst_0_2_U1  ( .A(\Red_MCInst_MC1_v0_3 [2]), .B(\Red_MCInst_MC1_v1_3 [2]), .Z(\Red_MCInst_MC1_r3Inst_XORInst_0_2_n5 ) );
  XOR2_X1 \Red_MCInst_MC2_v0_2Inst_0_U3  ( .A(\MCInst_MC2_v0_3 [3]), .B(
        \Red_MCInst_MC2_v0_1 [0]), .Z(\Red_MCInst_MC2_v0_2 [0]) );
  XOR2_X1 \Red_MCInst_MC2_v0_3Inst_0_U3  ( .A(\Red_MCInst_MC2_v0_0 [0]), .B(
        \Red_MCInst_MC2_v0_2 [2]), .Z(\Red_MCInst_MC2_v0_3 [0]) );
  XNOR2_X1 \Red_MCInst_MC2_v1_0Inst_0_U4  ( .A(\Red_MCInst_MC2_v1_0Inst_0_n2 ), 
        .B(\Red_MCInst_MC2_v1_2 [1]), .ZN(\Red_MCInst_MC2_v1_0 [0]) );
  XNOR2_X1 \Red_MCInst_MC2_v1_0Inst_0_U3  ( .A(\MCInst_MC2_v1_3 [3]), .B(
        \MCInst_MC2_v1_0 [0]), .ZN(\Red_MCInst_MC2_v1_0Inst_0_n2 ) );
  XOR2_X1 \Red_MCInst_MC2_v1_2Inst_0_U3  ( .A(\Red_MCInst_MC2_v1_2 [1]), .B(
        \Red_MCInst_MC2_v1_1 [2]), .Z(\Red_MCInst_MC2_v1_2 [0]) );
  XOR2_X1 \Red_MCInst_MC2_v1_3Inst_0_U3  ( .A(\MCInst_MC2_v1_0 [0]), .B(
        \Red_MCInst_MC2_v1_2 [1]), .Z(\Red_MCInst_MC2_v1_3 [0]) );
  XOR2_X1 \Red_MCInst_MC2_v2_0Inst_0_U3  ( .A(\Red_MCInst_MC2_v2_1 [1]), .B(
        \MCInst_MC2_v2_0 [2]), .Z(\Red_MCInst_MC2_v2_0 [0]) );
  XOR2_X1 \Red_MCInst_MC2_v2_1Inst_0_U3  ( .A(\MCInst_MC2_v2_0 [2]), .B(
        \MCInst_MC2_v2_0 [3]), .Z(\Red_MCInst_MC2_v2_1 [0]) );
  XNOR2_X1 \Red_MCInst_MC2_v2_2Inst_0_U4  ( .A(\Red_MCInst_MC2_v2_2Inst_0_n2 ), 
        .B(\MCInst_MC2_v2_0 [2]), .ZN(\Red_MCInst_MC2_v2_2 [0]) );
  XNOR2_X1 \Red_MCInst_MC2_v2_2Inst_0_U3  ( .A(\Red_MCInst_MC2_v2_2 [1]), .B(
        \Red_MCInst_MC2_v2_1 [1]), .ZN(\Red_MCInst_MC2_v2_2Inst_0_n2 ) );
  XNOR2_X1 \Red_MCInst_MC2_v2_3Inst_0_U4  ( .A(\Red_MCInst_MC2_v2_3Inst_0_n2 ), 
        .B(\MCInst_MC2_v2_0 [3]), .ZN(\Red_MCInst_MC2_v2_3 [0]) );
  XNOR2_X1 \Red_MCInst_MC2_v2_3Inst_0_U3  ( .A(\Red_MCInst_MC2_v2_2 [1]), .B(
        \Red_MCInst_MC2_v2_1 [1]), .ZN(\Red_MCInst_MC2_v2_3Inst_0_n2 ) );
  XOR2_X1 \Red_MCInst_MC2_v3_0Inst_0_U3  ( .A(\MCInst_MC2_v3_2 [3]), .B(
        \Red_MCInst_MC2_v3_3 [2]), .Z(\Red_MCInst_MC2_v3_0 [0]) );
  XNOR2_X1 \Red_MCInst_MC2_v3_2Inst_0_U5  ( .A(\Red_MCInst_MC2_v3_2Inst_0_n4 ), 
        .B(\Red_MCInst_MC2_v3_2Inst_0_n3 ), .ZN(\Red_MCInst_MC2_v3_2 [0]) );
  XNOR2_X1 \Red_MCInst_MC2_v3_2Inst_0_U4  ( .A(\Red_MCInst_MC2_v3_3 [2]), .B(
        \MCInst_MC2_v3_2 [3]), .ZN(\Red_MCInst_MC2_v3_2Inst_0_n3 ) );
  XOR2_X1 \Red_MCInst_MC2_v3_2Inst_0_U3  ( .A(\MCInst_MC2_v3_0 [3]), .B(
        \Red_MCInst_MC2_v3_1 [2]), .Z(\Red_MCInst_MC2_v3_2Inst_0_n4 ) );
  XOR2_X1 \Red_MCInst_MC2_v3_3Inst_0_U3  ( .A(\MCInst_MC2_v3_0 [3]), .B(
        \Red_MCInst_MC2_v3_1 [2]), .Z(\Red_MCInst_MC2_v3_3 [0]) );
  XOR2_X1 \Red_MCInst_MC2_v0_0Inst_1_U3  ( .A(\Red_MCInst_MC2_v0_2 [2]), .B(
        \Red_MCInst_MC2_v0_1 [0]), .Z(\Red_MCInst_MC2_v0_0 [1]) );
  XNOR2_X1 \Red_MCInst_MC2_v0_1Inst_1_U4  ( .A(\Red_MCInst_MC2_v0_1Inst_1_n2 ), 
        .B(\MCInst_MC2_v0_3 [3]), .ZN(\Red_MCInst_MC2_v0_1 [1]) );
  XNOR2_X1 \Red_MCInst_MC2_v0_1Inst_1_U3  ( .A(\Red_MCInst_MC2_v0_1 [0]), .B(
        \Red_MCInst_MC2_v0_0 [0]), .ZN(\Red_MCInst_MC2_v0_1Inst_1_n2 ) );
  XOR2_X1 \Red_MCInst_MC2_v0_2Inst_1_U3  ( .A(\Red_MCInst_MC2_v0_0 [0]), .B(
        \Red_MCInst_MC2_v0_2 [2]), .Z(\Red_MCInst_MC2_v0_2 [1]) );
  XOR2_X1 \Red_MCInst_MC2_v0_3Inst_1_U3  ( .A(\Red_MCInst_MC2_v0_0 [0]), .B(
        \MCInst_MC2_v0_3 [3]), .Z(\Red_MCInst_MC2_v0_3 [1]) );
  XNOR2_X1 \Red_MCInst_MC2_v1_0Inst_1_U4  ( .A(\Red_MCInst_MC2_v1_0Inst_1_n2 ), 
        .B(\Red_MCInst_MC2_v1_2 [1]), .ZN(\Red_MCInst_MC2_v1_0 [1]) );
  XNOR2_X1 \Red_MCInst_MC2_v1_0Inst_1_U3  ( .A(\Red_MCInst_MC2_v1_1 [2]), .B(
        \MCInst_MC2_v1_0 [0]), .ZN(\Red_MCInst_MC2_v1_0Inst_1_n2 ) );
  XNOR2_X1 \Red_MCInst_MC2_v1_1Inst_1_U5  ( .A(\Red_MCInst_MC2_v1_1Inst_1_n4 ), 
        .B(\Red_MCInst_MC2_v1_1Inst_1_n3 ), .ZN(\Red_MCInst_MC2_v1_1 [1]) );
  XNOR2_X1 \Red_MCInst_MC2_v1_1Inst_1_U4  ( .A(\Red_MCInst_MC2_v1_2 [1]), .B(
        \MCInst_MC2_v1_0 [0]), .ZN(\Red_MCInst_MC2_v1_1Inst_1_n3 ) );
  XOR2_X1 \Red_MCInst_MC2_v1_1Inst_1_U3  ( .A(\MCInst_MC2_v1_3 [3]), .B(
        \Red_MCInst_MC2_v1_1 [2]), .Z(\Red_MCInst_MC2_v1_1Inst_1_n4 ) );
  XOR2_X1 \Red_MCInst_MC2_v1_3Inst_1_U3  ( .A(\MCInst_MC2_v1_0 [0]), .B(
        \MCInst_MC2_v1_3 [3]), .Z(\Red_MCInst_MC2_v1_3 [1]) );
  XOR2_X1 \Red_MCInst_MC2_v2_0Inst_1_U3  ( .A(\Red_MCInst_MC2_v2_1 [1]), .B(
        \MCInst_MC2_v2_0 [3]), .Z(\Red_MCInst_MC2_v2_0 [1]) );
  XOR2_X1 \Red_MCInst_MC2_v2_3Inst_1_U3  ( .A(\Red_MCInst_MC2_v2_1 [1]), .B(
        \Red_MCInst_MC2_v2_2 [1]), .Z(\Red_MCInst_MC2_v2_3 [1]) );
  XOR2_X1 \Red_MCInst_MC2_v3_0Inst_1_U3  ( .A(\MCInst_MC2_v3_2 [3]), .B(
        \MCInst_MC2_v3_0 [3]), .Z(\Red_MCInst_MC2_v3_0 [1]) );
  XNOR2_X1 \Red_MCInst_MC2_v3_1Inst_1_U5  ( .A(\Red_MCInst_MC2_v3_1Inst_1_n4 ), 
        .B(\Red_MCInst_MC2_v3_1Inst_1_n3 ), .ZN(\Red_MCInst_MC2_v3_1 [1]) );
  XNOR2_X1 \Red_MCInst_MC2_v3_1Inst_1_U4  ( .A(\Red_MCInst_MC2_v3_3 [2]), .B(
        \MCInst_MC2_v3_2 [3]), .ZN(\Red_MCInst_MC2_v3_1Inst_1_n3 ) );
  XOR2_X1 \Red_MCInst_MC2_v3_1Inst_1_U3  ( .A(\MCInst_MC2_v3_0 [3]), .B(
        \Red_MCInst_MC2_v3_1 [2]), .Z(\Red_MCInst_MC2_v3_1Inst_1_n4 ) );
  XOR2_X1 \Red_MCInst_MC2_v3_2Inst_1_U3  ( .A(\Red_MCInst_MC2_v3_3 [2]), .B(
        \MCInst_MC2_v3_0 [3]), .Z(\Red_MCInst_MC2_v3_2 [1]) );
  XOR2_X1 \Red_MCInst_MC2_v3_3Inst_1_U3  ( .A(\MCInst_MC2_v3_2 [3]), .B(
        \Red_MCInst_MC2_v3_3 [2]), .Z(\Red_MCInst_MC2_v3_3 [1]) );
  XNOR2_X1 \Red_MCInst_MC2_v0_0Inst_2_U4  ( .A(\Red_MCInst_MC2_v0_0Inst_2_n2 ), 
        .B(\Red_MCInst_MC2_v0_2 [2]), .ZN(\Red_MCInst_MC2_v0_0 [2]) );
  XNOR2_X1 \Red_MCInst_MC2_v0_0Inst_2_U3  ( .A(\MCInst_MC2_v0_3 [3]), .B(
        \Red_MCInst_MC2_v0_0 [0]), .ZN(\Red_MCInst_MC2_v0_0Inst_2_n2 ) );
  XOR2_X1 \Red_MCInst_MC2_v0_1Inst_2_U3  ( .A(\Red_MCInst_MC2_v0_0 [0]), .B(
        \Red_MCInst_MC2_v0_2 [2]), .Z(\Red_MCInst_MC2_v0_1 [2]) );
  XNOR2_X1 \Red_MCInst_MC2_v0_3Inst_2_U5  ( .A(\Red_MCInst_MC2_v0_3Inst_2_n4 ), 
        .B(\Red_MCInst_MC2_v0_3Inst_2_n3 ), .ZN(\Red_MCInst_MC2_v0_3 [2]) );
  XNOR2_X1 \Red_MCInst_MC2_v0_3Inst_2_U4  ( .A(\Red_MCInst_MC2_v0_2 [2]), .B(
        \Red_MCInst_MC2_v0_0 [0]), .ZN(\Red_MCInst_MC2_v0_3Inst_2_n3 ) );
  XOR2_X1 \Red_MCInst_MC2_v0_3Inst_2_U3  ( .A(\MCInst_MC2_v0_3 [3]), .B(
        \Red_MCInst_MC2_v0_1 [0]), .Z(\Red_MCInst_MC2_v0_3Inst_2_n4 ) );
  XNOR2_X1 \Red_MCInst_MC2_v1_0Inst_2_U4  ( .A(\Red_MCInst_MC2_v1_0Inst_2_n2 ), 
        .B(\MCInst_MC2_v1_3 [3]), .ZN(\Red_MCInst_MC2_v1_0 [2]) );
  XNOR2_X1 \Red_MCInst_MC2_v1_0Inst_2_U3  ( .A(\Red_MCInst_MC2_v1_1 [2]), .B(
        \Red_MCInst_MC2_v1_2 [1]), .ZN(\Red_MCInst_MC2_v1_0Inst_2_n2 ) );
  XNOR2_X1 \Red_MCInst_MC2_v1_2Inst_2_U4  ( .A(\Red_MCInst_MC2_v1_2Inst_2_n2 ), 
        .B(\Red_MCInst_MC2_v1_2 [1]), .ZN(\Red_MCInst_MC2_v1_2 [2]) );
  XNOR2_X1 \Red_MCInst_MC2_v1_2Inst_2_U3  ( .A(\Red_MCInst_MC2_v1_1 [2]), .B(
        \MCInst_MC2_v1_0 [0]), .ZN(\Red_MCInst_MC2_v1_2Inst_2_n2 ) );
  XNOR2_X1 \Red_MCInst_MC2_v1_3Inst_2_U5  ( .A(\Red_MCInst_MC2_v1_3Inst_2_n4 ), 
        .B(\Red_MCInst_MC2_v1_3Inst_2_n3 ), .ZN(\Red_MCInst_MC2_v1_3 [2]) );
  XNOR2_X1 \Red_MCInst_MC2_v1_3Inst_2_U4  ( .A(\Red_MCInst_MC2_v1_2 [1]), .B(
        \MCInst_MC2_v1_0 [0]), .ZN(\Red_MCInst_MC2_v1_3Inst_2_n3 ) );
  XOR2_X1 \Red_MCInst_MC2_v1_3Inst_2_U3  ( .A(\MCInst_MC2_v1_3 [3]), .B(
        \Red_MCInst_MC2_v1_1 [2]), .Z(\Red_MCInst_MC2_v1_3Inst_2_n4 ) );
  XNOR2_X1 \Red_MCInst_MC2_v2_0Inst_2_U5  ( .A(\Red_MCInst_MC2_v2_0Inst_2_n4 ), 
        .B(\Red_MCInst_MC2_v2_0Inst_2_n3 ), .ZN(\Red_MCInst_MC2_v2_0 [2]) );
  XNOR2_X1 \Red_MCInst_MC2_v2_0Inst_2_U4  ( .A(\MCInst_MC2_v2_0 [2]), .B(
        \Red_MCInst_MC2_v2_1 [1]), .ZN(\Red_MCInst_MC2_v2_0Inst_2_n3 ) );
  XOR2_X1 \Red_MCInst_MC2_v2_0Inst_2_U3  ( .A(\MCInst_MC2_v2_0 [3]), .B(
        \Red_MCInst_MC2_v2_2 [1]), .Z(\Red_MCInst_MC2_v2_0Inst_2_n4 ) );
  XOR2_X1 \Red_MCInst_MC2_v2_1Inst_2_U3  ( .A(\Red_MCInst_MC2_v2_1 [1]), .B(
        \Red_MCInst_MC2_v2_2 [1]), .Z(\Red_MCInst_MC2_v2_1 [2]) );
  XOR2_X1 \Red_MCInst_MC2_v2_2Inst_2_U3  ( .A(\MCInst_MC2_v2_0 [3]), .B(
        \Red_MCInst_MC2_v2_2 [1]), .Z(\Red_MCInst_MC2_v2_2 [2]) );
  XOR2_X1 \Red_MCInst_MC2_v2_3Inst_2_U3  ( .A(\Red_MCInst_MC2_v2_1 [1]), .B(
        \MCInst_MC2_v2_0 [3]), .Z(\Red_MCInst_MC2_v2_3 [2]) );
  XNOR2_X1 \Red_MCInst_MC2_v3_0Inst_2_U5  ( .A(\Red_MCInst_MC2_v3_0Inst_2_n4 ), 
        .B(\Red_MCInst_MC2_v3_0Inst_2_n3 ), .ZN(\Red_MCInst_MC2_v3_0 [2]) );
  XNOR2_X1 \Red_MCInst_MC2_v3_0Inst_2_U4  ( .A(\Red_MCInst_MC2_v3_3 [2]), .B(
        \MCInst_MC2_v3_2 [3]), .ZN(\Red_MCInst_MC2_v3_0Inst_2_n3 ) );
  XOR2_X1 \Red_MCInst_MC2_v3_0Inst_2_U3  ( .A(\MCInst_MC2_v3_0 [3]), .B(
        \Red_MCInst_MC2_v3_1 [2]), .Z(\Red_MCInst_MC2_v3_0Inst_2_n4 ) );
  XNOR2_X1 \Red_MCInst_MC2_v3_2Inst_2_U4  ( .A(\Red_MCInst_MC2_v3_2Inst_2_n2 ), 
        .B(\MCInst_MC2_v3_0 [3]), .ZN(\Red_MCInst_MC2_v3_2 [2]) );
  XNOR2_X1 \Red_MCInst_MC2_v3_2Inst_2_U3  ( .A(\Red_MCInst_MC2_v3_1 [2]), .B(
        \MCInst_MC2_v3_2 [3]), .ZN(\Red_MCInst_MC2_v3_2Inst_2_n2 ) );
  XNOR2_X1 \Red_MCInst_MC2_r0Inst_XORInst_0_0_U3  ( .A(
        \Red_MCInst_MC2_r0Inst_XORInst_0_0_n5 ), .B(
        \Red_MCInst_MC2_r0Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback[39]) );
  XNOR2_X1 \Red_MCInst_MC2_r0Inst_XORInst_0_0_U2  ( .A(
        \Red_MCInst_MC2_v3_0 [0]), .B(\Red_MCInst_MC2_v2_0 [0]), .ZN(
        \Red_MCInst_MC2_r0Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \Red_MCInst_MC2_r0Inst_XORInst_0_0_U1  ( .A(\Red_MCInst_MC2_v0_0 [0]), .B(\Red_MCInst_MC2_v1_0 [0]), .Z(\Red_MCInst_MC2_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \Red_MCInst_MC2_r0Inst_XORInst_0_1_U3  ( .A(
        \Red_MCInst_MC2_r0Inst_XORInst_0_1_n5 ), .B(
        \Red_MCInst_MC2_r0Inst_XORInst_0_1_n4 ), .ZN(Red_Feedback[40]) );
  XNOR2_X1 \Red_MCInst_MC2_r0Inst_XORInst_0_1_U2  ( .A(
        \Red_MCInst_MC2_v3_0 [1]), .B(\Red_MCInst_MC2_v2_0 [1]), .ZN(
        \Red_MCInst_MC2_r0Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \Red_MCInst_MC2_r0Inst_XORInst_0_1_U1  ( .A(\Red_MCInst_MC2_v0_0 [1]), .B(\Red_MCInst_MC2_v1_0 [1]), .Z(\Red_MCInst_MC2_r0Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \Red_MCInst_MC2_r0Inst_XORInst_0_2_U3  ( .A(
        \Red_MCInst_MC2_r0Inst_XORInst_0_2_n5 ), .B(
        \Red_MCInst_MC2_r0Inst_XORInst_0_2_n4 ), .ZN(Red_Feedback[41]) );
  XNOR2_X1 \Red_MCInst_MC2_r0Inst_XORInst_0_2_U2  ( .A(
        \Red_MCInst_MC2_v3_0 [2]), .B(\Red_MCInst_MC2_v2_0 [2]), .ZN(
        \Red_MCInst_MC2_r0Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \Red_MCInst_MC2_r0Inst_XORInst_0_2_U1  ( .A(\Red_MCInst_MC2_v0_0 [2]), .B(\Red_MCInst_MC2_v1_0 [2]), .Z(\Red_MCInst_MC2_r0Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \Red_MCInst_MC2_r1Inst_XORInst_0_0_U3  ( .A(
        \Red_MCInst_MC2_r1Inst_XORInst_0_0_n5 ), .B(
        \Red_MCInst_MC2_r1Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback[27]) );
  XNOR2_X1 \Red_MCInst_MC2_r1Inst_XORInst_0_0_U2  ( .A(
        \Red_MCInst_MC2_v3_3 [2]), .B(\Red_MCInst_MC2_v2_1 [0]), .ZN(
        \Red_MCInst_MC2_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \Red_MCInst_MC2_r1Inst_XORInst_0_0_U1  ( .A(\Red_MCInst_MC2_v0_1 [0]), .B(\Red_MCInst_MC2_v1_2 [1]), .Z(\Red_MCInst_MC2_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \Red_MCInst_MC2_r1Inst_XORInst_0_1_U3  ( .A(
        \Red_MCInst_MC2_r1Inst_XORInst_0_1_n5 ), .B(
        \Red_MCInst_MC2_r1Inst_XORInst_0_1_n4 ), .ZN(Red_Feedback[28]) );
  XNOR2_X1 \Red_MCInst_MC2_r1Inst_XORInst_0_1_U2  ( .A(
        \Red_MCInst_MC2_v3_1 [1]), .B(\Red_MCInst_MC2_v2_1 [1]), .ZN(
        \Red_MCInst_MC2_r1Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \Red_MCInst_MC2_r1Inst_XORInst_0_1_U1  ( .A(\Red_MCInst_MC2_v0_1 [1]), .B(\Red_MCInst_MC2_v1_1 [1]), .Z(\Red_MCInst_MC2_r1Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \Red_MCInst_MC2_r1Inst_XORInst_0_2_U3  ( .A(
        \Red_MCInst_MC2_r1Inst_XORInst_0_2_n5 ), .B(
        \Red_MCInst_MC2_r1Inst_XORInst_0_2_n4 ), .ZN(Red_Feedback[29]) );
  XNOR2_X1 \Red_MCInst_MC2_r1Inst_XORInst_0_2_U2  ( .A(
        \Red_MCInst_MC2_v3_1 [2]), .B(\Red_MCInst_MC2_v2_1 [2]), .ZN(
        \Red_MCInst_MC2_r1Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \Red_MCInst_MC2_r1Inst_XORInst_0_2_U1  ( .A(\Red_MCInst_MC2_v0_1 [2]), .B(\Red_MCInst_MC2_v1_1 [2]), .Z(\Red_MCInst_MC2_r1Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \Red_MCInst_MC2_r2Inst_XORInst_0_0_U3  ( .A(
        \Red_MCInst_MC2_r2Inst_XORInst_0_0_n5 ), .B(
        \Red_MCInst_MC2_r2Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback[15]) );
  XNOR2_X1 \Red_MCInst_MC2_r2Inst_XORInst_0_0_U2  ( .A(
        \Red_MCInst_MC2_v3_2 [0]), .B(\Red_MCInst_MC2_v2_2 [0]), .ZN(
        \Red_MCInst_MC2_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \Red_MCInst_MC2_r2Inst_XORInst_0_0_U1  ( .A(\Red_MCInst_MC2_v0_2 [0]), .B(\Red_MCInst_MC2_v1_2 [0]), .Z(\Red_MCInst_MC2_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \Red_MCInst_MC2_r2Inst_XORInst_0_1_U3  ( .A(
        \Red_MCInst_MC2_r2Inst_XORInst_0_1_n5 ), .B(
        \Red_MCInst_MC2_r2Inst_XORInst_0_1_n4 ), .ZN(Red_Feedback[16]) );
  XNOR2_X1 \Red_MCInst_MC2_r2Inst_XORInst_0_1_U2  ( .A(
        \Red_MCInst_MC2_v3_2 [1]), .B(\Red_MCInst_MC2_v2_2 [1]), .ZN(
        \Red_MCInst_MC2_r2Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \Red_MCInst_MC2_r2Inst_XORInst_0_1_U1  ( .A(\Red_MCInst_MC2_v0_2 [1]), .B(\Red_MCInst_MC2_v1_2 [1]), .Z(\Red_MCInst_MC2_r2Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \Red_MCInst_MC2_r2Inst_XORInst_0_2_U3  ( .A(
        \Red_MCInst_MC2_r2Inst_XORInst_0_2_n5 ), .B(
        \Red_MCInst_MC2_r2Inst_XORInst_0_2_n4 ), .ZN(Red_Feedback[17]) );
  XNOR2_X1 \Red_MCInst_MC2_r2Inst_XORInst_0_2_U2  ( .A(
        \Red_MCInst_MC2_v3_2 [2]), .B(\Red_MCInst_MC2_v2_2 [2]), .ZN(
        \Red_MCInst_MC2_r2Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \Red_MCInst_MC2_r2Inst_XORInst_0_2_U1  ( .A(\Red_MCInst_MC2_v0_2 [2]), .B(\Red_MCInst_MC2_v1_2 [2]), .Z(\Red_MCInst_MC2_r2Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \Red_MCInst_MC2_r3Inst_XORInst_0_0_U3  ( .A(
        \Red_MCInst_MC2_r3Inst_XORInst_0_0_n5 ), .B(
        \Red_MCInst_MC2_r3Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback[3]) );
  XNOR2_X1 \Red_MCInst_MC2_r3Inst_XORInst_0_0_U2  ( .A(
        \Red_MCInst_MC2_v3_3 [0]), .B(\Red_MCInst_MC2_v2_3 [0]), .ZN(
        \Red_MCInst_MC2_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \Red_MCInst_MC2_r3Inst_XORInst_0_0_U1  ( .A(\Red_MCInst_MC2_v0_3 [0]), .B(\Red_MCInst_MC2_v1_3 [0]), .Z(\Red_MCInst_MC2_r3Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \Red_MCInst_MC2_r3Inst_XORInst_0_1_U3  ( .A(
        \Red_MCInst_MC2_r3Inst_XORInst_0_1_n5 ), .B(
        \Red_MCInst_MC2_r3Inst_XORInst_0_1_n4 ), .ZN(Red_Feedback[4]) );
  XNOR2_X1 \Red_MCInst_MC2_r3Inst_XORInst_0_1_U2  ( .A(
        \Red_MCInst_MC2_v3_3 [1]), .B(\Red_MCInst_MC2_v2_3 [1]), .ZN(
        \Red_MCInst_MC2_r3Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \Red_MCInst_MC2_r3Inst_XORInst_0_1_U1  ( .A(\Red_MCInst_MC2_v0_3 [1]), .B(\Red_MCInst_MC2_v1_3 [1]), .Z(\Red_MCInst_MC2_r3Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \Red_MCInst_MC2_r3Inst_XORInst_0_2_U3  ( .A(
        \Red_MCInst_MC2_r3Inst_XORInst_0_2_n5 ), .B(
        \Red_MCInst_MC2_r3Inst_XORInst_0_2_n4 ), .ZN(Red_Feedback[5]) );
  XNOR2_X1 \Red_MCInst_MC2_r3Inst_XORInst_0_2_U2  ( .A(
        \Red_MCInst_MC2_v3_3 [2]), .B(\Red_MCInst_MC2_v2_3 [2]), .ZN(
        \Red_MCInst_MC2_r3Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \Red_MCInst_MC2_r3Inst_XORInst_0_2_U1  ( .A(\Red_MCInst_MC2_v0_3 [2]), .B(\Red_MCInst_MC2_v1_3 [2]), .Z(\Red_MCInst_MC2_r3Inst_XORInst_0_2_n5 ) );
  XOR2_X1 \Red_MCInst_MC3_v0_2Inst_0_U3  ( .A(\MCInst_MC3_v0_3 [3]), .B(
        \Red_MCInst_MC3_v0_1 [0]), .Z(\Red_MCInst_MC3_v0_2 [0]) );
  XOR2_X1 \Red_MCInst_MC3_v0_3Inst_0_U3  ( .A(\Red_MCInst_MC3_v0_0 [0]), .B(
        \Red_MCInst_MC3_v0_2 [2]), .Z(\Red_MCInst_MC3_v0_3 [0]) );
  XNOR2_X1 \Red_MCInst_MC3_v1_0Inst_0_U4  ( .A(\Red_MCInst_MC3_v1_0Inst_0_n2 ), 
        .B(\Red_MCInst_MC3_v1_2 [1]), .ZN(\Red_MCInst_MC3_v1_0 [0]) );
  XNOR2_X1 \Red_MCInst_MC3_v1_0Inst_0_U3  ( .A(\MCInst_MC3_v1_3 [3]), .B(
        \MCInst_MC3_v1_0 [0]), .ZN(\Red_MCInst_MC3_v1_0Inst_0_n2 ) );
  XOR2_X1 \Red_MCInst_MC3_v1_2Inst_0_U3  ( .A(\Red_MCInst_MC3_v1_2 [1]), .B(
        \Red_MCInst_MC3_v1_1 [2]), .Z(\Red_MCInst_MC3_v1_2 [0]) );
  XOR2_X1 \Red_MCInst_MC3_v1_3Inst_0_U3  ( .A(\MCInst_MC3_v1_0 [0]), .B(
        \Red_MCInst_MC3_v1_2 [1]), .Z(\Red_MCInst_MC3_v1_3 [0]) );
  XOR2_X1 \Red_MCInst_MC3_v2_0Inst_0_U3  ( .A(\Red_MCInst_MC3_v2_1 [1]), .B(
        \MCInst_MC3_v2_0 [2]), .Z(\Red_MCInst_MC3_v2_0 [0]) );
  XOR2_X1 \Red_MCInst_MC3_v2_1Inst_0_U3  ( .A(\MCInst_MC3_v2_0 [2]), .B(
        \MCInst_MC3_v2_0 [3]), .Z(\Red_MCInst_MC3_v2_1 [0]) );
  XNOR2_X1 \Red_MCInst_MC3_v2_2Inst_0_U4  ( .A(\Red_MCInst_MC3_v2_2Inst_0_n2 ), 
        .B(\MCInst_MC3_v2_0 [2]), .ZN(\Red_MCInst_MC3_v2_2 [0]) );
  XNOR2_X1 \Red_MCInst_MC3_v2_2Inst_0_U3  ( .A(\Red_MCInst_MC3_v2_2 [1]), .B(
        \Red_MCInst_MC3_v2_1 [1]), .ZN(\Red_MCInst_MC3_v2_2Inst_0_n2 ) );
  XNOR2_X1 \Red_MCInst_MC3_v2_3Inst_0_U4  ( .A(\Red_MCInst_MC3_v2_3Inst_0_n2 ), 
        .B(\MCInst_MC3_v2_0 [3]), .ZN(\Red_MCInst_MC3_v2_3 [0]) );
  XNOR2_X1 \Red_MCInst_MC3_v2_3Inst_0_U3  ( .A(\Red_MCInst_MC3_v2_2 [1]), .B(
        \Red_MCInst_MC3_v2_1 [1]), .ZN(\Red_MCInst_MC3_v2_3Inst_0_n2 ) );
  XOR2_X1 \Red_MCInst_MC3_v3_0Inst_0_U3  ( .A(\MCInst_MC3_v3_2 [3]), .B(
        \Red_MCInst_MC3_v3_3 [2]), .Z(\Red_MCInst_MC3_v3_0 [0]) );
  XNOR2_X1 \Red_MCInst_MC3_v3_2Inst_0_U5  ( .A(\Red_MCInst_MC3_v3_2Inst_0_n4 ), 
        .B(\Red_MCInst_MC3_v3_2Inst_0_n3 ), .ZN(\Red_MCInst_MC3_v3_2 [0]) );
  XNOR2_X1 \Red_MCInst_MC3_v3_2Inst_0_U4  ( .A(\Red_MCInst_MC3_v3_3 [2]), .B(
        \MCInst_MC3_v3_2 [3]), .ZN(\Red_MCInst_MC3_v3_2Inst_0_n3 ) );
  XOR2_X1 \Red_MCInst_MC3_v3_2Inst_0_U3  ( .A(\MCInst_MC3_v3_0 [3]), .B(
        \Red_MCInst_MC3_v3_1 [2]), .Z(\Red_MCInst_MC3_v3_2Inst_0_n4 ) );
  XOR2_X1 \Red_MCInst_MC3_v3_3Inst_0_U3  ( .A(\MCInst_MC3_v3_0 [3]), .B(
        \Red_MCInst_MC3_v3_1 [2]), .Z(\Red_MCInst_MC3_v3_3 [0]) );
  XOR2_X1 \Red_MCInst_MC3_v0_0Inst_1_U3  ( .A(\Red_MCInst_MC3_v0_2 [2]), .B(
        \Red_MCInst_MC3_v0_1 [0]), .Z(\Red_MCInst_MC3_v0_0 [1]) );
  XNOR2_X1 \Red_MCInst_MC3_v0_1Inst_1_U4  ( .A(\Red_MCInst_MC3_v0_1Inst_1_n2 ), 
        .B(\MCInst_MC3_v0_3 [3]), .ZN(\Red_MCInst_MC3_v0_1 [1]) );
  XNOR2_X1 \Red_MCInst_MC3_v0_1Inst_1_U3  ( .A(\Red_MCInst_MC3_v0_1 [0]), .B(
        \Red_MCInst_MC3_v0_0 [0]), .ZN(\Red_MCInst_MC3_v0_1Inst_1_n2 ) );
  XOR2_X1 \Red_MCInst_MC3_v0_2Inst_1_U3  ( .A(\Red_MCInst_MC3_v0_0 [0]), .B(
        \Red_MCInst_MC3_v0_2 [2]), .Z(\Red_MCInst_MC3_v0_2 [1]) );
  XOR2_X1 \Red_MCInst_MC3_v0_3Inst_1_U3  ( .A(\Red_MCInst_MC3_v0_0 [0]), .B(
        \MCInst_MC3_v0_3 [3]), .Z(\Red_MCInst_MC3_v0_3 [1]) );
  XNOR2_X1 \Red_MCInst_MC3_v1_0Inst_1_U4  ( .A(\Red_MCInst_MC3_v1_0Inst_1_n2 ), 
        .B(\Red_MCInst_MC3_v1_2 [1]), .ZN(\Red_MCInst_MC3_v1_0 [1]) );
  XNOR2_X1 \Red_MCInst_MC3_v1_0Inst_1_U3  ( .A(\Red_MCInst_MC3_v1_1 [2]), .B(
        \MCInst_MC3_v1_0 [0]), .ZN(\Red_MCInst_MC3_v1_0Inst_1_n2 ) );
  XNOR2_X1 \Red_MCInst_MC3_v1_1Inst_1_U5  ( .A(\Red_MCInst_MC3_v1_1Inst_1_n4 ), 
        .B(\Red_MCInst_MC3_v1_1Inst_1_n3 ), .ZN(\Red_MCInst_MC3_v1_1 [1]) );
  XNOR2_X1 \Red_MCInst_MC3_v1_1Inst_1_U4  ( .A(\Red_MCInst_MC3_v1_2 [1]), .B(
        \MCInst_MC3_v1_0 [0]), .ZN(\Red_MCInst_MC3_v1_1Inst_1_n3 ) );
  XOR2_X1 \Red_MCInst_MC3_v1_1Inst_1_U3  ( .A(\MCInst_MC3_v1_3 [3]), .B(
        \Red_MCInst_MC3_v1_1 [2]), .Z(\Red_MCInst_MC3_v1_1Inst_1_n4 ) );
  XOR2_X1 \Red_MCInst_MC3_v1_3Inst_1_U3  ( .A(\MCInst_MC3_v1_0 [0]), .B(
        \MCInst_MC3_v1_3 [3]), .Z(\Red_MCInst_MC3_v1_3 [1]) );
  XOR2_X1 \Red_MCInst_MC3_v2_0Inst_1_U3  ( .A(\Red_MCInst_MC3_v2_1 [1]), .B(
        \MCInst_MC3_v2_0 [3]), .Z(\Red_MCInst_MC3_v2_0 [1]) );
  XOR2_X1 \Red_MCInst_MC3_v2_3Inst_1_U3  ( .A(\Red_MCInst_MC3_v2_1 [1]), .B(
        \Red_MCInst_MC3_v2_2 [1]), .Z(\Red_MCInst_MC3_v2_3 [1]) );
  XOR2_X1 \Red_MCInst_MC3_v3_0Inst_1_U3  ( .A(\MCInst_MC3_v3_2 [3]), .B(
        \MCInst_MC3_v3_0 [3]), .Z(\Red_MCInst_MC3_v3_0 [1]) );
  XNOR2_X1 \Red_MCInst_MC3_v3_1Inst_1_U5  ( .A(\Red_MCInst_MC3_v3_1Inst_1_n4 ), 
        .B(\Red_MCInst_MC3_v3_1Inst_1_n3 ), .ZN(\Red_MCInst_MC3_v3_1 [1]) );
  XNOR2_X1 \Red_MCInst_MC3_v3_1Inst_1_U4  ( .A(\Red_MCInst_MC3_v3_3 [2]), .B(
        \MCInst_MC3_v3_2 [3]), .ZN(\Red_MCInst_MC3_v3_1Inst_1_n3 ) );
  XOR2_X1 \Red_MCInst_MC3_v3_1Inst_1_U3  ( .A(\MCInst_MC3_v3_0 [3]), .B(
        \Red_MCInst_MC3_v3_1 [2]), .Z(\Red_MCInst_MC3_v3_1Inst_1_n4 ) );
  XOR2_X1 \Red_MCInst_MC3_v3_2Inst_1_U3  ( .A(\Red_MCInst_MC3_v3_3 [2]), .B(
        \MCInst_MC3_v3_0 [3]), .Z(\Red_MCInst_MC3_v3_2 [1]) );
  XOR2_X1 \Red_MCInst_MC3_v3_3Inst_1_U3  ( .A(\MCInst_MC3_v3_2 [3]), .B(
        \Red_MCInst_MC3_v3_3 [2]), .Z(\Red_MCInst_MC3_v3_3 [1]) );
  XNOR2_X1 \Red_MCInst_MC3_v0_0Inst_2_U4  ( .A(\Red_MCInst_MC3_v0_0Inst_2_n2 ), 
        .B(\Red_MCInst_MC3_v0_2 [2]), .ZN(\Red_MCInst_MC3_v0_0 [2]) );
  XNOR2_X1 \Red_MCInst_MC3_v0_0Inst_2_U3  ( .A(\MCInst_MC3_v0_3 [3]), .B(
        \Red_MCInst_MC3_v0_0 [0]), .ZN(\Red_MCInst_MC3_v0_0Inst_2_n2 ) );
  XOR2_X1 \Red_MCInst_MC3_v0_1Inst_2_U3  ( .A(\Red_MCInst_MC3_v0_0 [0]), .B(
        \Red_MCInst_MC3_v0_2 [2]), .Z(\Red_MCInst_MC3_v0_1 [2]) );
  XNOR2_X1 \Red_MCInst_MC3_v0_3Inst_2_U5  ( .A(\Red_MCInst_MC3_v0_3Inst_2_n4 ), 
        .B(\Red_MCInst_MC3_v0_3Inst_2_n3 ), .ZN(\Red_MCInst_MC3_v0_3 [2]) );
  XNOR2_X1 \Red_MCInst_MC3_v0_3Inst_2_U4  ( .A(\Red_MCInst_MC3_v0_2 [2]), .B(
        \Red_MCInst_MC3_v0_0 [0]), .ZN(\Red_MCInst_MC3_v0_3Inst_2_n3 ) );
  XOR2_X1 \Red_MCInst_MC3_v0_3Inst_2_U3  ( .A(\MCInst_MC3_v0_3 [3]), .B(
        \Red_MCInst_MC3_v0_1 [0]), .Z(\Red_MCInst_MC3_v0_3Inst_2_n4 ) );
  XNOR2_X1 \Red_MCInst_MC3_v1_0Inst_2_U4  ( .A(\Red_MCInst_MC3_v1_0Inst_2_n2 ), 
        .B(\MCInst_MC3_v1_3 [3]), .ZN(\Red_MCInst_MC3_v1_0 [2]) );
  XNOR2_X1 \Red_MCInst_MC3_v1_0Inst_2_U3  ( .A(\Red_MCInst_MC3_v1_1 [2]), .B(
        \Red_MCInst_MC3_v1_2 [1]), .ZN(\Red_MCInst_MC3_v1_0Inst_2_n2 ) );
  XNOR2_X1 \Red_MCInst_MC3_v1_2Inst_2_U4  ( .A(\Red_MCInst_MC3_v1_2Inst_2_n2 ), 
        .B(\Red_MCInst_MC3_v1_2 [1]), .ZN(\Red_MCInst_MC3_v1_2 [2]) );
  XNOR2_X1 \Red_MCInst_MC3_v1_2Inst_2_U3  ( .A(\Red_MCInst_MC3_v1_1 [2]), .B(
        \MCInst_MC3_v1_0 [0]), .ZN(\Red_MCInst_MC3_v1_2Inst_2_n2 ) );
  XNOR2_X1 \Red_MCInst_MC3_v1_3Inst_2_U5  ( .A(\Red_MCInst_MC3_v1_3Inst_2_n4 ), 
        .B(\Red_MCInst_MC3_v1_3Inst_2_n3 ), .ZN(\Red_MCInst_MC3_v1_3 [2]) );
  XNOR2_X1 \Red_MCInst_MC3_v1_3Inst_2_U4  ( .A(\Red_MCInst_MC3_v1_2 [1]), .B(
        \MCInst_MC3_v1_0 [0]), .ZN(\Red_MCInst_MC3_v1_3Inst_2_n3 ) );
  XOR2_X1 \Red_MCInst_MC3_v1_3Inst_2_U3  ( .A(\MCInst_MC3_v1_3 [3]), .B(
        \Red_MCInst_MC3_v1_1 [2]), .Z(\Red_MCInst_MC3_v1_3Inst_2_n4 ) );
  XNOR2_X1 \Red_MCInst_MC3_v2_0Inst_2_U5  ( .A(\Red_MCInst_MC3_v2_0Inst_2_n4 ), 
        .B(\Red_MCInst_MC3_v2_0Inst_2_n3 ), .ZN(\Red_MCInst_MC3_v2_0 [2]) );
  XNOR2_X1 \Red_MCInst_MC3_v2_0Inst_2_U4  ( .A(\MCInst_MC3_v2_0 [2]), .B(
        \Red_MCInst_MC3_v2_1 [1]), .ZN(\Red_MCInst_MC3_v2_0Inst_2_n3 ) );
  XOR2_X1 \Red_MCInst_MC3_v2_0Inst_2_U3  ( .A(\MCInst_MC3_v2_0 [3]), .B(
        \Red_MCInst_MC3_v2_2 [1]), .Z(\Red_MCInst_MC3_v2_0Inst_2_n4 ) );
  XOR2_X1 \Red_MCInst_MC3_v2_1Inst_2_U3  ( .A(\Red_MCInst_MC3_v2_1 [1]), .B(
        \Red_MCInst_MC3_v2_2 [1]), .Z(\Red_MCInst_MC3_v2_1 [2]) );
  XOR2_X1 \Red_MCInst_MC3_v2_2Inst_2_U3  ( .A(\MCInst_MC3_v2_0 [3]), .B(
        \Red_MCInst_MC3_v2_2 [1]), .Z(\Red_MCInst_MC3_v2_2 [2]) );
  XOR2_X1 \Red_MCInst_MC3_v2_3Inst_2_U3  ( .A(\Red_MCInst_MC3_v2_1 [1]), .B(
        \MCInst_MC3_v2_0 [3]), .Z(\Red_MCInst_MC3_v2_3 [2]) );
  XNOR2_X1 \Red_MCInst_MC3_v3_0Inst_2_U5  ( .A(\Red_MCInst_MC3_v3_0Inst_2_n4 ), 
        .B(\Red_MCInst_MC3_v3_0Inst_2_n3 ), .ZN(\Red_MCInst_MC3_v3_0 [2]) );
  XNOR2_X1 \Red_MCInst_MC3_v3_0Inst_2_U4  ( .A(\Red_MCInst_MC3_v3_3 [2]), .B(
        \MCInst_MC3_v3_2 [3]), .ZN(\Red_MCInst_MC3_v3_0Inst_2_n3 ) );
  XOR2_X1 \Red_MCInst_MC3_v3_0Inst_2_U3  ( .A(\MCInst_MC3_v3_0 [3]), .B(
        \Red_MCInst_MC3_v3_1 [2]), .Z(\Red_MCInst_MC3_v3_0Inst_2_n4 ) );
  XNOR2_X1 \Red_MCInst_MC3_v3_2Inst_2_U4  ( .A(\Red_MCInst_MC3_v3_2Inst_2_n2 ), 
        .B(\MCInst_MC3_v3_0 [3]), .ZN(\Red_MCInst_MC3_v3_2 [2]) );
  XNOR2_X1 \Red_MCInst_MC3_v3_2Inst_2_U3  ( .A(\Red_MCInst_MC3_v3_1 [2]), .B(
        \MCInst_MC3_v3_2 [3]), .ZN(\Red_MCInst_MC3_v3_2Inst_2_n2 ) );
  XNOR2_X1 \Red_MCInst_MC3_r0Inst_XORInst_0_0_U3  ( .A(
        \Red_MCInst_MC3_r0Inst_XORInst_0_0_n5 ), .B(
        \Red_MCInst_MC3_r0Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback[36]) );
  XNOR2_X1 \Red_MCInst_MC3_r0Inst_XORInst_0_0_U2  ( .A(
        \Red_MCInst_MC3_v3_0 [0]), .B(\Red_MCInst_MC3_v2_0 [0]), .ZN(
        \Red_MCInst_MC3_r0Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \Red_MCInst_MC3_r0Inst_XORInst_0_0_U1  ( .A(\Red_MCInst_MC3_v0_0 [0]), .B(\Red_MCInst_MC3_v1_0 [0]), .Z(\Red_MCInst_MC3_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \Red_MCInst_MC3_r0Inst_XORInst_0_1_U3  ( .A(
        \Red_MCInst_MC3_r0Inst_XORInst_0_1_n5 ), .B(
        \Red_MCInst_MC3_r0Inst_XORInst_0_1_n4 ), .ZN(Red_Feedback[37]) );
  XNOR2_X1 \Red_MCInst_MC3_r0Inst_XORInst_0_1_U2  ( .A(
        \Red_MCInst_MC3_v3_0 [1]), .B(\Red_MCInst_MC3_v2_0 [1]), .ZN(
        \Red_MCInst_MC3_r0Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \Red_MCInst_MC3_r0Inst_XORInst_0_1_U1  ( .A(\Red_MCInst_MC3_v0_0 [1]), .B(\Red_MCInst_MC3_v1_0 [1]), .Z(\Red_MCInst_MC3_r0Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \Red_MCInst_MC3_r0Inst_XORInst_0_2_U3  ( .A(
        \Red_MCInst_MC3_r0Inst_XORInst_0_2_n5 ), .B(
        \Red_MCInst_MC3_r0Inst_XORInst_0_2_n4 ), .ZN(Red_Feedback[38]) );
  XNOR2_X1 \Red_MCInst_MC3_r0Inst_XORInst_0_2_U2  ( .A(
        \Red_MCInst_MC3_v3_0 [2]), .B(\Red_MCInst_MC3_v2_0 [2]), .ZN(
        \Red_MCInst_MC3_r0Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \Red_MCInst_MC3_r0Inst_XORInst_0_2_U1  ( .A(\Red_MCInst_MC3_v0_0 [2]), .B(\Red_MCInst_MC3_v1_0 [2]), .Z(\Red_MCInst_MC3_r0Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \Red_MCInst_MC3_r1Inst_XORInst_0_0_U3  ( .A(
        \Red_MCInst_MC3_r1Inst_XORInst_0_0_n5 ), .B(
        \Red_MCInst_MC3_r1Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback[24]) );
  XNOR2_X1 \Red_MCInst_MC3_r1Inst_XORInst_0_0_U2  ( .A(
        \Red_MCInst_MC3_v3_3 [2]), .B(\Red_MCInst_MC3_v2_1 [0]), .ZN(
        \Red_MCInst_MC3_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \Red_MCInst_MC3_r1Inst_XORInst_0_0_U1  ( .A(\Red_MCInst_MC3_v0_1 [0]), .B(\Red_MCInst_MC3_v1_2 [1]), .Z(\Red_MCInst_MC3_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \Red_MCInst_MC3_r1Inst_XORInst_0_1_U3  ( .A(
        \Red_MCInst_MC3_r1Inst_XORInst_0_1_n5 ), .B(
        \Red_MCInst_MC3_r1Inst_XORInst_0_1_n4 ), .ZN(Red_Feedback[25]) );
  XNOR2_X1 \Red_MCInst_MC3_r1Inst_XORInst_0_1_U2  ( .A(
        \Red_MCInst_MC3_v3_1 [1]), .B(\Red_MCInst_MC3_v2_1 [1]), .ZN(
        \Red_MCInst_MC3_r1Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \Red_MCInst_MC3_r1Inst_XORInst_0_1_U1  ( .A(\Red_MCInst_MC3_v0_1 [1]), .B(\Red_MCInst_MC3_v1_1 [1]), .Z(\Red_MCInst_MC3_r1Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \Red_MCInst_MC3_r1Inst_XORInst_0_2_U3  ( .A(
        \Red_MCInst_MC3_r1Inst_XORInst_0_2_n5 ), .B(
        \Red_MCInst_MC3_r1Inst_XORInst_0_2_n4 ), .ZN(Red_Feedback[26]) );
  XNOR2_X1 \Red_MCInst_MC3_r1Inst_XORInst_0_2_U2  ( .A(
        \Red_MCInst_MC3_v3_1 [2]), .B(\Red_MCInst_MC3_v2_1 [2]), .ZN(
        \Red_MCInst_MC3_r1Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \Red_MCInst_MC3_r1Inst_XORInst_0_2_U1  ( .A(\Red_MCInst_MC3_v0_1 [2]), .B(\Red_MCInst_MC3_v1_1 [2]), .Z(\Red_MCInst_MC3_r1Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \Red_MCInst_MC3_r2Inst_XORInst_0_0_U3  ( .A(
        \Red_MCInst_MC3_r2Inst_XORInst_0_0_n5 ), .B(
        \Red_MCInst_MC3_r2Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback[12]) );
  XNOR2_X1 \Red_MCInst_MC3_r2Inst_XORInst_0_0_U2  ( .A(
        \Red_MCInst_MC3_v3_2 [0]), .B(\Red_MCInst_MC3_v2_2 [0]), .ZN(
        \Red_MCInst_MC3_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \Red_MCInst_MC3_r2Inst_XORInst_0_0_U1  ( .A(\Red_MCInst_MC3_v0_2 [0]), .B(\Red_MCInst_MC3_v1_2 [0]), .Z(\Red_MCInst_MC3_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \Red_MCInst_MC3_r2Inst_XORInst_0_1_U3  ( .A(
        \Red_MCInst_MC3_r2Inst_XORInst_0_1_n5 ), .B(
        \Red_MCInst_MC3_r2Inst_XORInst_0_1_n4 ), .ZN(Red_Feedback[13]) );
  XNOR2_X1 \Red_MCInst_MC3_r2Inst_XORInst_0_1_U2  ( .A(
        \Red_MCInst_MC3_v3_2 [1]), .B(\Red_MCInst_MC3_v2_2 [1]), .ZN(
        \Red_MCInst_MC3_r2Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \Red_MCInst_MC3_r2Inst_XORInst_0_1_U1  ( .A(\Red_MCInst_MC3_v0_2 [1]), .B(\Red_MCInst_MC3_v1_2 [1]), .Z(\Red_MCInst_MC3_r2Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \Red_MCInst_MC3_r2Inst_XORInst_0_2_U3  ( .A(
        \Red_MCInst_MC3_r2Inst_XORInst_0_2_n5 ), .B(
        \Red_MCInst_MC3_r2Inst_XORInst_0_2_n4 ), .ZN(Red_Feedback[14]) );
  XNOR2_X1 \Red_MCInst_MC3_r2Inst_XORInst_0_2_U2  ( .A(
        \Red_MCInst_MC3_v3_2 [2]), .B(\Red_MCInst_MC3_v2_2 [2]), .ZN(
        \Red_MCInst_MC3_r2Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \Red_MCInst_MC3_r2Inst_XORInst_0_2_U1  ( .A(\Red_MCInst_MC3_v0_2 [2]), .B(\Red_MCInst_MC3_v1_2 [2]), .Z(\Red_MCInst_MC3_r2Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \Red_MCInst_MC3_r3Inst_XORInst_0_0_U3  ( .A(
        \Red_MCInst_MC3_r3Inst_XORInst_0_0_n5 ), .B(
        \Red_MCInst_MC3_r3Inst_XORInst_0_0_n4 ), .ZN(Red_Feedback[0]) );
  XNOR2_X1 \Red_MCInst_MC3_r3Inst_XORInst_0_0_U2  ( .A(
        \Red_MCInst_MC3_v3_3 [0]), .B(\Red_MCInst_MC3_v2_3 [0]), .ZN(
        \Red_MCInst_MC3_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 \Red_MCInst_MC3_r3Inst_XORInst_0_0_U1  ( .A(\Red_MCInst_MC3_v0_3 [0]), .B(\Red_MCInst_MC3_v1_3 [0]), .Z(\Red_MCInst_MC3_r3Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 \Red_MCInst_MC3_r3Inst_XORInst_0_1_U3  ( .A(
        \Red_MCInst_MC3_r3Inst_XORInst_0_1_n5 ), .B(
        \Red_MCInst_MC3_r3Inst_XORInst_0_1_n4 ), .ZN(Red_Feedback[1]) );
  XNOR2_X1 \Red_MCInst_MC3_r3Inst_XORInst_0_1_U2  ( .A(
        \Red_MCInst_MC3_v3_3 [1]), .B(\Red_MCInst_MC3_v2_3 [1]), .ZN(
        \Red_MCInst_MC3_r3Inst_XORInst_0_1_n4 ) );
  XOR2_X1 \Red_MCInst_MC3_r3Inst_XORInst_0_1_U1  ( .A(\Red_MCInst_MC3_v0_3 [1]), .B(\Red_MCInst_MC3_v1_3 [1]), .Z(\Red_MCInst_MC3_r3Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 \Red_MCInst_MC3_r3Inst_XORInst_0_2_U3  ( .A(
        \Red_MCInst_MC3_r3Inst_XORInst_0_2_n5 ), .B(
        \Red_MCInst_MC3_r3Inst_XORInst_0_2_n4 ), .ZN(Red_Feedback[2]) );
  XNOR2_X1 \Red_MCInst_MC3_r3Inst_XORInst_0_2_U2  ( .A(
        \Red_MCInst_MC3_v3_3 [2]), .B(\Red_MCInst_MC3_v2_3 [2]), .ZN(
        \Red_MCInst_MC3_r3Inst_XORInst_0_2_n4 ) );
  XOR2_X1 \Red_MCInst_MC3_r3Inst_XORInst_0_2_U1  ( .A(\Red_MCInst_MC3_v0_3 [2]), .B(\Red_MCInst_MC3_v1_3 [2]), .Z(\Red_MCInst_MC3_r3Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 \Red_KeyInst_LFInst_0_LFInst_0_U4  ( .A(
        \Red_KeyInst_LFInst_0_LFInst_0_n2 ), .B(Key[1]), .ZN(Red_RoundKey[0])
         );
  XNOR2_X1 \Red_KeyInst_LFInst_0_LFInst_0_U3  ( .A(Key[2]), .B(Key[0]), .ZN(
        \Red_KeyInst_LFInst_0_LFInst_0_n2 ) );
  XNOR2_X1 \Red_KeyInst_LFInst_0_LFInst_1_U4  ( .A(
        \Red_KeyInst_LFInst_0_LFInst_1_n2 ), .B(Key[1]), .ZN(Red_RoundKey[1])
         );
  XNOR2_X1 \Red_KeyInst_LFInst_0_LFInst_1_U3  ( .A(Key[3]), .B(Key[0]), .ZN(
        \Red_KeyInst_LFInst_0_LFInst_1_n2 ) );
  XNOR2_X1 \Red_KeyInst_LFInst_0_LFInst_2_U4  ( .A(
        \Red_KeyInst_LFInst_0_LFInst_2_n2 ), .B(Key[2]), .ZN(Red_RoundKey[2])
         );
  XNOR2_X1 \Red_KeyInst_LFInst_0_LFInst_2_U3  ( .A(Key[3]), .B(Key[1]), .ZN(
        \Red_KeyInst_LFInst_0_LFInst_2_n2 ) );
  XNOR2_X1 \Red_KeyInst_LFInst_1_LFInst_0_U4  ( .A(
        \Red_KeyInst_LFInst_1_LFInst_0_n2 ), .B(Key[5]), .ZN(Red_RoundKey[3])
         );
  XNOR2_X1 \Red_KeyInst_LFInst_1_LFInst_0_U3  ( .A(Key[6]), .B(Key[4]), .ZN(
        \Red_KeyInst_LFInst_1_LFInst_0_n2 ) );
  XNOR2_X1 \Red_KeyInst_LFInst_1_LFInst_1_U4  ( .A(
        \Red_KeyInst_LFInst_1_LFInst_1_n2 ), .B(Key[5]), .ZN(Red_RoundKey[4])
         );
  XNOR2_X1 \Red_KeyInst_LFInst_1_LFInst_1_U3  ( .A(Key[7]), .B(Key[4]), .ZN(
        \Red_KeyInst_LFInst_1_LFInst_1_n2 ) );
  XNOR2_X1 \Red_KeyInst_LFInst_1_LFInst_2_U4  ( .A(
        \Red_KeyInst_LFInst_1_LFInst_2_n2 ), .B(Key[6]), .ZN(Red_RoundKey[5])
         );
  XNOR2_X1 \Red_KeyInst_LFInst_1_LFInst_2_U3  ( .A(Key[7]), .B(Key[5]), .ZN(
        \Red_KeyInst_LFInst_1_LFInst_2_n2 ) );
  XNOR2_X1 \Red_KeyInst_LFInst_2_LFInst_0_U4  ( .A(
        \Red_KeyInst_LFInst_2_LFInst_0_n2 ), .B(Key[9]), .ZN(Red_RoundKey[6])
         );
  XNOR2_X1 \Red_KeyInst_LFInst_2_LFInst_0_U3  ( .A(Key[10]), .B(Key[8]), .ZN(
        \Red_KeyInst_LFInst_2_LFInst_0_n2 ) );
  XNOR2_X1 \Red_KeyInst_LFInst_2_LFInst_1_U4  ( .A(
        \Red_KeyInst_LFInst_2_LFInst_1_n2 ), .B(Key[9]), .ZN(Red_RoundKey[7])
         );
  XNOR2_X1 \Red_KeyInst_LFInst_2_LFInst_1_U3  ( .A(Key[11]), .B(Key[8]), .ZN(
        \Red_KeyInst_LFInst_2_LFInst_1_n2 ) );
  XNOR2_X1 \Red_KeyInst_LFInst_2_LFInst_2_U4  ( .A(
        \Red_KeyInst_LFInst_2_LFInst_2_n2 ), .B(Key[10]), .ZN(Red_RoundKey[8])
         );
  XNOR2_X1 \Red_KeyInst_LFInst_2_LFInst_2_U3  ( .A(Key[11]), .B(Key[9]), .ZN(
        \Red_KeyInst_LFInst_2_LFInst_2_n2 ) );
  XNOR2_X1 \Red_KeyInst_LFInst_3_LFInst_0_U4  ( .A(
        \Red_KeyInst_LFInst_3_LFInst_0_n2 ), .B(Key[13]), .ZN(Red_RoundKey[9])
         );
  XNOR2_X1 \Red_KeyInst_LFInst_3_LFInst_0_U3  ( .A(Key[14]), .B(Key[12]), .ZN(
        \Red_KeyInst_LFInst_3_LFInst_0_n2 ) );
  XNOR2_X1 \Red_KeyInst_LFInst_3_LFInst_1_U4  ( .A(
        \Red_KeyInst_LFInst_3_LFInst_1_n2 ), .B(Key[13]), .ZN(Red_RoundKey[10]) );
  XNOR2_X1 \Red_KeyInst_LFInst_3_LFInst_1_U3  ( .A(Key[15]), .B(Key[12]), .ZN(
        \Red_KeyInst_LFInst_3_LFInst_1_n2 ) );
  XNOR2_X1 \Red_KeyInst_LFInst_3_LFInst_2_U4  ( .A(
        \Red_KeyInst_LFInst_3_LFInst_2_n2 ), .B(Key[14]), .ZN(Red_RoundKey[11]) );
  XNOR2_X1 \Red_KeyInst_LFInst_3_LFInst_2_U3  ( .A(Key[15]), .B(Key[13]), .ZN(
        \Red_KeyInst_LFInst_3_LFInst_2_n2 ) );
  XNOR2_X1 \Red_KeyInst_LFInst_4_LFInst_0_U4  ( .A(
        \Red_KeyInst_LFInst_4_LFInst_0_n2 ), .B(Key[17]), .ZN(Red_RoundKey[12]) );
  XNOR2_X1 \Red_KeyInst_LFInst_4_LFInst_0_U3  ( .A(Key[18]), .B(Key[16]), .ZN(
        \Red_KeyInst_LFInst_4_LFInst_0_n2 ) );
  XNOR2_X1 \Red_KeyInst_LFInst_4_LFInst_1_U4  ( .A(
        \Red_KeyInst_LFInst_4_LFInst_1_n2 ), .B(Key[17]), .ZN(Red_RoundKey[13]) );
  XNOR2_X1 \Red_KeyInst_LFInst_4_LFInst_1_U3  ( .A(Key[19]), .B(Key[16]), .ZN(
        \Red_KeyInst_LFInst_4_LFInst_1_n2 ) );
  XNOR2_X1 \Red_KeyInst_LFInst_4_LFInst_2_U4  ( .A(
        \Red_KeyInst_LFInst_4_LFInst_2_n2 ), .B(Key[18]), .ZN(Red_RoundKey[14]) );
  XNOR2_X1 \Red_KeyInst_LFInst_4_LFInst_2_U3  ( .A(Key[19]), .B(Key[17]), .ZN(
        \Red_KeyInst_LFInst_4_LFInst_2_n2 ) );
  XNOR2_X1 \Red_KeyInst_LFInst_5_LFInst_0_U4  ( .A(
        \Red_KeyInst_LFInst_5_LFInst_0_n2 ), .B(Key[21]), .ZN(Red_RoundKey[15]) );
  XNOR2_X1 \Red_KeyInst_LFInst_5_LFInst_0_U3  ( .A(Key[22]), .B(Key[20]), .ZN(
        \Red_KeyInst_LFInst_5_LFInst_0_n2 ) );
  XNOR2_X1 \Red_KeyInst_LFInst_5_LFInst_1_U4  ( .A(
        \Red_KeyInst_LFInst_5_LFInst_1_n2 ), .B(Key[21]), .ZN(Red_RoundKey[16]) );
  XNOR2_X1 \Red_KeyInst_LFInst_5_LFInst_1_U3  ( .A(Key[23]), .B(Key[20]), .ZN(
        \Red_KeyInst_LFInst_5_LFInst_1_n2 ) );
  XNOR2_X1 \Red_KeyInst_LFInst_5_LFInst_2_U4  ( .A(
        \Red_KeyInst_LFInst_5_LFInst_2_n2 ), .B(Key[22]), .ZN(Red_RoundKey[17]) );
  XNOR2_X1 \Red_KeyInst_LFInst_5_LFInst_2_U3  ( .A(Key[23]), .B(Key[21]), .ZN(
        \Red_KeyInst_LFInst_5_LFInst_2_n2 ) );
  XNOR2_X1 \Red_KeyInst_LFInst_6_LFInst_0_U4  ( .A(
        \Red_KeyInst_LFInst_6_LFInst_0_n2 ), .B(Key[25]), .ZN(Red_RoundKey[18]) );
  XNOR2_X1 \Red_KeyInst_LFInst_6_LFInst_0_U3  ( .A(Key[26]), .B(Key[24]), .ZN(
        \Red_KeyInst_LFInst_6_LFInst_0_n2 ) );
  XNOR2_X1 \Red_KeyInst_LFInst_6_LFInst_1_U4  ( .A(
        \Red_KeyInst_LFInst_6_LFInst_1_n2 ), .B(Key[25]), .ZN(Red_RoundKey[19]) );
  XNOR2_X1 \Red_KeyInst_LFInst_6_LFInst_1_U3  ( .A(Key[27]), .B(Key[24]), .ZN(
        \Red_KeyInst_LFInst_6_LFInst_1_n2 ) );
  XNOR2_X1 \Red_KeyInst_LFInst_6_LFInst_2_U4  ( .A(
        \Red_KeyInst_LFInst_6_LFInst_2_n2 ), .B(Key[26]), .ZN(Red_RoundKey[20]) );
  XNOR2_X1 \Red_KeyInst_LFInst_6_LFInst_2_U3  ( .A(Key[27]), .B(Key[25]), .ZN(
        \Red_KeyInst_LFInst_6_LFInst_2_n2 ) );
  XNOR2_X1 \Red_KeyInst_LFInst_7_LFInst_0_U4  ( .A(
        \Red_KeyInst_LFInst_7_LFInst_0_n2 ), .B(Key[29]), .ZN(Red_RoundKey[21]) );
  XNOR2_X1 \Red_KeyInst_LFInst_7_LFInst_0_U3  ( .A(Key[30]), .B(Key[28]), .ZN(
        \Red_KeyInst_LFInst_7_LFInst_0_n2 ) );
  XNOR2_X1 \Red_KeyInst_LFInst_7_LFInst_1_U4  ( .A(
        \Red_KeyInst_LFInst_7_LFInst_1_n2 ), .B(Key[29]), .ZN(Red_RoundKey[22]) );
  XNOR2_X1 \Red_KeyInst_LFInst_7_LFInst_1_U3  ( .A(Key[31]), .B(Key[28]), .ZN(
        \Red_KeyInst_LFInst_7_LFInst_1_n2 ) );
  XNOR2_X1 \Red_KeyInst_LFInst_7_LFInst_2_U4  ( .A(
        \Red_KeyInst_LFInst_7_LFInst_2_n2 ), .B(Key[30]), .ZN(Red_RoundKey[23]) );
  XNOR2_X1 \Red_KeyInst_LFInst_7_LFInst_2_U3  ( .A(Key[31]), .B(Key[29]), .ZN(
        \Red_KeyInst_LFInst_7_LFInst_2_n2 ) );
  XNOR2_X1 \Red_KeyInst_LFInst_8_LFInst_0_U4  ( .A(
        \Red_KeyInst_LFInst_8_LFInst_0_n2 ), .B(Key[33]), .ZN(Red_RoundKey[24]) );
  XNOR2_X1 \Red_KeyInst_LFInst_8_LFInst_0_U3  ( .A(Key[34]), .B(Key[32]), .ZN(
        \Red_KeyInst_LFInst_8_LFInst_0_n2 ) );
  XNOR2_X1 \Red_KeyInst_LFInst_8_LFInst_1_U4  ( .A(
        \Red_KeyInst_LFInst_8_LFInst_1_n2 ), .B(Key[33]), .ZN(Red_RoundKey[25]) );
  XNOR2_X1 \Red_KeyInst_LFInst_8_LFInst_1_U3  ( .A(Key[35]), .B(Key[32]), .ZN(
        \Red_KeyInst_LFInst_8_LFInst_1_n2 ) );
  XNOR2_X1 \Red_KeyInst_LFInst_8_LFInst_2_U4  ( .A(
        \Red_KeyInst_LFInst_8_LFInst_2_n2 ), .B(Key[34]), .ZN(Red_RoundKey[26]) );
  XNOR2_X1 \Red_KeyInst_LFInst_8_LFInst_2_U3  ( .A(Key[35]), .B(Key[33]), .ZN(
        \Red_KeyInst_LFInst_8_LFInst_2_n2 ) );
  XNOR2_X1 \Red_KeyInst_LFInst_9_LFInst_0_U4  ( .A(
        \Red_KeyInst_LFInst_9_LFInst_0_n2 ), .B(Key[37]), .ZN(Red_RoundKey[27]) );
  XNOR2_X1 \Red_KeyInst_LFInst_9_LFInst_0_U3  ( .A(Key[38]), .B(Key[36]), .ZN(
        \Red_KeyInst_LFInst_9_LFInst_0_n2 ) );
  XNOR2_X1 \Red_KeyInst_LFInst_9_LFInst_1_U4  ( .A(
        \Red_KeyInst_LFInst_9_LFInst_1_n2 ), .B(Key[37]), .ZN(Red_RoundKey[28]) );
  XNOR2_X1 \Red_KeyInst_LFInst_9_LFInst_1_U3  ( .A(Key[39]), .B(Key[36]), .ZN(
        \Red_KeyInst_LFInst_9_LFInst_1_n2 ) );
  XNOR2_X1 \Red_KeyInst_LFInst_9_LFInst_2_U4  ( .A(
        \Red_KeyInst_LFInst_9_LFInst_2_n2 ), .B(Key[38]), .ZN(Red_RoundKey[29]) );
  XNOR2_X1 \Red_KeyInst_LFInst_9_LFInst_2_U3  ( .A(Key[39]), .B(Key[37]), .ZN(
        \Red_KeyInst_LFInst_9_LFInst_2_n2 ) );
  XNOR2_X1 \Red_KeyInst_LFInst_10_LFInst_0_U4  ( .A(
        \Red_KeyInst_LFInst_10_LFInst_0_n2 ), .B(Key[41]), .ZN(
        Red_RoundKey[30]) );
  XNOR2_X1 \Red_KeyInst_LFInst_10_LFInst_0_U3  ( .A(Key[42]), .B(Key[40]), 
        .ZN(\Red_KeyInst_LFInst_10_LFInst_0_n2 ) );
  XNOR2_X1 \Red_KeyInst_LFInst_10_LFInst_1_U4  ( .A(
        \Red_KeyInst_LFInst_10_LFInst_1_n2 ), .B(Key[41]), .ZN(
        Red_RoundKey[31]) );
  XNOR2_X1 \Red_KeyInst_LFInst_10_LFInst_1_U3  ( .A(Key[43]), .B(Key[40]), 
        .ZN(\Red_KeyInst_LFInst_10_LFInst_1_n2 ) );
  XNOR2_X1 \Red_KeyInst_LFInst_10_LFInst_2_U4  ( .A(
        \Red_KeyInst_LFInst_10_LFInst_2_n2 ), .B(Key[42]), .ZN(
        Red_RoundKey[32]) );
  XNOR2_X1 \Red_KeyInst_LFInst_10_LFInst_2_U3  ( .A(Key[43]), .B(Key[41]), 
        .ZN(\Red_KeyInst_LFInst_10_LFInst_2_n2 ) );
  XNOR2_X1 \Red_KeyInst_LFInst_11_LFInst_0_U4  ( .A(
        \Red_KeyInst_LFInst_11_LFInst_0_n2 ), .B(Key[45]), .ZN(
        Red_RoundKey[33]) );
  XNOR2_X1 \Red_KeyInst_LFInst_11_LFInst_0_U3  ( .A(Key[46]), .B(Key[44]), 
        .ZN(\Red_KeyInst_LFInst_11_LFInst_0_n2 ) );
  XNOR2_X1 \Red_KeyInst_LFInst_11_LFInst_1_U4  ( .A(
        \Red_KeyInst_LFInst_11_LFInst_1_n2 ), .B(Key[45]), .ZN(
        Red_RoundKey[34]) );
  XNOR2_X1 \Red_KeyInst_LFInst_11_LFInst_1_U3  ( .A(Key[47]), .B(Key[44]), 
        .ZN(\Red_KeyInst_LFInst_11_LFInst_1_n2 ) );
  XNOR2_X1 \Red_KeyInst_LFInst_11_LFInst_2_U4  ( .A(
        \Red_KeyInst_LFInst_11_LFInst_2_n2 ), .B(Key[46]), .ZN(
        Red_RoundKey[35]) );
  XNOR2_X1 \Red_KeyInst_LFInst_11_LFInst_2_U3  ( .A(Key[47]), .B(Key[45]), 
        .ZN(\Red_KeyInst_LFInst_11_LFInst_2_n2 ) );
  XNOR2_X1 \Red_KeyInst_LFInst_12_LFInst_0_U4  ( .A(
        \Red_KeyInst_LFInst_12_LFInst_0_n2 ), .B(Key[49]), .ZN(
        Red_RoundKey[36]) );
  XNOR2_X1 \Red_KeyInst_LFInst_12_LFInst_0_U3  ( .A(Key[50]), .B(Key[48]), 
        .ZN(\Red_KeyInst_LFInst_12_LFInst_0_n2 ) );
  XNOR2_X1 \Red_KeyInst_LFInst_12_LFInst_1_U4  ( .A(
        \Red_KeyInst_LFInst_12_LFInst_1_n2 ), .B(Key[49]), .ZN(
        Red_RoundKey[37]) );
  XNOR2_X1 \Red_KeyInst_LFInst_12_LFInst_1_U3  ( .A(Key[51]), .B(Key[48]), 
        .ZN(\Red_KeyInst_LFInst_12_LFInst_1_n2 ) );
  XNOR2_X1 \Red_KeyInst_LFInst_12_LFInst_2_U4  ( .A(
        \Red_KeyInst_LFInst_12_LFInst_2_n2 ), .B(Key[50]), .ZN(
        Red_RoundKey[38]) );
  XNOR2_X1 \Red_KeyInst_LFInst_12_LFInst_2_U3  ( .A(Key[51]), .B(Key[49]), 
        .ZN(\Red_KeyInst_LFInst_12_LFInst_2_n2 ) );
  XNOR2_X1 \Red_KeyInst_LFInst_13_LFInst_0_U4  ( .A(
        \Red_KeyInst_LFInst_13_LFInst_0_n2 ), .B(Key[53]), .ZN(
        Red_RoundKey[39]) );
  XNOR2_X1 \Red_KeyInst_LFInst_13_LFInst_0_U3  ( .A(Key[54]), .B(Key[52]), 
        .ZN(\Red_KeyInst_LFInst_13_LFInst_0_n2 ) );
  XNOR2_X1 \Red_KeyInst_LFInst_13_LFInst_1_U4  ( .A(
        \Red_KeyInst_LFInst_13_LFInst_1_n2 ), .B(Key[53]), .ZN(
        Red_RoundKey[40]) );
  XNOR2_X1 \Red_KeyInst_LFInst_13_LFInst_1_U3  ( .A(Key[55]), .B(Key[52]), 
        .ZN(\Red_KeyInst_LFInst_13_LFInst_1_n2 ) );
  XNOR2_X1 \Red_KeyInst_LFInst_13_LFInst_2_U4  ( .A(
        \Red_KeyInst_LFInst_13_LFInst_2_n2 ), .B(Key[54]), .ZN(
        Red_RoundKey[41]) );
  XNOR2_X1 \Red_KeyInst_LFInst_13_LFInst_2_U3  ( .A(Key[55]), .B(Key[53]), 
        .ZN(\Red_KeyInst_LFInst_13_LFInst_2_n2 ) );
  XNOR2_X1 \Red_KeyInst_LFInst_14_LFInst_0_U4  ( .A(
        \Red_KeyInst_LFInst_14_LFInst_0_n2 ), .B(Key[57]), .ZN(
        Red_RoundKey[42]) );
  XNOR2_X1 \Red_KeyInst_LFInst_14_LFInst_0_U3  ( .A(Key[58]), .B(Key[56]), 
        .ZN(\Red_KeyInst_LFInst_14_LFInst_0_n2 ) );
  XNOR2_X1 \Red_KeyInst_LFInst_14_LFInst_1_U4  ( .A(
        \Red_KeyInst_LFInst_14_LFInst_1_n2 ), .B(Key[57]), .ZN(
        Red_RoundKey[43]) );
  XNOR2_X1 \Red_KeyInst_LFInst_14_LFInst_1_U3  ( .A(Key[59]), .B(Key[56]), 
        .ZN(\Red_KeyInst_LFInst_14_LFInst_1_n2 ) );
  XNOR2_X1 \Red_KeyInst_LFInst_14_LFInst_2_U4  ( .A(
        \Red_KeyInst_LFInst_14_LFInst_2_n2 ), .B(Key[58]), .ZN(
        Red_RoundKey[44]) );
  XNOR2_X1 \Red_KeyInst_LFInst_14_LFInst_2_U3  ( .A(Key[59]), .B(Key[57]), 
        .ZN(\Red_KeyInst_LFInst_14_LFInst_2_n2 ) );
  XNOR2_X1 \Red_KeyInst_LFInst_15_LFInst_0_U4  ( .A(
        \Red_KeyInst_LFInst_15_LFInst_0_n2 ), .B(Key[61]), .ZN(
        Red_RoundKey[45]) );
  XNOR2_X1 \Red_KeyInst_LFInst_15_LFInst_0_U3  ( .A(Key[62]), .B(Key[60]), 
        .ZN(\Red_KeyInst_LFInst_15_LFInst_0_n2 ) );
  XNOR2_X1 \Red_KeyInst_LFInst_15_LFInst_1_U4  ( .A(
        \Red_KeyInst_LFInst_15_LFInst_1_n2 ), .B(Key[61]), .ZN(
        Red_RoundKey[46]) );
  XNOR2_X1 \Red_KeyInst_LFInst_15_LFInst_1_U3  ( .A(Key[63]), .B(Key[60]), 
        .ZN(\Red_KeyInst_LFInst_15_LFInst_1_n2 ) );
  XNOR2_X1 \Red_KeyInst_LFInst_15_LFInst_2_U4  ( .A(
        \Red_KeyInst_LFInst_15_LFInst_2_n2 ), .B(Key[62]), .ZN(
        Red_RoundKey[47]) );
  XNOR2_X1 \Red_KeyInst_LFInst_15_LFInst_2_U3  ( .A(Key[63]), .B(Key[61]), 
        .ZN(\Red_KeyInst_LFInst_15_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_0_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_0_LFInst_0_n2 ), .B(AddRoundKeyOutput[1]), 
        .ZN(Red_SignaltoCheck[0]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_0_LFInst_0_U3  ( .A(AddRoundKeyOutput[2]), 
        .B(AddRoundKeyOutput[0]), .ZN(\Red_ToCheckInst_LFInst_0_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_0_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_0_LFInst_1_n2 ), .B(AddRoundKeyOutput[1]), 
        .ZN(Red_SignaltoCheck[1]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_0_LFInst_1_U3  ( .A(AddRoundKeyOutput[3]), 
        .B(AddRoundKeyOutput[0]), .ZN(\Red_ToCheckInst_LFInst_0_LFInst_1_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_0_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_0_LFInst_2_n2 ), .B(AddRoundKeyOutput[2]), 
        .ZN(Red_SignaltoCheck[2]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_0_LFInst_2_U3  ( .A(AddRoundKeyOutput[3]), 
        .B(AddRoundKeyOutput[1]), .ZN(\Red_ToCheckInst_LFInst_0_LFInst_2_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_1_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_1_LFInst_0_n2 ), .B(AddRoundKeyOutput[5]), 
        .ZN(Red_SignaltoCheck[3]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_1_LFInst_0_U3  ( .A(AddRoundKeyOutput[6]), 
        .B(AddRoundKeyOutput[4]), .ZN(\Red_ToCheckInst_LFInst_1_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_1_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_1_LFInst_1_n2 ), .B(AddRoundKeyOutput[5]), 
        .ZN(Red_SignaltoCheck[4]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_1_LFInst_1_U3  ( .A(AddRoundKeyOutput[7]), 
        .B(AddRoundKeyOutput[4]), .ZN(\Red_ToCheckInst_LFInst_1_LFInst_1_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_1_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_1_LFInst_2_n2 ), .B(AddRoundKeyOutput[6]), 
        .ZN(Red_SignaltoCheck[5]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_1_LFInst_2_U3  ( .A(AddRoundKeyOutput[7]), 
        .B(AddRoundKeyOutput[5]), .ZN(\Red_ToCheckInst_LFInst_1_LFInst_2_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_2_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_2_LFInst_0_n2 ), .B(AddRoundKeyOutput[9]), 
        .ZN(Red_SignaltoCheck[6]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_2_LFInst_0_U3  ( .A(AddRoundKeyOutput[10]), 
        .B(AddRoundKeyOutput[8]), .ZN(\Red_ToCheckInst_LFInst_2_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_2_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_2_LFInst_1_n2 ), .B(AddRoundKeyOutput[9]), 
        .ZN(Red_SignaltoCheck[7]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_2_LFInst_1_U3  ( .A(AddRoundKeyOutput[11]), 
        .B(AddRoundKeyOutput[8]), .ZN(\Red_ToCheckInst_LFInst_2_LFInst_1_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_2_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_2_LFInst_2_n2 ), .B(AddRoundKeyOutput[10]), 
        .ZN(Red_SignaltoCheck[8]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_2_LFInst_2_U3  ( .A(AddRoundKeyOutput[11]), 
        .B(AddRoundKeyOutput[9]), .ZN(\Red_ToCheckInst_LFInst_2_LFInst_2_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_3_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_3_LFInst_0_n2 ), .B(AddRoundKeyOutput[13]), 
        .ZN(Red_SignaltoCheck[9]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_3_LFInst_0_U3  ( .A(AddRoundKeyOutput[14]), 
        .B(AddRoundKeyOutput[12]), .ZN(\Red_ToCheckInst_LFInst_3_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_3_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_3_LFInst_1_n2 ), .B(AddRoundKeyOutput[13]), 
        .ZN(Red_SignaltoCheck[10]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_3_LFInst_1_U3  ( .A(AddRoundKeyOutput[15]), 
        .B(AddRoundKeyOutput[12]), .ZN(\Red_ToCheckInst_LFInst_3_LFInst_1_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_3_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_3_LFInst_2_n2 ), .B(AddRoundKeyOutput[14]), 
        .ZN(Red_SignaltoCheck[11]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_3_LFInst_2_U3  ( .A(AddRoundKeyOutput[15]), 
        .B(AddRoundKeyOutput[13]), .ZN(\Red_ToCheckInst_LFInst_3_LFInst_2_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_4_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_4_LFInst_0_n2 ), .B(AddRoundKeyOutput[17]), 
        .ZN(Red_SignaltoCheck[12]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_4_LFInst_0_U3  ( .A(AddRoundKeyOutput[18]), 
        .B(AddRoundKeyOutput[16]), .ZN(\Red_ToCheckInst_LFInst_4_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_4_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_4_LFInst_1_n2 ), .B(AddRoundKeyOutput[17]), 
        .ZN(Red_SignaltoCheck[13]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_4_LFInst_1_U3  ( .A(AddRoundKeyOutput[19]), 
        .B(AddRoundKeyOutput[16]), .ZN(\Red_ToCheckInst_LFInst_4_LFInst_1_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_4_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_4_LFInst_2_n2 ), .B(AddRoundKeyOutput[18]), 
        .ZN(Red_SignaltoCheck[14]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_4_LFInst_2_U3  ( .A(AddRoundKeyOutput[19]), 
        .B(AddRoundKeyOutput[17]), .ZN(\Red_ToCheckInst_LFInst_4_LFInst_2_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_5_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_5_LFInst_0_n2 ), .B(AddRoundKeyOutput[21]), 
        .ZN(Red_SignaltoCheck[15]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_5_LFInst_0_U3  ( .A(AddRoundKeyOutput[22]), 
        .B(AddRoundKeyOutput[20]), .ZN(\Red_ToCheckInst_LFInst_5_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_5_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_5_LFInst_1_n2 ), .B(AddRoundKeyOutput[21]), 
        .ZN(Red_SignaltoCheck[16]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_5_LFInst_1_U3  ( .A(AddRoundKeyOutput[23]), 
        .B(AddRoundKeyOutput[20]), .ZN(\Red_ToCheckInst_LFInst_5_LFInst_1_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_5_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_5_LFInst_2_n2 ), .B(AddRoundKeyOutput[22]), 
        .ZN(Red_SignaltoCheck[17]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_5_LFInst_2_U3  ( .A(AddRoundKeyOutput[23]), 
        .B(AddRoundKeyOutput[21]), .ZN(\Red_ToCheckInst_LFInst_5_LFInst_2_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_6_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_6_LFInst_0_n2 ), .B(AddRoundKeyOutput[25]), 
        .ZN(Red_SignaltoCheck[18]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_6_LFInst_0_U3  ( .A(AddRoundKeyOutput[26]), 
        .B(AddRoundKeyOutput[24]), .ZN(\Red_ToCheckInst_LFInst_6_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_6_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_6_LFInst_1_n2 ), .B(AddRoundKeyOutput[25]), 
        .ZN(Red_SignaltoCheck[19]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_6_LFInst_1_U3  ( .A(AddRoundKeyOutput[27]), 
        .B(AddRoundKeyOutput[24]), .ZN(\Red_ToCheckInst_LFInst_6_LFInst_1_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_6_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_6_LFInst_2_n2 ), .B(AddRoundKeyOutput[26]), 
        .ZN(Red_SignaltoCheck[20]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_6_LFInst_2_U3  ( .A(AddRoundKeyOutput[27]), 
        .B(AddRoundKeyOutput[25]), .ZN(\Red_ToCheckInst_LFInst_6_LFInst_2_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_7_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_7_LFInst_0_n2 ), .B(AddRoundKeyOutput[29]), 
        .ZN(Red_SignaltoCheck[21]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_7_LFInst_0_U3  ( .A(AddRoundKeyOutput[30]), 
        .B(AddRoundKeyOutput[28]), .ZN(\Red_ToCheckInst_LFInst_7_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_7_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_7_LFInst_1_n2 ), .B(AddRoundKeyOutput[29]), 
        .ZN(Red_SignaltoCheck[22]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_7_LFInst_1_U3  ( .A(AddRoundKeyOutput[31]), 
        .B(AddRoundKeyOutput[28]), .ZN(\Red_ToCheckInst_LFInst_7_LFInst_1_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_7_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_7_LFInst_2_n2 ), .B(AddRoundKeyOutput[30]), 
        .ZN(Red_SignaltoCheck[23]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_7_LFInst_2_U3  ( .A(AddRoundKeyOutput[31]), 
        .B(AddRoundKeyOutput[29]), .ZN(\Red_ToCheckInst_LFInst_7_LFInst_2_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_8_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_8_LFInst_0_n2 ), .B(AddRoundKeyOutput[33]), 
        .ZN(Red_SignaltoCheck[24]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_8_LFInst_0_U3  ( .A(AddRoundKeyOutput[34]), 
        .B(AddRoundKeyOutput[32]), .ZN(\Red_ToCheckInst_LFInst_8_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_8_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_8_LFInst_1_n2 ), .B(AddRoundKeyOutput[33]), 
        .ZN(Red_SignaltoCheck[25]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_8_LFInst_1_U3  ( .A(AddRoundKeyOutput[35]), 
        .B(AddRoundKeyOutput[32]), .ZN(\Red_ToCheckInst_LFInst_8_LFInst_1_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_8_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_8_LFInst_2_n2 ), .B(AddRoundKeyOutput[34]), 
        .ZN(Red_SignaltoCheck[26]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_8_LFInst_2_U3  ( .A(AddRoundKeyOutput[35]), 
        .B(AddRoundKeyOutput[33]), .ZN(\Red_ToCheckInst_LFInst_8_LFInst_2_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_9_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_9_LFInst_0_n2 ), .B(AddRoundKeyOutput[37]), 
        .ZN(Red_SignaltoCheck[27]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_9_LFInst_0_U3  ( .A(AddRoundKeyOutput[38]), 
        .B(AddRoundKeyOutput[36]), .ZN(\Red_ToCheckInst_LFInst_9_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_9_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_9_LFInst_1_n2 ), .B(AddRoundKeyOutput[37]), 
        .ZN(Red_SignaltoCheck[28]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_9_LFInst_1_U3  ( .A(AddRoundKeyOutput[39]), 
        .B(AddRoundKeyOutput[36]), .ZN(\Red_ToCheckInst_LFInst_9_LFInst_1_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_9_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_9_LFInst_2_n2 ), .B(AddRoundKeyOutput[38]), 
        .ZN(Red_SignaltoCheck[29]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_9_LFInst_2_U3  ( .A(AddRoundKeyOutput[39]), 
        .B(AddRoundKeyOutput[37]), .ZN(\Red_ToCheckInst_LFInst_9_LFInst_2_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_10_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_10_LFInst_0_n2 ), .B(AddRoundKeyOutput[41]), 
        .ZN(Red_SignaltoCheck[30]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_10_LFInst_0_U3  ( .A(AddRoundKeyOutput[42]), 
        .B(AddRoundKeyOutput[40]), .ZN(\Red_ToCheckInst_LFInst_10_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_10_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_10_LFInst_1_n2 ), .B(AddRoundKeyOutput[41]), 
        .ZN(Red_SignaltoCheck[31]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_10_LFInst_1_U3  ( .A(AddRoundKeyOutput[43]), 
        .B(AddRoundKeyOutput[40]), .ZN(\Red_ToCheckInst_LFInst_10_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_10_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_10_LFInst_2_n2 ), .B(AddRoundKeyOutput[42]), 
        .ZN(Red_SignaltoCheck[32]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_10_LFInst_2_U3  ( .A(AddRoundKeyOutput[43]), 
        .B(AddRoundKeyOutput[41]), .ZN(\Red_ToCheckInst_LFInst_10_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_11_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_11_LFInst_0_n2 ), .B(AddRoundKeyOutput[45]), 
        .ZN(Red_SignaltoCheck[33]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_11_LFInst_0_U3  ( .A(AddRoundKeyOutput[46]), 
        .B(AddRoundKeyOutput[44]), .ZN(\Red_ToCheckInst_LFInst_11_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_11_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_11_LFInst_1_n2 ), .B(AddRoundKeyOutput[45]), 
        .ZN(Red_SignaltoCheck[34]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_11_LFInst_1_U3  ( .A(AddRoundKeyOutput[47]), 
        .B(AddRoundKeyOutput[44]), .ZN(\Red_ToCheckInst_LFInst_11_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_11_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_11_LFInst_2_n2 ), .B(AddRoundKeyOutput[46]), 
        .ZN(Red_SignaltoCheck[35]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_11_LFInst_2_U3  ( .A(AddRoundKeyOutput[47]), 
        .B(AddRoundKeyOutput[45]), .ZN(\Red_ToCheckInst_LFInst_11_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_12_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_12_LFInst_0_n2 ), .B(AddRoundKeyOutput[49]), 
        .ZN(Red_SignaltoCheck[36]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_12_LFInst_0_U3  ( .A(AddRoundKeyOutput[50]), 
        .B(AddRoundKeyOutput[48]), .ZN(\Red_ToCheckInst_LFInst_12_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_12_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_12_LFInst_1_n2 ), .B(AddRoundKeyOutput[49]), 
        .ZN(Red_SignaltoCheck[37]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_12_LFInst_1_U3  ( .A(AddRoundKeyOutput[51]), 
        .B(AddRoundKeyOutput[48]), .ZN(\Red_ToCheckInst_LFInst_12_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_12_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_12_LFInst_2_n2 ), .B(AddRoundKeyOutput[50]), 
        .ZN(Red_SignaltoCheck[38]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_12_LFInst_2_U3  ( .A(AddRoundKeyOutput[51]), 
        .B(AddRoundKeyOutput[49]), .ZN(\Red_ToCheckInst_LFInst_12_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_13_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_13_LFInst_0_n2 ), .B(AddRoundKeyOutput[53]), 
        .ZN(Red_SignaltoCheck[39]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_13_LFInst_0_U3  ( .A(AddRoundKeyOutput[54]), 
        .B(AddRoundKeyOutput[52]), .ZN(\Red_ToCheckInst_LFInst_13_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_13_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_13_LFInst_1_n2 ), .B(AddRoundKeyOutput[53]), 
        .ZN(Red_SignaltoCheck[40]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_13_LFInst_1_U3  ( .A(AddRoundKeyOutput[55]), 
        .B(AddRoundKeyOutput[52]), .ZN(\Red_ToCheckInst_LFInst_13_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_13_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_13_LFInst_2_n2 ), .B(AddRoundKeyOutput[54]), 
        .ZN(Red_SignaltoCheck[41]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_13_LFInst_2_U3  ( .A(AddRoundKeyOutput[55]), 
        .B(AddRoundKeyOutput[53]), .ZN(\Red_ToCheckInst_LFInst_13_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_14_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_14_LFInst_0_n2 ), .B(AddRoundKeyOutput[57]), 
        .ZN(Red_SignaltoCheck[42]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_14_LFInst_0_U3  ( .A(AddRoundKeyOutput[58]), 
        .B(AddRoundKeyOutput[56]), .ZN(\Red_ToCheckInst_LFInst_14_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_14_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_14_LFInst_1_n2 ), .B(AddRoundKeyOutput[57]), 
        .ZN(Red_SignaltoCheck[43]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_14_LFInst_1_U3  ( .A(AddRoundKeyOutput[59]), 
        .B(AddRoundKeyOutput[56]), .ZN(\Red_ToCheckInst_LFInst_14_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_14_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_14_LFInst_2_n2 ), .B(AddRoundKeyOutput[58]), 
        .ZN(Red_SignaltoCheck[44]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_14_LFInst_2_U3  ( .A(AddRoundKeyOutput[59]), 
        .B(AddRoundKeyOutput[57]), .ZN(\Red_ToCheckInst_LFInst_14_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_15_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_15_LFInst_0_n2 ), .B(AddRoundKeyOutput[61]), 
        .ZN(Red_SignaltoCheck[45]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_15_LFInst_0_U3  ( .A(AddRoundKeyOutput[62]), 
        .B(AddRoundKeyOutput[60]), .ZN(\Red_ToCheckInst_LFInst_15_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_15_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_15_LFInst_1_n2 ), .B(AddRoundKeyOutput[61]), 
        .ZN(Red_SignaltoCheck[46]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_15_LFInst_1_U3  ( .A(AddRoundKeyOutput[63]), 
        .B(AddRoundKeyOutput[60]), .ZN(\Red_ToCheckInst_LFInst_15_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_15_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_15_LFInst_2_n2 ), .B(AddRoundKeyOutput[62]), 
        .ZN(Red_SignaltoCheck[47]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_15_LFInst_2_U3  ( .A(AddRoundKeyOutput[63]), 
        .B(AddRoundKeyOutput[61]), .ZN(\Red_ToCheckInst_LFInst_15_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_16_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_16_LFInst_0_n2 ), .B(Ciphertext[1]), .ZN(
        Red_SignaltoCheck[48]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_16_LFInst_0_U3  ( .A(Ciphertext[2]), .B(
        Ciphertext[0]), .ZN(\Red_ToCheckInst_LFInst_16_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_16_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_16_LFInst_1_n2 ), .B(Ciphertext[1]), .ZN(
        Red_SignaltoCheck[49]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_16_LFInst_1_U3  ( .A(Ciphertext[3]), .B(
        Ciphertext[0]), .ZN(\Red_ToCheckInst_LFInst_16_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_16_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_16_LFInst_2_n2 ), .B(Ciphertext[2]), .ZN(
        Red_SignaltoCheck[50]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_16_LFInst_2_U3  ( .A(Ciphertext[3]), .B(
        Ciphertext[1]), .ZN(\Red_ToCheckInst_LFInst_16_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_17_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_17_LFInst_0_n2 ), .B(Ciphertext[5]), .ZN(
        Red_SignaltoCheck[51]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_17_LFInst_0_U3  ( .A(Ciphertext[6]), .B(
        Ciphertext[4]), .ZN(\Red_ToCheckInst_LFInst_17_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_17_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_17_LFInst_1_n2 ), .B(Ciphertext[5]), .ZN(
        Red_SignaltoCheck[52]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_17_LFInst_1_U3  ( .A(Ciphertext[7]), .B(
        Ciphertext[4]), .ZN(\Red_ToCheckInst_LFInst_17_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_17_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_17_LFInst_2_n2 ), .B(Ciphertext[6]), .ZN(
        Red_SignaltoCheck[53]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_17_LFInst_2_U3  ( .A(Ciphertext[7]), .B(
        Ciphertext[5]), .ZN(\Red_ToCheckInst_LFInst_17_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_18_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_18_LFInst_0_n2 ), .B(Ciphertext[9]), .ZN(
        Red_SignaltoCheck[54]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_18_LFInst_0_U3  ( .A(Ciphertext[10]), .B(
        Ciphertext[8]), .ZN(\Red_ToCheckInst_LFInst_18_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_18_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_18_LFInst_1_n2 ), .B(Ciphertext[9]), .ZN(
        Red_SignaltoCheck[55]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_18_LFInst_1_U3  ( .A(Ciphertext[11]), .B(
        Ciphertext[8]), .ZN(\Red_ToCheckInst_LFInst_18_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_18_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_18_LFInst_2_n2 ), .B(Ciphertext[10]), .ZN(
        Red_SignaltoCheck[56]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_18_LFInst_2_U3  ( .A(Ciphertext[11]), .B(
        Ciphertext[9]), .ZN(\Red_ToCheckInst_LFInst_18_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_19_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_19_LFInst_0_n2 ), .B(Ciphertext[13]), .ZN(
        Red_SignaltoCheck[57]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_19_LFInst_0_U3  ( .A(Ciphertext[14]), .B(
        Ciphertext[12]), .ZN(\Red_ToCheckInst_LFInst_19_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_19_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_19_LFInst_1_n2 ), .B(Ciphertext[13]), .ZN(
        Red_SignaltoCheck[58]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_19_LFInst_1_U3  ( .A(Ciphertext[15]), .B(
        Ciphertext[12]), .ZN(\Red_ToCheckInst_LFInst_19_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_19_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_19_LFInst_2_n2 ), .B(Ciphertext[14]), .ZN(
        Red_SignaltoCheck[59]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_19_LFInst_2_U3  ( .A(Ciphertext[15]), .B(
        Ciphertext[13]), .ZN(\Red_ToCheckInst_LFInst_19_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_20_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_20_LFInst_0_n2 ), .B(Ciphertext[17]), .ZN(
        Red_SignaltoCheck[60]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_20_LFInst_0_U3  ( .A(Ciphertext[18]), .B(
        Ciphertext[16]), .ZN(\Red_ToCheckInst_LFInst_20_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_20_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_20_LFInst_1_n2 ), .B(Ciphertext[17]), .ZN(
        Red_SignaltoCheck[61]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_20_LFInst_1_U3  ( .A(Ciphertext[19]), .B(
        Ciphertext[16]), .ZN(\Red_ToCheckInst_LFInst_20_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_20_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_20_LFInst_2_n2 ), .B(Ciphertext[18]), .ZN(
        Red_SignaltoCheck[62]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_20_LFInst_2_U3  ( .A(Ciphertext[19]), .B(
        Ciphertext[17]), .ZN(\Red_ToCheckInst_LFInst_20_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_21_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_21_LFInst_0_n2 ), .B(Ciphertext[21]), .ZN(
        Red_SignaltoCheck[63]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_21_LFInst_0_U3  ( .A(Ciphertext[22]), .B(
        Ciphertext[20]), .ZN(\Red_ToCheckInst_LFInst_21_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_21_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_21_LFInst_1_n2 ), .B(Ciphertext[21]), .ZN(
        Red_SignaltoCheck[64]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_21_LFInst_1_U3  ( .A(Ciphertext[23]), .B(
        Ciphertext[20]), .ZN(\Red_ToCheckInst_LFInst_21_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_21_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_21_LFInst_2_n2 ), .B(Ciphertext[22]), .ZN(
        Red_SignaltoCheck[65]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_21_LFInst_2_U3  ( .A(Ciphertext[23]), .B(
        Ciphertext[21]), .ZN(\Red_ToCheckInst_LFInst_21_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_22_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_22_LFInst_0_n2 ), .B(Ciphertext[25]), .ZN(
        Red_SignaltoCheck[66]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_22_LFInst_0_U3  ( .A(Ciphertext[26]), .B(
        Ciphertext[24]), .ZN(\Red_ToCheckInst_LFInst_22_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_22_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_22_LFInst_1_n2 ), .B(Ciphertext[25]), .ZN(
        Red_SignaltoCheck[67]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_22_LFInst_1_U3  ( .A(Ciphertext[27]), .B(
        Ciphertext[24]), .ZN(\Red_ToCheckInst_LFInst_22_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_22_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_22_LFInst_2_n2 ), .B(Ciphertext[26]), .ZN(
        Red_SignaltoCheck[68]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_22_LFInst_2_U3  ( .A(Ciphertext[27]), .B(
        Ciphertext[25]), .ZN(\Red_ToCheckInst_LFInst_22_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_23_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_23_LFInst_0_n2 ), .B(Ciphertext[29]), .ZN(
        Red_SignaltoCheck[69]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_23_LFInst_0_U3  ( .A(Ciphertext[30]), .B(
        Ciphertext[28]), .ZN(\Red_ToCheckInst_LFInst_23_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_23_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_23_LFInst_1_n2 ), .B(Ciphertext[29]), .ZN(
        Red_SignaltoCheck[70]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_23_LFInst_1_U3  ( .A(Ciphertext[31]), .B(
        Ciphertext[28]), .ZN(\Red_ToCheckInst_LFInst_23_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_23_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_23_LFInst_2_n2 ), .B(Ciphertext[30]), .ZN(
        Red_SignaltoCheck[71]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_23_LFInst_2_U3  ( .A(Ciphertext[31]), .B(
        Ciphertext[29]), .ZN(\Red_ToCheckInst_LFInst_23_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_24_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_24_LFInst_0_n2 ), .B(Ciphertext[33]), .ZN(
        Red_SignaltoCheck[72]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_24_LFInst_0_U3  ( .A(Ciphertext[34]), .B(
        Ciphertext[32]), .ZN(\Red_ToCheckInst_LFInst_24_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_24_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_24_LFInst_1_n2 ), .B(Ciphertext[33]), .ZN(
        Red_SignaltoCheck[73]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_24_LFInst_1_U3  ( .A(Ciphertext[35]), .B(
        Ciphertext[32]), .ZN(\Red_ToCheckInst_LFInst_24_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_24_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_24_LFInst_2_n2 ), .B(Ciphertext[34]), .ZN(
        Red_SignaltoCheck[74]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_24_LFInst_2_U3  ( .A(Ciphertext[35]), .B(
        Ciphertext[33]), .ZN(\Red_ToCheckInst_LFInst_24_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_25_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_25_LFInst_0_n2 ), .B(Ciphertext[37]), .ZN(
        Red_SignaltoCheck[75]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_25_LFInst_0_U3  ( .A(Ciphertext[38]), .B(
        Ciphertext[36]), .ZN(\Red_ToCheckInst_LFInst_25_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_25_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_25_LFInst_1_n2 ), .B(Ciphertext[37]), .ZN(
        Red_SignaltoCheck[76]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_25_LFInst_1_U3  ( .A(Ciphertext[39]), .B(
        Ciphertext[36]), .ZN(\Red_ToCheckInst_LFInst_25_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_25_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_25_LFInst_2_n2 ), .B(Ciphertext[38]), .ZN(
        Red_SignaltoCheck[77]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_25_LFInst_2_U3  ( .A(Ciphertext[39]), .B(
        Ciphertext[37]), .ZN(\Red_ToCheckInst_LFInst_25_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_26_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_26_LFInst_0_n2 ), .B(Ciphertext[41]), .ZN(
        Red_SignaltoCheck[78]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_26_LFInst_0_U3  ( .A(Ciphertext[42]), .B(
        Ciphertext[40]), .ZN(\Red_ToCheckInst_LFInst_26_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_26_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_26_LFInst_1_n2 ), .B(Ciphertext[41]), .ZN(
        Red_SignaltoCheck[79]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_26_LFInst_1_U3  ( .A(Ciphertext[43]), .B(
        Ciphertext[40]), .ZN(\Red_ToCheckInst_LFInst_26_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_26_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_26_LFInst_2_n2 ), .B(Ciphertext[42]), .ZN(
        Red_SignaltoCheck[80]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_26_LFInst_2_U3  ( .A(Ciphertext[43]), .B(
        Ciphertext[41]), .ZN(\Red_ToCheckInst_LFInst_26_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_27_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_27_LFInst_0_n2 ), .B(Ciphertext[45]), .ZN(
        Red_SignaltoCheck[81]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_27_LFInst_0_U3  ( .A(Ciphertext[46]), .B(
        Ciphertext[44]), .ZN(\Red_ToCheckInst_LFInst_27_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_27_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_27_LFInst_1_n2 ), .B(Ciphertext[45]), .ZN(
        Red_SignaltoCheck[82]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_27_LFInst_1_U3  ( .A(Ciphertext[47]), .B(
        Ciphertext[44]), .ZN(\Red_ToCheckInst_LFInst_27_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_27_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_27_LFInst_2_n2 ), .B(Ciphertext[46]), .ZN(
        Red_SignaltoCheck[83]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_27_LFInst_2_U3  ( .A(Ciphertext[47]), .B(
        Ciphertext[45]), .ZN(\Red_ToCheckInst_LFInst_27_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_28_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_28_LFInst_0_n2 ), .B(Ciphertext[49]), .ZN(
        Red_SignaltoCheck[84]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_28_LFInst_0_U3  ( .A(Ciphertext[50]), .B(
        Ciphertext[48]), .ZN(\Red_ToCheckInst_LFInst_28_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_28_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_28_LFInst_1_n2 ), .B(Ciphertext[49]), .ZN(
        Red_SignaltoCheck[85]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_28_LFInst_1_U3  ( .A(Ciphertext[51]), .B(
        Ciphertext[48]), .ZN(\Red_ToCheckInst_LFInst_28_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_28_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_28_LFInst_2_n2 ), .B(Ciphertext[50]), .ZN(
        Red_SignaltoCheck[86]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_28_LFInst_2_U3  ( .A(Ciphertext[51]), .B(
        Ciphertext[49]), .ZN(\Red_ToCheckInst_LFInst_28_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_29_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_29_LFInst_0_n2 ), .B(Ciphertext[53]), .ZN(
        Red_SignaltoCheck[87]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_29_LFInst_0_U3  ( .A(Ciphertext[54]), .B(
        Ciphertext[52]), .ZN(\Red_ToCheckInst_LFInst_29_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_29_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_29_LFInst_1_n2 ), .B(Ciphertext[53]), .ZN(
        Red_SignaltoCheck[88]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_29_LFInst_1_U3  ( .A(Ciphertext[55]), .B(
        Ciphertext[52]), .ZN(\Red_ToCheckInst_LFInst_29_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_29_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_29_LFInst_2_n2 ), .B(Ciphertext[54]), .ZN(
        Red_SignaltoCheck[89]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_29_LFInst_2_U3  ( .A(Ciphertext[55]), .B(
        Ciphertext[53]), .ZN(\Red_ToCheckInst_LFInst_29_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_30_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_30_LFInst_0_n2 ), .B(Ciphertext[57]), .ZN(
        Red_SignaltoCheck[90]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_30_LFInst_0_U3  ( .A(Ciphertext[58]), .B(
        Ciphertext[56]), .ZN(\Red_ToCheckInst_LFInst_30_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_30_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_30_LFInst_1_n2 ), .B(Ciphertext[57]), .ZN(
        Red_SignaltoCheck[91]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_30_LFInst_1_U3  ( .A(Ciphertext[59]), .B(
        Ciphertext[56]), .ZN(\Red_ToCheckInst_LFInst_30_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_30_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_30_LFInst_2_n2 ), .B(Ciphertext[58]), .ZN(
        Red_SignaltoCheck[92]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_30_LFInst_2_U3  ( .A(Ciphertext[59]), .B(
        Ciphertext[57]), .ZN(\Red_ToCheckInst_LFInst_30_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_31_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_31_LFInst_0_n2 ), .B(Ciphertext[61]), .ZN(
        Red_SignaltoCheck[93]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_31_LFInst_0_U3  ( .A(Ciphertext[62]), .B(
        Ciphertext[60]), .ZN(\Red_ToCheckInst_LFInst_31_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_31_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_31_LFInst_1_n2 ), .B(Ciphertext[61]), .ZN(
        Red_SignaltoCheck[94]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_31_LFInst_1_U3  ( .A(Ciphertext[63]), .B(
        Ciphertext[60]), .ZN(\Red_ToCheckInst_LFInst_31_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_31_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_31_LFInst_2_n2 ), .B(Ciphertext[62]), .ZN(
        Red_SignaltoCheck[95]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_31_LFInst_2_U3  ( .A(Ciphertext[63]), .B(
        Ciphertext[61]), .ZN(\Red_ToCheckInst_LFInst_31_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_32_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_32_LFInst_0_n2 ), .B(\Red_MCInst_MC3_v3_3 [2]), 
        .ZN(Red_SignaltoCheck[96]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_32_LFInst_0_U3  ( .A(\MCInst_MC3_v3_0 [3]), 
        .B(\MCInst_MC3_v3_2 [3]), .ZN(\Red_ToCheckInst_LFInst_32_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_32_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_32_LFInst_1_n2 ), .B(\Red_MCInst_MC3_v3_3 [2]), 
        .ZN(Red_SignaltoCheck[97]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_32_LFInst_1_U3  ( .A(
        \Red_MCInst_MC3_v3_1 [2]), .B(\MCInst_MC3_v3_2 [3]), .ZN(
        \Red_ToCheckInst_LFInst_32_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_32_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_32_LFInst_2_n2 ), .B(\MCInst_MC3_v3_0 [3]), 
        .ZN(Red_SignaltoCheck[98]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_32_LFInst_2_U3  ( .A(
        \Red_MCInst_MC3_v3_1 [2]), .B(\Red_MCInst_MC3_v3_3 [2]), .ZN(
        \Red_ToCheckInst_LFInst_32_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_33_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_33_LFInst_0_n2 ), .B(\Red_MCInst_MC2_v3_3 [2]), 
        .ZN(Red_SignaltoCheck[99]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_33_LFInst_0_U3  ( .A(\MCInst_MC2_v3_0 [3]), 
        .B(\MCInst_MC2_v3_2 [3]), .ZN(\Red_ToCheckInst_LFInst_33_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_33_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_33_LFInst_1_n2 ), .B(\Red_MCInst_MC2_v3_3 [2]), 
        .ZN(Red_SignaltoCheck[100]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_33_LFInst_1_U3  ( .A(
        \Red_MCInst_MC2_v3_1 [2]), .B(\MCInst_MC2_v3_2 [3]), .ZN(
        \Red_ToCheckInst_LFInst_33_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_33_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_33_LFInst_2_n2 ), .B(\MCInst_MC2_v3_0 [3]), 
        .ZN(Red_SignaltoCheck[101]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_33_LFInst_2_U3  ( .A(
        \Red_MCInst_MC2_v3_1 [2]), .B(\Red_MCInst_MC2_v3_3 [2]), .ZN(
        \Red_ToCheckInst_LFInst_33_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_34_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_34_LFInst_0_n2 ), .B(\Red_MCInst_MC1_v3_3 [2]), 
        .ZN(Red_SignaltoCheck[102]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_34_LFInst_0_U3  ( .A(\MCInst_MC1_v3_0 [3]), 
        .B(\MCInst_MC1_v3_2 [3]), .ZN(\Red_ToCheckInst_LFInst_34_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_34_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_34_LFInst_1_n2 ), .B(\Red_MCInst_MC1_v3_3 [2]), 
        .ZN(Red_SignaltoCheck[103]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_34_LFInst_1_U3  ( .A(
        \Red_MCInst_MC1_v3_1 [2]), .B(\MCInst_MC1_v3_2 [3]), .ZN(
        \Red_ToCheckInst_LFInst_34_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_34_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_34_LFInst_2_n2 ), .B(\MCInst_MC1_v3_0 [3]), 
        .ZN(Red_SignaltoCheck[104]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_34_LFInst_2_U3  ( .A(
        \Red_MCInst_MC1_v3_1 [2]), .B(\Red_MCInst_MC1_v3_3 [2]), .ZN(
        \Red_ToCheckInst_LFInst_34_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_35_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_35_LFInst_0_n2 ), .B(\Red_MCInst_MC0_v3_3 [2]), 
        .ZN(Red_SignaltoCheck[105]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_35_LFInst_0_U3  ( .A(\MCInst_MC0_v3_0 [3]), 
        .B(\MCInst_MC0_v3_2 [3]), .ZN(\Red_ToCheckInst_LFInst_35_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_35_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_35_LFInst_1_n2 ), .B(\Red_MCInst_MC0_v3_3 [2]), 
        .ZN(Red_SignaltoCheck[106]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_35_LFInst_1_U3  ( .A(
        \Red_MCInst_MC0_v3_1 [2]), .B(\MCInst_MC0_v3_2 [3]), .ZN(
        \Red_ToCheckInst_LFInst_35_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_35_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_35_LFInst_2_n2 ), .B(\MCInst_MC0_v3_0 [3]), 
        .ZN(Red_SignaltoCheck[107]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_35_LFInst_2_U3  ( .A(
        \Red_MCInst_MC0_v3_1 [2]), .B(\Red_MCInst_MC0_v3_3 [2]), .ZN(
        \Red_ToCheckInst_LFInst_35_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_36_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_36_LFInst_0_n2 ), .B(\MCInst_MC3_v2_0 [2]), 
        .ZN(Red_SignaltoCheck[108]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_36_LFInst_0_U3  ( .A(\MCInst_MC3_v2_0 [3]), 
        .B(\Red_MCInst_MC3_v2_1 [1]), .ZN(
        \Red_ToCheckInst_LFInst_36_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_36_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_36_LFInst_1_n2 ), .B(\MCInst_MC3_v2_0 [2]), 
        .ZN(Red_SignaltoCheck[109]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_36_LFInst_1_U3  ( .A(
        \Red_MCInst_MC3_v2_2 [1]), .B(\Red_MCInst_MC3_v2_1 [1]), .ZN(
        \Red_ToCheckInst_LFInst_36_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_36_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_36_LFInst_2_n2 ), .B(\MCInst_MC3_v2_0 [3]), 
        .ZN(Red_SignaltoCheck[110]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_36_LFInst_2_U3  ( .A(
        \Red_MCInst_MC3_v2_2 [1]), .B(\MCInst_MC3_v2_0 [2]), .ZN(
        \Red_ToCheckInst_LFInst_36_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_37_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_37_LFInst_0_n2 ), .B(\MCInst_MC2_v2_0 [2]), 
        .ZN(Red_SignaltoCheck[111]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_37_LFInst_0_U3  ( .A(\MCInst_MC2_v2_0 [3]), 
        .B(\Red_MCInst_MC2_v2_1 [1]), .ZN(
        \Red_ToCheckInst_LFInst_37_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_37_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_37_LFInst_1_n2 ), .B(\MCInst_MC2_v2_0 [2]), 
        .ZN(Red_SignaltoCheck[112]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_37_LFInst_1_U3  ( .A(
        \Red_MCInst_MC2_v2_2 [1]), .B(\Red_MCInst_MC2_v2_1 [1]), .ZN(
        \Red_ToCheckInst_LFInst_37_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_37_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_37_LFInst_2_n2 ), .B(\MCInst_MC2_v2_0 [3]), 
        .ZN(Red_SignaltoCheck[113]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_37_LFInst_2_U3  ( .A(
        \Red_MCInst_MC2_v2_2 [1]), .B(\MCInst_MC2_v2_0 [2]), .ZN(
        \Red_ToCheckInst_LFInst_37_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_38_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_38_LFInst_0_n2 ), .B(\MCInst_MC1_v2_0 [2]), 
        .ZN(Red_SignaltoCheck[114]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_38_LFInst_0_U3  ( .A(\MCInst_MC1_v2_0 [3]), 
        .B(\Red_MCInst_MC1_v2_1 [1]), .ZN(
        \Red_ToCheckInst_LFInst_38_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_38_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_38_LFInst_1_n2 ), .B(\MCInst_MC1_v2_0 [2]), 
        .ZN(Red_SignaltoCheck[115]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_38_LFInst_1_U3  ( .A(
        \Red_MCInst_MC1_v2_2 [1]), .B(\Red_MCInst_MC1_v2_1 [1]), .ZN(
        \Red_ToCheckInst_LFInst_38_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_38_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_38_LFInst_2_n2 ), .B(\MCInst_MC1_v2_0 [3]), 
        .ZN(Red_SignaltoCheck[116]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_38_LFInst_2_U3  ( .A(
        \Red_MCInst_MC1_v2_2 [1]), .B(\MCInst_MC1_v2_0 [2]), .ZN(
        \Red_ToCheckInst_LFInst_38_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_39_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_39_LFInst_0_n2 ), .B(\MCInst_MC0_v2_0 [2]), 
        .ZN(Red_SignaltoCheck[117]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_39_LFInst_0_U3  ( .A(\MCInst_MC0_v2_0 [3]), 
        .B(\Red_MCInst_MC0_v2_1 [1]), .ZN(
        \Red_ToCheckInst_LFInst_39_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_39_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_39_LFInst_1_n2 ), .B(\MCInst_MC0_v2_0 [2]), 
        .ZN(Red_SignaltoCheck[118]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_39_LFInst_1_U3  ( .A(
        \Red_MCInst_MC0_v2_2 [1]), .B(\Red_MCInst_MC0_v2_1 [1]), .ZN(
        \Red_ToCheckInst_LFInst_39_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_39_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_39_LFInst_2_n2 ), .B(\MCInst_MC0_v2_0 [3]), 
        .ZN(Red_SignaltoCheck[119]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_39_LFInst_2_U3  ( .A(
        \Red_MCInst_MC0_v2_2 [1]), .B(\MCInst_MC0_v2_0 [2]), .ZN(
        \Red_ToCheckInst_LFInst_39_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_40_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_40_LFInst_0_n2 ), .B(\Red_MCInst_MC3_v1_2 [1]), 
        .ZN(Red_SignaltoCheck[120]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_40_LFInst_0_U3  ( .A(\MCInst_MC3_v1_3 [3]), 
        .B(\MCInst_MC3_v1_0 [0]), .ZN(\Red_ToCheckInst_LFInst_40_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_40_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_40_LFInst_1_n2 ), .B(\Red_MCInst_MC3_v1_2 [1]), 
        .ZN(Red_SignaltoCheck[121]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_40_LFInst_1_U3  ( .A(
        \Red_MCInst_MC3_v1_1 [2]), .B(\MCInst_MC3_v1_0 [0]), .ZN(
        \Red_ToCheckInst_LFInst_40_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_40_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_40_LFInst_2_n2 ), .B(\MCInst_MC3_v1_3 [3]), 
        .ZN(Red_SignaltoCheck[122]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_40_LFInst_2_U3  ( .A(
        \Red_MCInst_MC3_v1_1 [2]), .B(\Red_MCInst_MC3_v1_2 [1]), .ZN(
        \Red_ToCheckInst_LFInst_40_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_41_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_41_LFInst_0_n2 ), .B(\Red_MCInst_MC2_v1_2 [1]), 
        .ZN(Red_SignaltoCheck[123]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_41_LFInst_0_U3  ( .A(\MCInst_MC2_v1_3 [3]), 
        .B(\MCInst_MC2_v1_0 [0]), .ZN(\Red_ToCheckInst_LFInst_41_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_41_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_41_LFInst_1_n2 ), .B(\Red_MCInst_MC2_v1_2 [1]), 
        .ZN(Red_SignaltoCheck[124]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_41_LFInst_1_U3  ( .A(
        \Red_MCInst_MC2_v1_1 [2]), .B(\MCInst_MC2_v1_0 [0]), .ZN(
        \Red_ToCheckInst_LFInst_41_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_41_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_41_LFInst_2_n2 ), .B(\MCInst_MC2_v1_3 [3]), 
        .ZN(Red_SignaltoCheck[125]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_41_LFInst_2_U3  ( .A(
        \Red_MCInst_MC2_v1_1 [2]), .B(\Red_MCInst_MC2_v1_2 [1]), .ZN(
        \Red_ToCheckInst_LFInst_41_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_42_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_42_LFInst_0_n2 ), .B(\Red_MCInst_MC1_v1_2 [1]), 
        .ZN(Red_SignaltoCheck[126]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_42_LFInst_0_U3  ( .A(\MCInst_MC1_v1_3 [3]), 
        .B(\MCInst_MC1_v1_0 [0]), .ZN(\Red_ToCheckInst_LFInst_42_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_42_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_42_LFInst_1_n2 ), .B(\Red_MCInst_MC1_v1_2 [1]), 
        .ZN(Red_SignaltoCheck[127]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_42_LFInst_1_U3  ( .A(
        \Red_MCInst_MC1_v1_1 [2]), .B(\MCInst_MC1_v1_0 [0]), .ZN(
        \Red_ToCheckInst_LFInst_42_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_42_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_42_LFInst_2_n2 ), .B(\MCInst_MC1_v1_3 [3]), 
        .ZN(Red_SignaltoCheck[128]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_42_LFInst_2_U3  ( .A(
        \Red_MCInst_MC1_v1_1 [2]), .B(\Red_MCInst_MC1_v1_2 [1]), .ZN(
        \Red_ToCheckInst_LFInst_42_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_43_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_43_LFInst_0_n2 ), .B(\Red_MCInst_MC0_v1_2 [1]), 
        .ZN(Red_SignaltoCheck[129]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_43_LFInst_0_U3  ( .A(\MCInst_MC0_v1_3 [3]), 
        .B(\MCInst_MC0_v1_0 [0]), .ZN(\Red_ToCheckInst_LFInst_43_LFInst_0_n2 )
         );
  XNOR2_X1 \Red_ToCheckInst_LFInst_43_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_43_LFInst_1_n2 ), .B(\Red_MCInst_MC0_v1_2 [1]), 
        .ZN(Red_SignaltoCheck[130]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_43_LFInst_1_U3  ( .A(
        \Red_MCInst_MC0_v1_1 [2]), .B(\MCInst_MC0_v1_0 [0]), .ZN(
        \Red_ToCheckInst_LFInst_43_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_43_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_43_LFInst_2_n2 ), .B(\MCInst_MC0_v1_3 [3]), 
        .ZN(Red_SignaltoCheck[131]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_43_LFInst_2_U3  ( .A(
        \Red_MCInst_MC0_v1_1 [2]), .B(\Red_MCInst_MC0_v1_2 [1]), .ZN(
        \Red_ToCheckInst_LFInst_43_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_44_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_44_LFInst_0_n2 ), .B(\Red_MCInst_MC3_v0_2 [2]), 
        .ZN(Red_SignaltoCheck[132]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_44_LFInst_0_U3  ( .A(\MCInst_MC3_v0_3 [3]), 
        .B(\Red_MCInst_MC3_v0_0 [0]), .ZN(
        \Red_ToCheckInst_LFInst_44_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_44_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_44_LFInst_1_n2 ), .B(\Red_MCInst_MC3_v0_2 [2]), 
        .ZN(Red_SignaltoCheck[133]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_44_LFInst_1_U3  ( .A(
        \Red_MCInst_MC3_v0_1 [0]), .B(\Red_MCInst_MC3_v0_0 [0]), .ZN(
        \Red_ToCheckInst_LFInst_44_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_44_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_44_LFInst_2_n2 ), .B(\MCInst_MC3_v0_3 [3]), 
        .ZN(Red_SignaltoCheck[134]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_44_LFInst_2_U3  ( .A(
        \Red_MCInst_MC3_v0_1 [0]), .B(\Red_MCInst_MC3_v0_2 [2]), .ZN(
        \Red_ToCheckInst_LFInst_44_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_45_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_45_LFInst_0_n2 ), .B(\Red_MCInst_MC2_v0_2 [2]), 
        .ZN(Red_SignaltoCheck[135]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_45_LFInst_0_U3  ( .A(\MCInst_MC2_v0_3 [3]), 
        .B(\Red_MCInst_MC2_v0_0 [0]), .ZN(
        \Red_ToCheckInst_LFInst_45_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_45_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_45_LFInst_1_n2 ), .B(\Red_MCInst_MC2_v0_2 [2]), 
        .ZN(Red_SignaltoCheck[136]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_45_LFInst_1_U3  ( .A(
        \Red_MCInst_MC2_v0_1 [0]), .B(\Red_MCInst_MC2_v0_0 [0]), .ZN(
        \Red_ToCheckInst_LFInst_45_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_45_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_45_LFInst_2_n2 ), .B(\MCInst_MC2_v0_3 [3]), 
        .ZN(Red_SignaltoCheck[137]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_45_LFInst_2_U3  ( .A(
        \Red_MCInst_MC2_v0_1 [0]), .B(\Red_MCInst_MC2_v0_2 [2]), .ZN(
        \Red_ToCheckInst_LFInst_45_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_46_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_46_LFInst_0_n2 ), .B(\Red_MCInst_MC1_v0_2 [2]), 
        .ZN(Red_SignaltoCheck[138]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_46_LFInst_0_U3  ( .A(\MCInst_MC1_v0_3 [3]), 
        .B(\Red_MCInst_MC1_v0_0 [0]), .ZN(
        \Red_ToCheckInst_LFInst_46_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_46_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_46_LFInst_1_n2 ), .B(\Red_MCInst_MC1_v0_2 [2]), 
        .ZN(Red_SignaltoCheck[139]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_46_LFInst_1_U3  ( .A(
        \Red_MCInst_MC1_v0_1 [0]), .B(\Red_MCInst_MC1_v0_0 [0]), .ZN(
        \Red_ToCheckInst_LFInst_46_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_46_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_46_LFInst_2_n2 ), .B(\MCInst_MC1_v0_3 [3]), 
        .ZN(Red_SignaltoCheck[140]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_46_LFInst_2_U3  ( .A(
        \Red_MCInst_MC1_v0_1 [0]), .B(\Red_MCInst_MC1_v0_2 [2]), .ZN(
        \Red_ToCheckInst_LFInst_46_LFInst_2_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_47_LFInst_0_U4  ( .A(
        \Red_ToCheckInst_LFInst_47_LFInst_0_n2 ), .B(\Red_MCInst_MC0_v0_2 [2]), 
        .ZN(Red_SignaltoCheck[141]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_47_LFInst_0_U3  ( .A(\MCInst_MC0_v0_3 [3]), 
        .B(\Red_MCInst_MC0_v0_0 [0]), .ZN(
        \Red_ToCheckInst_LFInst_47_LFInst_0_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_47_LFInst_1_U4  ( .A(
        \Red_ToCheckInst_LFInst_47_LFInst_1_n2 ), .B(\Red_MCInst_MC0_v0_2 [2]), 
        .ZN(Red_SignaltoCheck[142]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_47_LFInst_1_U3  ( .A(
        \Red_MCInst_MC0_v0_1 [0]), .B(\Red_MCInst_MC0_v0_0 [0]), .ZN(
        \Red_ToCheckInst_LFInst_47_LFInst_1_n2 ) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_47_LFInst_2_U4  ( .A(
        \Red_ToCheckInst_LFInst_47_LFInst_2_n2 ), .B(\MCInst_MC0_v0_3 [3]), 
        .ZN(Red_SignaltoCheck[143]) );
  XNOR2_X1 \Red_ToCheckInst_LFInst_47_LFInst_2_U3  ( .A(
        \Red_MCInst_MC0_v0_1 [0]), .B(\Red_MCInst_MC0_v0_2 [2]), .ZN(
        \Red_ToCheckInst_LFInst_47_LFInst_2_n2 ) );
  NOR2_X1 \Check1_CheckInst_0_U79  ( .A1(\Check1_CheckInst_0_n95 ), .A2(
        \Check1_CheckInst_0_n94 ), .ZN(Error[0]) );
  NAND2_X1 \Check1_CheckInst_0_U78  ( .A1(\Check1_CheckInst_0_n93 ), .A2(
        \Check1_CheckInst_0_n92 ), .ZN(\Check1_CheckInst_0_n94 ) );
  NOR2_X1 \Check1_CheckInst_0_U77  ( .A1(\Check1_CheckInst_0_n91 ), .A2(
        \Check1_CheckInst_0_n90 ), .ZN(\Check1_CheckInst_0_n92 ) );
  NAND2_X1 \Check1_CheckInst_0_U76  ( .A1(\Check1_CheckInst_0_n89 ), .A2(
        \Check1_CheckInst_0_n88 ), .ZN(\Check1_CheckInst_0_n90 ) );
  NOR2_X1 \Check1_CheckInst_0_U75  ( .A1(\Check1_CheckInst_0_n87 ), .A2(
        \Check1_CheckInst_0_n86 ), .ZN(\Check1_CheckInst_0_n88 ) );
  NAND2_X1 \Check1_CheckInst_0_U74  ( .A1(\Check1_CheckInst_0_n85 ), .A2(
        \Check1_CheckInst_0_n84 ), .ZN(\Check1_CheckInst_0_n86 ) );
  NOR2_X1 \Check1_CheckInst_0_U73  ( .A1(\Check1_CheckInst_0_n83 ), .A2(
        \Check1_CheckInst_0_n82 ), .ZN(\Check1_CheckInst_0_n84 ) );
  NAND2_X1 \Check1_CheckInst_0_U72  ( .A1(\Check1_CheckInst_0_n81 ), .A2(
        \Check1_CheckInst_0_n80 ), .ZN(\Check1_CheckInst_0_n82 ) );
  XNOR2_X1 \Check1_CheckInst_0_U71  ( .A(Red_AddRoundKeyOutput[24]), .B(
        Red_SignaltoCheck[24]), .ZN(\Check1_CheckInst_0_n80 ) );
  XNOR2_X1 \Check1_CheckInst_0_U70  ( .A(Red_AddRoundKeyOutput[0]), .B(
        Red_SignaltoCheck[0]), .ZN(\Check1_CheckInst_0_n81 ) );
  NAND2_X1 \Check1_CheckInst_0_U69  ( .A1(\Check1_CheckInst_0_n79 ), .A2(
        \Check1_CheckInst_0_n78 ), .ZN(\Check1_CheckInst_0_n83 ) );
  XNOR2_X1 \Check1_CheckInst_0_U68  ( .A(Red_AddRoundKeyOutput[30]), .B(
        Red_SignaltoCheck[30]), .ZN(\Check1_CheckInst_0_n78 ) );
  XNOR2_X1 \Check1_CheckInst_0_U67  ( .A(Red_SignaltoCheck[3]), .B(
        Red_AddRoundKeyOutput[3]), .ZN(\Check1_CheckInst_0_n79 ) );
  NOR2_X1 \Check1_CheckInst_0_U66  ( .A1(\Check1_CheckInst_0_n77 ), .A2(
        \Check1_CheckInst_0_n76 ), .ZN(\Check1_CheckInst_0_n85 ) );
  NAND2_X1 \Check1_CheckInst_0_U65  ( .A1(\Check1_CheckInst_0_n75 ), .A2(
        \Check1_CheckInst_0_n74 ), .ZN(\Check1_CheckInst_0_n76 ) );
  NOR2_X1 \Check1_CheckInst_0_U64  ( .A1(Red_SignaltoCheck[135]), .A2(
        Red_SignaltoCheck[141]), .ZN(\Check1_CheckInst_0_n74 ) );
  NOR2_X1 \Check1_CheckInst_0_U63  ( .A1(Red_SignaltoCheck[126]), .A2(
        Red_SignaltoCheck[120]), .ZN(\Check1_CheckInst_0_n75 ) );
  NAND2_X1 \Check1_CheckInst_0_U62  ( .A1(\Check1_CheckInst_0_n73 ), .A2(
        \Check1_CheckInst_0_n72 ), .ZN(\Check1_CheckInst_0_n77 ) );
  NOR2_X1 \Check1_CheckInst_0_U61  ( .A1(Red_SignaltoCheck[138]), .A2(
        Red_SignaltoCheck[102]), .ZN(\Check1_CheckInst_0_n72 ) );
  NOR2_X1 \Check1_CheckInst_0_U60  ( .A1(Red_SignaltoCheck[129]), .A2(
        Red_SignaltoCheck[111]), .ZN(\Check1_CheckInst_0_n73 ) );
  NAND2_X1 \Check1_CheckInst_0_U59  ( .A1(\Check1_CheckInst_0_n71 ), .A2(
        \Check1_CheckInst_0_n70 ), .ZN(\Check1_CheckInst_0_n87 ) );
  NOR2_X1 \Check1_CheckInst_0_U58  ( .A1(\Check1_CheckInst_0_n69 ), .A2(
        \Check1_CheckInst_0_n68 ), .ZN(\Check1_CheckInst_0_n70 ) );
  XOR2_X1 \Check1_CheckInst_0_U57  ( .A(Red_AddRoundKeyOutput[18]), .B(
        Red_SignaltoCheck[18]), .Z(\Check1_CheckInst_0_n68 ) );
  XOR2_X1 \Check1_CheckInst_0_U56  ( .A(Red_AddRoundKeyOutput[15]), .B(
        Red_SignaltoCheck[15]), .Z(\Check1_CheckInst_0_n69 ) );
  NOR2_X1 \Check1_CheckInst_0_U55  ( .A1(\Check1_CheckInst_0_n67 ), .A2(
        \Check1_CheckInst_0_n66 ), .ZN(\Check1_CheckInst_0_n71 ) );
  XOR2_X1 \Check1_CheckInst_0_U54  ( .A(Red_AddRoundKeyOutput[27]), .B(
        Red_SignaltoCheck[27]), .Z(\Check1_CheckInst_0_n66 ) );
  XOR2_X1 \Check1_CheckInst_0_U53  ( .A(Red_AddRoundKeyOutput[21]), .B(
        Red_SignaltoCheck[21]), .Z(\Check1_CheckInst_0_n67 ) );
  NOR2_X1 \Check1_CheckInst_0_U52  ( .A1(\Check1_CheckInst_0_n65 ), .A2(
        \Check1_CheckInst_0_n64 ), .ZN(\Check1_CheckInst_0_n89 ) );
  NAND2_X1 \Check1_CheckInst_0_U51  ( .A1(\Check1_CheckInst_0_n63 ), .A2(
        \Check1_CheckInst_0_n62 ), .ZN(\Check1_CheckInst_0_n64 ) );
  NOR2_X1 \Check1_CheckInst_0_U50  ( .A1(Red_SignaltoCheck[99]), .A2(
        Red_SignaltoCheck[117]), .ZN(\Check1_CheckInst_0_n62 ) );
  NOR2_X1 \Check1_CheckInst_0_U49  ( .A1(Red_SignaltoCheck[105]), .A2(
        Red_SignaltoCheck[96]), .ZN(\Check1_CheckInst_0_n63 ) );
  NAND2_X1 \Check1_CheckInst_0_U48  ( .A1(\Check1_CheckInst_0_n61 ), .A2(
        \Check1_CheckInst_0_n60 ), .ZN(\Check1_CheckInst_0_n65 ) );
  NOR2_X1 \Check1_CheckInst_0_U47  ( .A1(Red_SignaltoCheck[132]), .A2(
        Red_SignaltoCheck[123]), .ZN(\Check1_CheckInst_0_n60 ) );
  NOR2_X1 \Check1_CheckInst_0_U46  ( .A1(Red_SignaltoCheck[108]), .A2(
        Red_SignaltoCheck[114]), .ZN(\Check1_CheckInst_0_n61 ) );
  NAND2_X1 \Check1_CheckInst_0_U45  ( .A1(\Check1_CheckInst_0_n59 ), .A2(
        \Check1_CheckInst_0_n58 ), .ZN(\Check1_CheckInst_0_n91 ) );
  NOR2_X1 \Check1_CheckInst_0_U44  ( .A1(\Check1_CheckInst_0_n57 ), .A2(
        \Check1_CheckInst_0_n56 ), .ZN(\Check1_CheckInst_0_n58 ) );
  NAND2_X1 \Check1_CheckInst_0_U43  ( .A1(\Check1_CheckInst_0_n55 ), .A2(
        \Check1_CheckInst_0_n54 ), .ZN(\Check1_CheckInst_0_n56 ) );
  NOR2_X1 \Check1_CheckInst_0_U42  ( .A1(\Check1_CheckInst_0_n53 ), .A2(
        \Check1_CheckInst_0_n52 ), .ZN(\Check1_CheckInst_0_n54 ) );
  XOR2_X1 \Check1_CheckInst_0_U41  ( .A(Red_Feedback[30]), .B(
        Red_SignaltoCheck[78]), .Z(\Check1_CheckInst_0_n52 ) );
  XOR2_X1 \Check1_CheckInst_0_U40  ( .A(Red_Feedback[33]), .B(
        Red_SignaltoCheck[81]), .Z(\Check1_CheckInst_0_n53 ) );
  NOR2_X1 \Check1_CheckInst_0_U39  ( .A1(\Check1_CheckInst_0_n51 ), .A2(
        \Check1_CheckInst_0_n50 ), .ZN(\Check1_CheckInst_0_n55 ) );
  XOR2_X1 \Check1_CheckInst_0_U38  ( .A(Red_Feedback[24]), .B(
        Red_SignaltoCheck[72]), .Z(\Check1_CheckInst_0_n50 ) );
  XOR2_X1 \Check1_CheckInst_0_U37  ( .A(Red_Feedback[36]), .B(
        Red_SignaltoCheck[84]), .Z(\Check1_CheckInst_0_n51 ) );
  NAND2_X1 \Check1_CheckInst_0_U36  ( .A1(\Check1_CheckInst_0_n49 ), .A2(
        \Check1_CheckInst_0_n48 ), .ZN(\Check1_CheckInst_0_n57 ) );
  XNOR2_X1 \Check1_CheckInst_0_U35  ( .A(Red_Feedback[27]), .B(
        Red_SignaltoCheck[75]), .ZN(\Check1_CheckInst_0_n48 ) );
  XNOR2_X1 \Check1_CheckInst_0_U34  ( .A(Red_Feedback[21]), .B(
        Red_SignaltoCheck[69]), .ZN(\Check1_CheckInst_0_n49 ) );
  NOR2_X1 \Check1_CheckInst_0_U33  ( .A1(\Check1_CheckInst_0_n47 ), .A2(
        \Check1_CheckInst_0_n46 ), .ZN(\Check1_CheckInst_0_n59 ) );
  XOR2_X1 \Check1_CheckInst_0_U32  ( .A(Red_Feedback[39]), .B(
        Red_SignaltoCheck[87]), .Z(\Check1_CheckInst_0_n46 ) );
  XOR2_X1 \Check1_CheckInst_0_U31  ( .A(Red_Feedback[42]), .B(
        Red_SignaltoCheck[90]), .Z(\Check1_CheckInst_0_n47 ) );
  NOR2_X1 \Check1_CheckInst_0_U30  ( .A1(\Check1_CheckInst_0_n45 ), .A2(
        \Check1_CheckInst_0_n44 ), .ZN(\Check1_CheckInst_0_n93 ) );
  NAND2_X1 \Check1_CheckInst_0_U29  ( .A1(\Check1_CheckInst_0_n43 ), .A2(
        \Check1_CheckInst_0_n42 ), .ZN(\Check1_CheckInst_0_n44 ) );
  NOR2_X1 \Check1_CheckInst_0_U28  ( .A1(\Check1_CheckInst_0_n41 ), .A2(
        \Check1_CheckInst_0_n40 ), .ZN(\Check1_CheckInst_0_n42 ) );
  NAND2_X1 \Check1_CheckInst_0_U27  ( .A1(\Check1_CheckInst_0_n39 ), .A2(
        \Check1_CheckInst_0_n38 ), .ZN(\Check1_CheckInst_0_n40 ) );
  XNOR2_X1 \Check1_CheckInst_0_U26  ( .A(Red_AddRoundKeyOutput[45]), .B(
        Red_SignaltoCheck[45]), .ZN(\Check1_CheckInst_0_n38 ) );
  XNOR2_X1 \Check1_CheckInst_0_U25  ( .A(Red_Feedback[45]), .B(
        Red_SignaltoCheck[93]), .ZN(\Check1_CheckInst_0_n39 ) );
  NAND2_X1 \Check1_CheckInst_0_U24  ( .A1(\Check1_CheckInst_0_n37 ), .A2(
        \Check1_CheckInst_0_n36 ), .ZN(\Check1_CheckInst_0_n41 ) );
  XNOR2_X1 \Check1_CheckInst_0_U23  ( .A(Red_Feedback[0]), .B(
        Red_SignaltoCheck[48]), .ZN(\Check1_CheckInst_0_n36 ) );
  XNOR2_X1 \Check1_CheckInst_0_U22  ( .A(Red_AddRoundKeyOutput[42]), .B(
        Red_SignaltoCheck[42]), .ZN(\Check1_CheckInst_0_n37 ) );
  NOR2_X1 \Check1_CheckInst_0_U21  ( .A1(\Check1_CheckInst_0_n35 ), .A2(
        \Check1_CheckInst_0_n34 ), .ZN(\Check1_CheckInst_0_n43 ) );
  XOR2_X1 \Check1_CheckInst_0_U20  ( .A(Red_AddRoundKeyOutput[33]), .B(
        Red_SignaltoCheck[33]), .Z(\Check1_CheckInst_0_n34 ) );
  XOR2_X1 \Check1_CheckInst_0_U19  ( .A(Red_AddRoundKeyOutput[36]), .B(
        Red_SignaltoCheck[36]), .Z(\Check1_CheckInst_0_n35 ) );
  NAND2_X1 \Check1_CheckInst_0_U18  ( .A1(\Check1_CheckInst_0_n33 ), .A2(
        \Check1_CheckInst_0_n32 ), .ZN(\Check1_CheckInst_0_n45 ) );
  XNOR2_X1 \Check1_CheckInst_0_U17  ( .A(Red_Feedback[15]), .B(
        Red_SignaltoCheck[63]), .ZN(\Check1_CheckInst_0_n32 ) );
  XNOR2_X1 \Check1_CheckInst_0_U16  ( .A(Red_AddRoundKeyOutput[39]), .B(
        Red_SignaltoCheck[39]), .ZN(\Check1_CheckInst_0_n33 ) );
  NAND2_X1 \Check1_CheckInst_0_U15  ( .A1(\Check1_CheckInst_0_n31 ), .A2(
        \Check1_CheckInst_0_n30 ), .ZN(\Check1_CheckInst_0_n95 ) );
  NOR2_X1 \Check1_CheckInst_0_U14  ( .A1(\Check1_CheckInst_0_n29 ), .A2(
        \Check1_CheckInst_0_n28 ), .ZN(\Check1_CheckInst_0_n30 ) );
  NAND2_X1 \Check1_CheckInst_0_U13  ( .A1(\Check1_CheckInst_0_n27 ), .A2(
        \Check1_CheckInst_0_n26 ), .ZN(\Check1_CheckInst_0_n28 ) );
  NOR2_X1 \Check1_CheckInst_0_U12  ( .A1(\Check1_CheckInst_0_n25 ), .A2(
        \Check1_CheckInst_0_n24 ), .ZN(\Check1_CheckInst_0_n26 ) );
  XOR2_X1 \Check1_CheckInst_0_U11  ( .A(Red_Feedback[18]), .B(
        Red_SignaltoCheck[66]), .Z(\Check1_CheckInst_0_n24 ) );
  XOR2_X1 \Check1_CheckInst_0_U10  ( .A(Red_Feedback[12]), .B(
        Red_SignaltoCheck[60]), .Z(\Check1_CheckInst_0_n25 ) );
  NOR2_X1 \Check1_CheckInst_0_U9  ( .A1(\Check1_CheckInst_0_n23 ), .A2(
        \Check1_CheckInst_0_n22 ), .ZN(\Check1_CheckInst_0_n27 ) );
  XOR2_X1 \Check1_CheckInst_0_U8  ( .A(Red_Feedback[3]), .B(
        Red_SignaltoCheck[51]), .Z(\Check1_CheckInst_0_n22 ) );
  XOR2_X1 \Check1_CheckInst_0_U7  ( .A(Red_Feedback[6]), .B(
        Red_SignaltoCheck[54]), .Z(\Check1_CheckInst_0_n23 ) );
  NAND2_X1 \Check1_CheckInst_0_U6  ( .A1(\Check1_CheckInst_0_n21 ), .A2(
        \Check1_CheckInst_0_n20 ), .ZN(\Check1_CheckInst_0_n29 ) );
  XNOR2_X1 \Check1_CheckInst_0_U5  ( .A(Red_AddRoundKeyOutput[9]), .B(
        Red_SignaltoCheck[9]), .ZN(\Check1_CheckInst_0_n20 ) );
  XNOR2_X1 \Check1_CheckInst_0_U4  ( .A(Red_Feedback[9]), .B(
        Red_SignaltoCheck[57]), .ZN(\Check1_CheckInst_0_n21 ) );
  NOR2_X1 \Check1_CheckInst_0_U3  ( .A1(\Check1_CheckInst_0_n19 ), .A2(
        \Check1_CheckInst_0_n18 ), .ZN(\Check1_CheckInst_0_n31 ) );
  XOR2_X1 \Check1_CheckInst_0_U2  ( .A(Red_AddRoundKeyOutput[12]), .B(
        Red_SignaltoCheck[12]), .Z(\Check1_CheckInst_0_n18 ) );
  XOR2_X1 \Check1_CheckInst_0_U1  ( .A(Red_AddRoundKeyOutput[6]), .B(
        Red_SignaltoCheck[6]), .Z(\Check1_CheckInst_0_n19 ) );
  NOR2_X1 \Check1_CheckInst_1_U79  ( .A1(\Check1_CheckInst_1_n96 ), .A2(
        \Check1_CheckInst_1_n95 ), .ZN(Error[1]) );
  NAND2_X1 \Check1_CheckInst_1_U78  ( .A1(\Check1_CheckInst_1_n94 ), .A2(
        \Check1_CheckInst_1_n93 ), .ZN(\Check1_CheckInst_1_n95 ) );
  NOR2_X1 \Check1_CheckInst_1_U77  ( .A1(\Check1_CheckInst_1_n92 ), .A2(
        \Check1_CheckInst_1_n91 ), .ZN(\Check1_CheckInst_1_n93 ) );
  NAND2_X1 \Check1_CheckInst_1_U76  ( .A1(\Check1_CheckInst_1_n90 ), .A2(
        \Check1_CheckInst_1_n89 ), .ZN(\Check1_CheckInst_1_n91 ) );
  NOR2_X1 \Check1_CheckInst_1_U75  ( .A1(\Check1_CheckInst_1_n88 ), .A2(
        \Check1_CheckInst_1_n87 ), .ZN(\Check1_CheckInst_1_n89 ) );
  NAND2_X1 \Check1_CheckInst_1_U74  ( .A1(\Check1_CheckInst_1_n86 ), .A2(
        \Check1_CheckInst_1_n85 ), .ZN(\Check1_CheckInst_1_n87 ) );
  NOR2_X1 \Check1_CheckInst_1_U73  ( .A1(\Check1_CheckInst_1_n84 ), .A2(
        \Check1_CheckInst_1_n83 ), .ZN(\Check1_CheckInst_1_n85 ) );
  NAND2_X1 \Check1_CheckInst_1_U72  ( .A1(\Check1_CheckInst_1_n82 ), .A2(
        \Check1_CheckInst_1_n81 ), .ZN(\Check1_CheckInst_1_n83 ) );
  XNOR2_X1 \Check1_CheckInst_1_U71  ( .A(Red_AddRoundKeyOutput[25]), .B(
        Red_SignaltoCheck[25]), .ZN(\Check1_CheckInst_1_n81 ) );
  XNOR2_X1 \Check1_CheckInst_1_U70  ( .A(Red_AddRoundKeyOutput[1]), .B(
        Red_SignaltoCheck[1]), .ZN(\Check1_CheckInst_1_n82 ) );
  NAND2_X1 \Check1_CheckInst_1_U69  ( .A1(\Check1_CheckInst_1_n80 ), .A2(
        \Check1_CheckInst_1_n79 ), .ZN(\Check1_CheckInst_1_n84 ) );
  XNOR2_X1 \Check1_CheckInst_1_U68  ( .A(Red_AddRoundKeyOutput[31]), .B(
        Red_SignaltoCheck[31]), .ZN(\Check1_CheckInst_1_n79 ) );
  XNOR2_X1 \Check1_CheckInst_1_U67  ( .A(Red_SignaltoCheck[4]), .B(
        Red_AddRoundKeyOutput[4]), .ZN(\Check1_CheckInst_1_n80 ) );
  NOR2_X1 \Check1_CheckInst_1_U66  ( .A1(\Check1_CheckInst_1_n78 ), .A2(
        \Check1_CheckInst_1_n77 ), .ZN(\Check1_CheckInst_1_n86 ) );
  NAND2_X1 \Check1_CheckInst_1_U65  ( .A1(\Check1_CheckInst_1_n76 ), .A2(
        \Check1_CheckInst_1_n75 ), .ZN(\Check1_CheckInst_1_n77 ) );
  NOR2_X1 \Check1_CheckInst_1_U64  ( .A1(Red_SignaltoCheck[136]), .A2(
        Red_SignaltoCheck[142]), .ZN(\Check1_CheckInst_1_n75 ) );
  NOR2_X1 \Check1_CheckInst_1_U63  ( .A1(Red_SignaltoCheck[127]), .A2(
        Red_SignaltoCheck[121]), .ZN(\Check1_CheckInst_1_n76 ) );
  NAND2_X1 \Check1_CheckInst_1_U62  ( .A1(\Check1_CheckInst_1_n74 ), .A2(
        \Check1_CheckInst_1_n73 ), .ZN(\Check1_CheckInst_1_n78 ) );
  NOR2_X1 \Check1_CheckInst_1_U61  ( .A1(Red_SignaltoCheck[139]), .A2(
        Red_SignaltoCheck[103]), .ZN(\Check1_CheckInst_1_n73 ) );
  NOR2_X1 \Check1_CheckInst_1_U60  ( .A1(Red_SignaltoCheck[130]), .A2(
        Red_SignaltoCheck[112]), .ZN(\Check1_CheckInst_1_n74 ) );
  NAND2_X1 \Check1_CheckInst_1_U59  ( .A1(\Check1_CheckInst_1_n72 ), .A2(
        \Check1_CheckInst_1_n71 ), .ZN(\Check1_CheckInst_1_n88 ) );
  NOR2_X1 \Check1_CheckInst_1_U58  ( .A1(\Check1_CheckInst_1_n70 ), .A2(
        \Check1_CheckInst_1_n69 ), .ZN(\Check1_CheckInst_1_n71 ) );
  XOR2_X1 \Check1_CheckInst_1_U57  ( .A(Red_AddRoundKeyOutput[19]), .B(
        Red_SignaltoCheck[19]), .Z(\Check1_CheckInst_1_n69 ) );
  XOR2_X1 \Check1_CheckInst_1_U56  ( .A(Red_AddRoundKeyOutput[16]), .B(
        Red_SignaltoCheck[16]), .Z(\Check1_CheckInst_1_n70 ) );
  NOR2_X1 \Check1_CheckInst_1_U55  ( .A1(\Check1_CheckInst_1_n68 ), .A2(
        \Check1_CheckInst_1_n67 ), .ZN(\Check1_CheckInst_1_n72 ) );
  XOR2_X1 \Check1_CheckInst_1_U54  ( .A(Red_AddRoundKeyOutput[28]), .B(
        Red_SignaltoCheck[28]), .Z(\Check1_CheckInst_1_n67 ) );
  XOR2_X1 \Check1_CheckInst_1_U53  ( .A(Red_AddRoundKeyOutput[22]), .B(
        Red_SignaltoCheck[22]), .Z(\Check1_CheckInst_1_n68 ) );
  NOR2_X1 \Check1_CheckInst_1_U52  ( .A1(\Check1_CheckInst_1_n66 ), .A2(
        \Check1_CheckInst_1_n65 ), .ZN(\Check1_CheckInst_1_n90 ) );
  NAND2_X1 \Check1_CheckInst_1_U51  ( .A1(\Check1_CheckInst_1_n64 ), .A2(
        \Check1_CheckInst_1_n63 ), .ZN(\Check1_CheckInst_1_n65 ) );
  NOR2_X1 \Check1_CheckInst_1_U50  ( .A1(Red_SignaltoCheck[100]), .A2(
        Red_SignaltoCheck[118]), .ZN(\Check1_CheckInst_1_n63 ) );
  NOR2_X1 \Check1_CheckInst_1_U49  ( .A1(Red_SignaltoCheck[106]), .A2(
        Red_SignaltoCheck[97]), .ZN(\Check1_CheckInst_1_n64 ) );
  NAND2_X1 \Check1_CheckInst_1_U48  ( .A1(\Check1_CheckInst_1_n62 ), .A2(
        \Check1_CheckInst_1_n61 ), .ZN(\Check1_CheckInst_1_n66 ) );
  NOR2_X1 \Check1_CheckInst_1_U47  ( .A1(Red_SignaltoCheck[133]), .A2(
        Red_SignaltoCheck[124]), .ZN(\Check1_CheckInst_1_n61 ) );
  NOR2_X1 \Check1_CheckInst_1_U46  ( .A1(Red_SignaltoCheck[109]), .A2(
        Red_SignaltoCheck[115]), .ZN(\Check1_CheckInst_1_n62 ) );
  NAND2_X1 \Check1_CheckInst_1_U45  ( .A1(\Check1_CheckInst_1_n60 ), .A2(
        \Check1_CheckInst_1_n59 ), .ZN(\Check1_CheckInst_1_n92 ) );
  NOR2_X1 \Check1_CheckInst_1_U44  ( .A1(\Check1_CheckInst_1_n58 ), .A2(
        \Check1_CheckInst_1_n57 ), .ZN(\Check1_CheckInst_1_n59 ) );
  NAND2_X1 \Check1_CheckInst_1_U43  ( .A1(\Check1_CheckInst_1_n56 ), .A2(
        \Check1_CheckInst_1_n55 ), .ZN(\Check1_CheckInst_1_n57 ) );
  NOR2_X1 \Check1_CheckInst_1_U42  ( .A1(\Check1_CheckInst_1_n54 ), .A2(
        \Check1_CheckInst_1_n53 ), .ZN(\Check1_CheckInst_1_n55 ) );
  XOR2_X1 \Check1_CheckInst_1_U41  ( .A(Red_Feedback[31]), .B(
        Red_SignaltoCheck[79]), .Z(\Check1_CheckInst_1_n53 ) );
  XOR2_X1 \Check1_CheckInst_1_U40  ( .A(Red_Feedback[34]), .B(
        Red_SignaltoCheck[82]), .Z(\Check1_CheckInst_1_n54 ) );
  NOR2_X1 \Check1_CheckInst_1_U39  ( .A1(\Check1_CheckInst_1_n52 ), .A2(
        \Check1_CheckInst_1_n51 ), .ZN(\Check1_CheckInst_1_n56 ) );
  XOR2_X1 \Check1_CheckInst_1_U38  ( .A(Red_Feedback[25]), .B(
        Red_SignaltoCheck[73]), .Z(\Check1_CheckInst_1_n51 ) );
  XOR2_X1 \Check1_CheckInst_1_U37  ( .A(Red_Feedback[37]), .B(
        Red_SignaltoCheck[85]), .Z(\Check1_CheckInst_1_n52 ) );
  NAND2_X1 \Check1_CheckInst_1_U36  ( .A1(\Check1_CheckInst_1_n50 ), .A2(
        \Check1_CheckInst_1_n49 ), .ZN(\Check1_CheckInst_1_n58 ) );
  XNOR2_X1 \Check1_CheckInst_1_U35  ( .A(Red_Feedback[28]), .B(
        Red_SignaltoCheck[76]), .ZN(\Check1_CheckInst_1_n49 ) );
  XNOR2_X1 \Check1_CheckInst_1_U34  ( .A(Red_Feedback[22]), .B(
        Red_SignaltoCheck[70]), .ZN(\Check1_CheckInst_1_n50 ) );
  NOR2_X1 \Check1_CheckInst_1_U33  ( .A1(\Check1_CheckInst_1_n48 ), .A2(
        \Check1_CheckInst_1_n47 ), .ZN(\Check1_CheckInst_1_n60 ) );
  XOR2_X1 \Check1_CheckInst_1_U32  ( .A(Red_Feedback[40]), .B(
        Red_SignaltoCheck[88]), .Z(\Check1_CheckInst_1_n47 ) );
  XOR2_X1 \Check1_CheckInst_1_U31  ( .A(Red_Feedback[43]), .B(
        Red_SignaltoCheck[91]), .Z(\Check1_CheckInst_1_n48 ) );
  NOR2_X1 \Check1_CheckInst_1_U30  ( .A1(\Check1_CheckInst_1_n46 ), .A2(
        \Check1_CheckInst_1_n45 ), .ZN(\Check1_CheckInst_1_n94 ) );
  NAND2_X1 \Check1_CheckInst_1_U29  ( .A1(\Check1_CheckInst_1_n44 ), .A2(
        \Check1_CheckInst_1_n43 ), .ZN(\Check1_CheckInst_1_n45 ) );
  NOR2_X1 \Check1_CheckInst_1_U28  ( .A1(\Check1_CheckInst_1_n42 ), .A2(
        \Check1_CheckInst_1_n41 ), .ZN(\Check1_CheckInst_1_n43 ) );
  NAND2_X1 \Check1_CheckInst_1_U27  ( .A1(\Check1_CheckInst_1_n40 ), .A2(
        \Check1_CheckInst_1_n39 ), .ZN(\Check1_CheckInst_1_n41 ) );
  XNOR2_X1 \Check1_CheckInst_1_U26  ( .A(Red_AddRoundKeyOutput[46]), .B(
        Red_SignaltoCheck[46]), .ZN(\Check1_CheckInst_1_n39 ) );
  XNOR2_X1 \Check1_CheckInst_1_U25  ( .A(Red_Feedback[46]), .B(
        Red_SignaltoCheck[94]), .ZN(\Check1_CheckInst_1_n40 ) );
  NAND2_X1 \Check1_CheckInst_1_U24  ( .A1(\Check1_CheckInst_1_n38 ), .A2(
        \Check1_CheckInst_1_n37 ), .ZN(\Check1_CheckInst_1_n42 ) );
  XNOR2_X1 \Check1_CheckInst_1_U23  ( .A(Red_Feedback[1]), .B(
        Red_SignaltoCheck[49]), .ZN(\Check1_CheckInst_1_n37 ) );
  XNOR2_X1 \Check1_CheckInst_1_U22  ( .A(Red_AddRoundKeyOutput[43]), .B(
        Red_SignaltoCheck[43]), .ZN(\Check1_CheckInst_1_n38 ) );
  NOR2_X1 \Check1_CheckInst_1_U21  ( .A1(\Check1_CheckInst_1_n36 ), .A2(
        \Check1_CheckInst_1_n35 ), .ZN(\Check1_CheckInst_1_n44 ) );
  XOR2_X1 \Check1_CheckInst_1_U20  ( .A(Red_AddRoundKeyOutput[34]), .B(
        Red_SignaltoCheck[34]), .Z(\Check1_CheckInst_1_n35 ) );
  XOR2_X1 \Check1_CheckInst_1_U19  ( .A(Red_AddRoundKeyOutput[37]), .B(
        Red_SignaltoCheck[37]), .Z(\Check1_CheckInst_1_n36 ) );
  NAND2_X1 \Check1_CheckInst_1_U18  ( .A1(\Check1_CheckInst_1_n34 ), .A2(
        \Check1_CheckInst_1_n33 ), .ZN(\Check1_CheckInst_1_n46 ) );
  XNOR2_X1 \Check1_CheckInst_1_U17  ( .A(Red_Feedback[16]), .B(
        Red_SignaltoCheck[64]), .ZN(\Check1_CheckInst_1_n33 ) );
  XNOR2_X1 \Check1_CheckInst_1_U16  ( .A(Red_AddRoundKeyOutput[40]), .B(
        Red_SignaltoCheck[40]), .ZN(\Check1_CheckInst_1_n34 ) );
  NAND2_X1 \Check1_CheckInst_1_U15  ( .A1(\Check1_CheckInst_1_n32 ), .A2(
        \Check1_CheckInst_1_n31 ), .ZN(\Check1_CheckInst_1_n96 ) );
  NOR2_X1 \Check1_CheckInst_1_U14  ( .A1(\Check1_CheckInst_1_n30 ), .A2(
        \Check1_CheckInst_1_n29 ), .ZN(\Check1_CheckInst_1_n31 ) );
  NAND2_X1 \Check1_CheckInst_1_U13  ( .A1(\Check1_CheckInst_1_n28 ), .A2(
        \Check1_CheckInst_1_n27 ), .ZN(\Check1_CheckInst_1_n29 ) );
  NOR2_X1 \Check1_CheckInst_1_U12  ( .A1(\Check1_CheckInst_1_n26 ), .A2(
        \Check1_CheckInst_1_n25 ), .ZN(\Check1_CheckInst_1_n27 ) );
  XOR2_X1 \Check1_CheckInst_1_U11  ( .A(Red_Feedback[19]), .B(
        Red_SignaltoCheck[67]), .Z(\Check1_CheckInst_1_n25 ) );
  XOR2_X1 \Check1_CheckInst_1_U10  ( .A(Red_Feedback[13]), .B(
        Red_SignaltoCheck[61]), .Z(\Check1_CheckInst_1_n26 ) );
  NOR2_X1 \Check1_CheckInst_1_U9  ( .A1(\Check1_CheckInst_1_n24 ), .A2(
        \Check1_CheckInst_1_n23 ), .ZN(\Check1_CheckInst_1_n28 ) );
  XOR2_X1 \Check1_CheckInst_1_U8  ( .A(Red_Feedback[4]), .B(
        Red_SignaltoCheck[52]), .Z(\Check1_CheckInst_1_n23 ) );
  XOR2_X1 \Check1_CheckInst_1_U7  ( .A(Red_Feedback[7]), .B(
        Red_SignaltoCheck[55]), .Z(\Check1_CheckInst_1_n24 ) );
  NAND2_X1 \Check1_CheckInst_1_U6  ( .A1(\Check1_CheckInst_1_n22 ), .A2(
        \Check1_CheckInst_1_n21 ), .ZN(\Check1_CheckInst_1_n30 ) );
  XNOR2_X1 \Check1_CheckInst_1_U5  ( .A(Red_AddRoundKeyOutput[10]), .B(
        Red_SignaltoCheck[10]), .ZN(\Check1_CheckInst_1_n21 ) );
  XNOR2_X1 \Check1_CheckInst_1_U4  ( .A(Red_Feedback[10]), .B(
        Red_SignaltoCheck[58]), .ZN(\Check1_CheckInst_1_n22 ) );
  NOR2_X1 \Check1_CheckInst_1_U3  ( .A1(\Check1_CheckInst_1_n20 ), .A2(
        \Check1_CheckInst_1_n19 ), .ZN(\Check1_CheckInst_1_n32 ) );
  XOR2_X1 \Check1_CheckInst_1_U2  ( .A(Red_AddRoundKeyOutput[13]), .B(
        Red_SignaltoCheck[13]), .Z(\Check1_CheckInst_1_n19 ) );
  XOR2_X1 \Check1_CheckInst_1_U1  ( .A(Red_AddRoundKeyOutput[7]), .B(
        Red_SignaltoCheck[7]), .Z(\Check1_CheckInst_1_n20 ) );
  NOR2_X1 \Check1_CheckInst_2_U79  ( .A1(\Check1_CheckInst_2_n96 ), .A2(
        \Check1_CheckInst_2_n95 ), .ZN(Error[2]) );
  NAND2_X1 \Check1_CheckInst_2_U78  ( .A1(\Check1_CheckInst_2_n94 ), .A2(
        \Check1_CheckInst_2_n93 ), .ZN(\Check1_CheckInst_2_n95 ) );
  NOR2_X1 \Check1_CheckInst_2_U77  ( .A1(\Check1_CheckInst_2_n92 ), .A2(
        \Check1_CheckInst_2_n91 ), .ZN(\Check1_CheckInst_2_n93 ) );
  NAND2_X1 \Check1_CheckInst_2_U76  ( .A1(\Check1_CheckInst_2_n90 ), .A2(
        \Check1_CheckInst_2_n89 ), .ZN(\Check1_CheckInst_2_n91 ) );
  NOR2_X1 \Check1_CheckInst_2_U75  ( .A1(\Check1_CheckInst_2_n88 ), .A2(
        \Check1_CheckInst_2_n87 ), .ZN(\Check1_CheckInst_2_n89 ) );
  NAND2_X1 \Check1_CheckInst_2_U74  ( .A1(\Check1_CheckInst_2_n86 ), .A2(
        \Check1_CheckInst_2_n85 ), .ZN(\Check1_CheckInst_2_n87 ) );
  NOR2_X1 \Check1_CheckInst_2_U73  ( .A1(\Check1_CheckInst_2_n84 ), .A2(
        \Check1_CheckInst_2_n83 ), .ZN(\Check1_CheckInst_2_n85 ) );
  NAND2_X1 \Check1_CheckInst_2_U72  ( .A1(\Check1_CheckInst_2_n82 ), .A2(
        \Check1_CheckInst_2_n81 ), .ZN(\Check1_CheckInst_2_n83 ) );
  XNOR2_X1 \Check1_CheckInst_2_U71  ( .A(Red_AddRoundKeyOutput[26]), .B(
        Red_SignaltoCheck[26]), .ZN(\Check1_CheckInst_2_n81 ) );
  XNOR2_X1 \Check1_CheckInst_2_U70  ( .A(Red_AddRoundKeyOutput[2]), .B(
        Red_SignaltoCheck[2]), .ZN(\Check1_CheckInst_2_n82 ) );
  NAND2_X1 \Check1_CheckInst_2_U69  ( .A1(\Check1_CheckInst_2_n80 ), .A2(
        \Check1_CheckInst_2_n79 ), .ZN(\Check1_CheckInst_2_n84 ) );
  XNOR2_X1 \Check1_CheckInst_2_U68  ( .A(Red_AddRoundKeyOutput[32]), .B(
        Red_SignaltoCheck[32]), .ZN(\Check1_CheckInst_2_n79 ) );
  XNOR2_X1 \Check1_CheckInst_2_U67  ( .A(Red_SignaltoCheck[5]), .B(
        Red_AddRoundKeyOutput[5]), .ZN(\Check1_CheckInst_2_n80 ) );
  NOR2_X1 \Check1_CheckInst_2_U66  ( .A1(\Check1_CheckInst_2_n78 ), .A2(
        \Check1_CheckInst_2_n77 ), .ZN(\Check1_CheckInst_2_n86 ) );
  NAND2_X1 \Check1_CheckInst_2_U65  ( .A1(\Check1_CheckInst_2_n76 ), .A2(
        \Check1_CheckInst_2_n75 ), .ZN(\Check1_CheckInst_2_n77 ) );
  NOR2_X1 \Check1_CheckInst_2_U64  ( .A1(Red_SignaltoCheck[137]), .A2(
        Red_SignaltoCheck[143]), .ZN(\Check1_CheckInst_2_n75 ) );
  NOR2_X1 \Check1_CheckInst_2_U63  ( .A1(Red_SignaltoCheck[128]), .A2(
        Red_SignaltoCheck[122]), .ZN(\Check1_CheckInst_2_n76 ) );
  NAND2_X1 \Check1_CheckInst_2_U62  ( .A1(\Check1_CheckInst_2_n74 ), .A2(
        \Check1_CheckInst_2_n73 ), .ZN(\Check1_CheckInst_2_n78 ) );
  NOR2_X1 \Check1_CheckInst_2_U61  ( .A1(Red_SignaltoCheck[140]), .A2(
        Red_SignaltoCheck[104]), .ZN(\Check1_CheckInst_2_n73 ) );
  NOR2_X1 \Check1_CheckInst_2_U60  ( .A1(Red_SignaltoCheck[131]), .A2(
        Red_SignaltoCheck[113]), .ZN(\Check1_CheckInst_2_n74 ) );
  NAND2_X1 \Check1_CheckInst_2_U59  ( .A1(\Check1_CheckInst_2_n72 ), .A2(
        \Check1_CheckInst_2_n71 ), .ZN(\Check1_CheckInst_2_n88 ) );
  NOR2_X1 \Check1_CheckInst_2_U58  ( .A1(\Check1_CheckInst_2_n70 ), .A2(
        \Check1_CheckInst_2_n69 ), .ZN(\Check1_CheckInst_2_n71 ) );
  XOR2_X1 \Check1_CheckInst_2_U57  ( .A(Red_AddRoundKeyOutput[20]), .B(
        Red_SignaltoCheck[20]), .Z(\Check1_CheckInst_2_n69 ) );
  XOR2_X1 \Check1_CheckInst_2_U56  ( .A(Red_AddRoundKeyOutput[17]), .B(
        Red_SignaltoCheck[17]), .Z(\Check1_CheckInst_2_n70 ) );
  NOR2_X1 \Check1_CheckInst_2_U55  ( .A1(\Check1_CheckInst_2_n68 ), .A2(
        \Check1_CheckInst_2_n67 ), .ZN(\Check1_CheckInst_2_n72 ) );
  XOR2_X1 \Check1_CheckInst_2_U54  ( .A(Red_AddRoundKeyOutput[29]), .B(
        Red_SignaltoCheck[29]), .Z(\Check1_CheckInst_2_n67 ) );
  XOR2_X1 \Check1_CheckInst_2_U53  ( .A(Red_AddRoundKeyOutput[23]), .B(
        Red_SignaltoCheck[23]), .Z(\Check1_CheckInst_2_n68 ) );
  NOR2_X1 \Check1_CheckInst_2_U52  ( .A1(\Check1_CheckInst_2_n66 ), .A2(
        \Check1_CheckInst_2_n65 ), .ZN(\Check1_CheckInst_2_n90 ) );
  NAND2_X1 \Check1_CheckInst_2_U51  ( .A1(\Check1_CheckInst_2_n64 ), .A2(
        \Check1_CheckInst_2_n63 ), .ZN(\Check1_CheckInst_2_n65 ) );
  NOR2_X1 \Check1_CheckInst_2_U50  ( .A1(Red_SignaltoCheck[101]), .A2(
        Red_SignaltoCheck[119]), .ZN(\Check1_CheckInst_2_n63 ) );
  NOR2_X1 \Check1_CheckInst_2_U49  ( .A1(Red_SignaltoCheck[107]), .A2(
        Red_SignaltoCheck[98]), .ZN(\Check1_CheckInst_2_n64 ) );
  NAND2_X1 \Check1_CheckInst_2_U48  ( .A1(\Check1_CheckInst_2_n62 ), .A2(
        \Check1_CheckInst_2_n61 ), .ZN(\Check1_CheckInst_2_n66 ) );
  NOR2_X1 \Check1_CheckInst_2_U47  ( .A1(Red_SignaltoCheck[134]), .A2(
        Red_SignaltoCheck[125]), .ZN(\Check1_CheckInst_2_n61 ) );
  NOR2_X1 \Check1_CheckInst_2_U46  ( .A1(Red_SignaltoCheck[110]), .A2(
        Red_SignaltoCheck[116]), .ZN(\Check1_CheckInst_2_n62 ) );
  NAND2_X1 \Check1_CheckInst_2_U45  ( .A1(\Check1_CheckInst_2_n60 ), .A2(
        \Check1_CheckInst_2_n59 ), .ZN(\Check1_CheckInst_2_n92 ) );
  NOR2_X1 \Check1_CheckInst_2_U44  ( .A1(\Check1_CheckInst_2_n58 ), .A2(
        \Check1_CheckInst_2_n57 ), .ZN(\Check1_CheckInst_2_n59 ) );
  NAND2_X1 \Check1_CheckInst_2_U43  ( .A1(\Check1_CheckInst_2_n56 ), .A2(
        \Check1_CheckInst_2_n55 ), .ZN(\Check1_CheckInst_2_n57 ) );
  NOR2_X1 \Check1_CheckInst_2_U42  ( .A1(\Check1_CheckInst_2_n54 ), .A2(
        \Check1_CheckInst_2_n53 ), .ZN(\Check1_CheckInst_2_n55 ) );
  XOR2_X1 \Check1_CheckInst_2_U41  ( .A(Red_Feedback[32]), .B(
        Red_SignaltoCheck[80]), .Z(\Check1_CheckInst_2_n53 ) );
  XOR2_X1 \Check1_CheckInst_2_U40  ( .A(Red_Feedback[35]), .B(
        Red_SignaltoCheck[83]), .Z(\Check1_CheckInst_2_n54 ) );
  NOR2_X1 \Check1_CheckInst_2_U39  ( .A1(\Check1_CheckInst_2_n52 ), .A2(
        \Check1_CheckInst_2_n51 ), .ZN(\Check1_CheckInst_2_n56 ) );
  XOR2_X1 \Check1_CheckInst_2_U38  ( .A(Red_Feedback[26]), .B(
        Red_SignaltoCheck[74]), .Z(\Check1_CheckInst_2_n51 ) );
  XOR2_X1 \Check1_CheckInst_2_U37  ( .A(Red_Feedback[38]), .B(
        Red_SignaltoCheck[86]), .Z(\Check1_CheckInst_2_n52 ) );
  NAND2_X1 \Check1_CheckInst_2_U36  ( .A1(\Check1_CheckInst_2_n50 ), .A2(
        \Check1_CheckInst_2_n49 ), .ZN(\Check1_CheckInst_2_n58 ) );
  XNOR2_X1 \Check1_CheckInst_2_U35  ( .A(Red_Feedback[29]), .B(
        Red_SignaltoCheck[77]), .ZN(\Check1_CheckInst_2_n49 ) );
  XNOR2_X1 \Check1_CheckInst_2_U34  ( .A(Red_Feedback[23]), .B(
        Red_SignaltoCheck[71]), .ZN(\Check1_CheckInst_2_n50 ) );
  NOR2_X1 \Check1_CheckInst_2_U33  ( .A1(\Check1_CheckInst_2_n48 ), .A2(
        \Check1_CheckInst_2_n47 ), .ZN(\Check1_CheckInst_2_n60 ) );
  XOR2_X1 \Check1_CheckInst_2_U32  ( .A(Red_Feedback[41]), .B(
        Red_SignaltoCheck[89]), .Z(\Check1_CheckInst_2_n47 ) );
  XOR2_X1 \Check1_CheckInst_2_U31  ( .A(Red_Feedback[44]), .B(
        Red_SignaltoCheck[92]), .Z(\Check1_CheckInst_2_n48 ) );
  NOR2_X1 \Check1_CheckInst_2_U30  ( .A1(\Check1_CheckInst_2_n46 ), .A2(
        \Check1_CheckInst_2_n45 ), .ZN(\Check1_CheckInst_2_n94 ) );
  NAND2_X1 \Check1_CheckInst_2_U29  ( .A1(\Check1_CheckInst_2_n44 ), .A2(
        \Check1_CheckInst_2_n43 ), .ZN(\Check1_CheckInst_2_n45 ) );
  NOR2_X1 \Check1_CheckInst_2_U28  ( .A1(\Check1_CheckInst_2_n42 ), .A2(
        \Check1_CheckInst_2_n41 ), .ZN(\Check1_CheckInst_2_n43 ) );
  NAND2_X1 \Check1_CheckInst_2_U27  ( .A1(\Check1_CheckInst_2_n40 ), .A2(
        \Check1_CheckInst_2_n39 ), .ZN(\Check1_CheckInst_2_n41 ) );
  XNOR2_X1 \Check1_CheckInst_2_U26  ( .A(Red_AddRoundKeyOutput[47]), .B(
        Red_SignaltoCheck[47]), .ZN(\Check1_CheckInst_2_n39 ) );
  XNOR2_X1 \Check1_CheckInst_2_U25  ( .A(Red_Feedback[47]), .B(
        Red_SignaltoCheck[95]), .ZN(\Check1_CheckInst_2_n40 ) );
  NAND2_X1 \Check1_CheckInst_2_U24  ( .A1(\Check1_CheckInst_2_n38 ), .A2(
        \Check1_CheckInst_2_n37 ), .ZN(\Check1_CheckInst_2_n42 ) );
  XNOR2_X1 \Check1_CheckInst_2_U23  ( .A(Red_Feedback[2]), .B(
        Red_SignaltoCheck[50]), .ZN(\Check1_CheckInst_2_n37 ) );
  XNOR2_X1 \Check1_CheckInst_2_U22  ( .A(Red_AddRoundKeyOutput[44]), .B(
        Red_SignaltoCheck[44]), .ZN(\Check1_CheckInst_2_n38 ) );
  NOR2_X1 \Check1_CheckInst_2_U21  ( .A1(\Check1_CheckInst_2_n36 ), .A2(
        \Check1_CheckInst_2_n35 ), .ZN(\Check1_CheckInst_2_n44 ) );
  XOR2_X1 \Check1_CheckInst_2_U20  ( .A(Red_AddRoundKeyOutput[35]), .B(
        Red_SignaltoCheck[35]), .Z(\Check1_CheckInst_2_n35 ) );
  XOR2_X1 \Check1_CheckInst_2_U19  ( .A(Red_AddRoundKeyOutput[38]), .B(
        Red_SignaltoCheck[38]), .Z(\Check1_CheckInst_2_n36 ) );
  NAND2_X1 \Check1_CheckInst_2_U18  ( .A1(\Check1_CheckInst_2_n34 ), .A2(
        \Check1_CheckInst_2_n33 ), .ZN(\Check1_CheckInst_2_n46 ) );
  XNOR2_X1 \Check1_CheckInst_2_U17  ( .A(Red_Feedback[17]), .B(
        Red_SignaltoCheck[65]), .ZN(\Check1_CheckInst_2_n33 ) );
  XNOR2_X1 \Check1_CheckInst_2_U16  ( .A(Red_AddRoundKeyOutput[41]), .B(
        Red_SignaltoCheck[41]), .ZN(\Check1_CheckInst_2_n34 ) );
  NAND2_X1 \Check1_CheckInst_2_U15  ( .A1(\Check1_CheckInst_2_n32 ), .A2(
        \Check1_CheckInst_2_n31 ), .ZN(\Check1_CheckInst_2_n96 ) );
  NOR2_X1 \Check1_CheckInst_2_U14  ( .A1(\Check1_CheckInst_2_n30 ), .A2(
        \Check1_CheckInst_2_n29 ), .ZN(\Check1_CheckInst_2_n31 ) );
  NAND2_X1 \Check1_CheckInst_2_U13  ( .A1(\Check1_CheckInst_2_n28 ), .A2(
        \Check1_CheckInst_2_n27 ), .ZN(\Check1_CheckInst_2_n29 ) );
  NOR2_X1 \Check1_CheckInst_2_U12  ( .A1(\Check1_CheckInst_2_n26 ), .A2(
        \Check1_CheckInst_2_n25 ), .ZN(\Check1_CheckInst_2_n27 ) );
  XOR2_X1 \Check1_CheckInst_2_U11  ( .A(Red_Feedback[20]), .B(
        Red_SignaltoCheck[68]), .Z(\Check1_CheckInst_2_n25 ) );
  XOR2_X1 \Check1_CheckInst_2_U10  ( .A(Red_Feedback[14]), .B(
        Red_SignaltoCheck[62]), .Z(\Check1_CheckInst_2_n26 ) );
  NOR2_X1 \Check1_CheckInst_2_U9  ( .A1(\Check1_CheckInst_2_n24 ), .A2(
        \Check1_CheckInst_2_n23 ), .ZN(\Check1_CheckInst_2_n28 ) );
  XOR2_X1 \Check1_CheckInst_2_U8  ( .A(Red_Feedback[5]), .B(
        Red_SignaltoCheck[53]), .Z(\Check1_CheckInst_2_n23 ) );
  XOR2_X1 \Check1_CheckInst_2_U7  ( .A(Red_Feedback[8]), .B(
        Red_SignaltoCheck[56]), .Z(\Check1_CheckInst_2_n24 ) );
  NAND2_X1 \Check1_CheckInst_2_U6  ( .A1(\Check1_CheckInst_2_n22 ), .A2(
        \Check1_CheckInst_2_n21 ), .ZN(\Check1_CheckInst_2_n30 ) );
  XNOR2_X1 \Check1_CheckInst_2_U5  ( .A(Red_AddRoundKeyOutput[11]), .B(
        Red_SignaltoCheck[11]), .ZN(\Check1_CheckInst_2_n21 ) );
  XNOR2_X1 \Check1_CheckInst_2_U4  ( .A(Red_Feedback[11]), .B(
        Red_SignaltoCheck[59]), .ZN(\Check1_CheckInst_2_n22 ) );
  NOR2_X1 \Check1_CheckInst_2_U3  ( .A1(\Check1_CheckInst_2_n20 ), .A2(
        \Check1_CheckInst_2_n19 ), .ZN(\Check1_CheckInst_2_n32 ) );
  XOR2_X1 \Check1_CheckInst_2_U2  ( .A(Red_AddRoundKeyOutput[14]), .B(
        Red_SignaltoCheck[14]), .Z(\Check1_CheckInst_2_n19 ) );
  XOR2_X1 \Check1_CheckInst_2_U1  ( .A(Red_AddRoundKeyOutput[8]), .B(
        Red_SignaltoCheck[8]), .Z(\Check1_CheckInst_2_n20 ) );
endmodule

