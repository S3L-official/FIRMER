module LED64Enc ( clk, rst, Plaintext, Key, Ciphertext );
  input [63:0] Plaintext;
  input [63:0] Key;
  output [63:0] Ciphertext;
  (* FIRMER="clock" *)input clk;
  (* FIRMER="control" *)input rst;
  wire   SubCellInst_LFInst_0_LFInst_3_n16 ,
         SubCellInst_LFInst_0_LFInst_3_n15 ,
         SubCellInst_LFInst_0_LFInst_3_n14 ,
         SubCellInst_LFInst_0_LFInst_3_n13 ,
         SubCellInst_LFInst_0_LFInst_3_n12 ,
         SubCellInst_LFInst_0_LFInst_3_n11 ,
         SubCellInst_LFInst_0_LFInst_2_n22 ,
         SubCellInst_LFInst_0_LFInst_2_n21 ,
         SubCellInst_LFInst_0_LFInst_2_n20 ,
         SubCellInst_LFInst_0_LFInst_2_n19 ,
         SubCellInst_LFInst_0_LFInst_2_n18 ,
         SubCellInst_LFInst_0_LFInst_2_n17 ,
         SubCellInst_LFInst_0_LFInst_2_n16 ,
         SubCellInst_LFInst_0_LFInst_2_n15 ,
         SubCellInst_LFInst_0_LFInst_1_n18 ,
         SubCellInst_LFInst_0_LFInst_1_n17 ,
         SubCellInst_LFInst_0_LFInst_1_n16 ,
         SubCellInst_LFInst_0_LFInst_1_n15 ,
         SubCellInst_LFInst_0_LFInst_1_n14 ,
         SubCellInst_LFInst_0_LFInst_1_n13 ,
         SubCellInst_LFInst_0_LFInst_1_n12 ,
         SubCellInst_LFInst_0_LFInst_1_n11 ,
         SubCellInst_LFInst_0_LFInst_1_n10 ,
         SubCellInst_LFInst_0_LFInst_0_n6 ,
         SubCellInst_LFInst_0_LFInst_0_n5 ,
         SubCellInst_LFInst_0_LFInst_0_n4 ,
         SubCellInst_LFInst_1_LFInst_3_n16 ,
         SubCellInst_LFInst_1_LFInst_3_n15 ,
         SubCellInst_LFInst_1_LFInst_3_n14 ,
         SubCellInst_LFInst_1_LFInst_3_n13 ,
         SubCellInst_LFInst_1_LFInst_3_n12 ,
         SubCellInst_LFInst_1_LFInst_3_n11 ,
         SubCellInst_LFInst_1_LFInst_2_n22 ,
         SubCellInst_LFInst_1_LFInst_2_n21 ,
         SubCellInst_LFInst_1_LFInst_2_n20 ,
         SubCellInst_LFInst_1_LFInst_2_n19 ,
         SubCellInst_LFInst_1_LFInst_2_n18 ,
         SubCellInst_LFInst_1_LFInst_2_n17 ,
         SubCellInst_LFInst_1_LFInst_2_n16 ,
         SubCellInst_LFInst_1_LFInst_2_n15 ,
         SubCellInst_LFInst_1_LFInst_1_n18 ,
         SubCellInst_LFInst_1_LFInst_1_n17 ,
         SubCellInst_LFInst_1_LFInst_1_n16 ,
         SubCellInst_LFInst_1_LFInst_1_n15 ,
         SubCellInst_LFInst_1_LFInst_1_n14 ,
         SubCellInst_LFInst_1_LFInst_1_n13 ,
         SubCellInst_LFInst_1_LFInst_1_n12 ,
         SubCellInst_LFInst_1_LFInst_1_n11 ,
         SubCellInst_LFInst_1_LFInst_1_n10 ,
         SubCellInst_LFInst_1_LFInst_0_n6 ,
         SubCellInst_LFInst_1_LFInst_0_n5 ,
         SubCellInst_LFInst_1_LFInst_0_n4 ,
         SubCellInst_LFInst_2_LFInst_3_n16 ,
         SubCellInst_LFInst_2_LFInst_3_n15 ,
         SubCellInst_LFInst_2_LFInst_3_n14 ,
         SubCellInst_LFInst_2_LFInst_3_n13 ,
         SubCellInst_LFInst_2_LFInst_3_n12 ,
         SubCellInst_LFInst_2_LFInst_3_n11 ,
         SubCellInst_LFInst_2_LFInst_2_n22 ,
         SubCellInst_LFInst_2_LFInst_2_n21 ,
         SubCellInst_LFInst_2_LFInst_2_n20 ,
         SubCellInst_LFInst_2_LFInst_2_n19 ,
         SubCellInst_LFInst_2_LFInst_2_n18 ,
         SubCellInst_LFInst_2_LFInst_2_n17 ,
         SubCellInst_LFInst_2_LFInst_2_n16 ,
         SubCellInst_LFInst_2_LFInst_2_n15 ,
         SubCellInst_LFInst_2_LFInst_1_n18 ,
         SubCellInst_LFInst_2_LFInst_1_n17 ,
         SubCellInst_LFInst_2_LFInst_1_n16 ,
         SubCellInst_LFInst_2_LFInst_1_n15 ,
         SubCellInst_LFInst_2_LFInst_1_n14 ,
         SubCellInst_LFInst_2_LFInst_1_n13 ,
         SubCellInst_LFInst_2_LFInst_1_n12 ,
         SubCellInst_LFInst_2_LFInst_1_n11 ,
         SubCellInst_LFInst_2_LFInst_1_n10 ,
         SubCellInst_LFInst_2_LFInst_0_n6 ,
         SubCellInst_LFInst_2_LFInst_0_n5 ,
         SubCellInst_LFInst_2_LFInst_0_n4 ,
         SubCellInst_LFInst_3_LFInst_3_n16 ,
         SubCellInst_LFInst_3_LFInst_3_n15 ,
         SubCellInst_LFInst_3_LFInst_3_n14 ,
         SubCellInst_LFInst_3_LFInst_3_n13 ,
         SubCellInst_LFInst_3_LFInst_3_n12 ,
         SubCellInst_LFInst_3_LFInst_3_n11 ,
         SubCellInst_LFInst_3_LFInst_2_n22 ,
         SubCellInst_LFInst_3_LFInst_2_n21 ,
         SubCellInst_LFInst_3_LFInst_2_n20 ,
         SubCellInst_LFInst_3_LFInst_2_n19 ,
         SubCellInst_LFInst_3_LFInst_2_n18 ,
         SubCellInst_LFInst_3_LFInst_2_n17 ,
         SubCellInst_LFInst_3_LFInst_2_n16 ,
         SubCellInst_LFInst_3_LFInst_2_n15 ,
         SubCellInst_LFInst_3_LFInst_1_n18 ,
         SubCellInst_LFInst_3_LFInst_1_n17 ,
         SubCellInst_LFInst_3_LFInst_1_n16 ,
         SubCellInst_LFInst_3_LFInst_1_n15 ,
         SubCellInst_LFInst_3_LFInst_1_n14 ,
         SubCellInst_LFInst_3_LFInst_1_n13 ,
         SubCellInst_LFInst_3_LFInst_1_n12 ,
         SubCellInst_LFInst_3_LFInst_1_n11 ,
         SubCellInst_LFInst_3_LFInst_1_n10 ,
         SubCellInst_LFInst_3_LFInst_0_n6 ,
         SubCellInst_LFInst_3_LFInst_0_n5 ,
         SubCellInst_LFInst_3_LFInst_0_n4 ,
         SubCellInst_LFInst_4_LFInst_3_n16 ,
         SubCellInst_LFInst_4_LFInst_3_n15 ,
         SubCellInst_LFInst_4_LFInst_3_n14 ,
         SubCellInst_LFInst_4_LFInst_3_n13 ,
         SubCellInst_LFInst_4_LFInst_3_n12 ,
         SubCellInst_LFInst_4_LFInst_3_n11 ,
         SubCellInst_LFInst_4_LFInst_2_n22 ,
         SubCellInst_LFInst_4_LFInst_2_n21 ,
         SubCellInst_LFInst_4_LFInst_2_n20 ,
         SubCellInst_LFInst_4_LFInst_2_n19 ,
         SubCellInst_LFInst_4_LFInst_2_n18 ,
         SubCellInst_LFInst_4_LFInst_2_n17 ,
         SubCellInst_LFInst_4_LFInst_2_n16 ,
         SubCellInst_LFInst_4_LFInst_2_n15 ,
         SubCellInst_LFInst_4_LFInst_1_n18 ,
         SubCellInst_LFInst_4_LFInst_1_n17 ,
         SubCellInst_LFInst_4_LFInst_1_n16 ,
         SubCellInst_LFInst_4_LFInst_1_n15 ,
         SubCellInst_LFInst_4_LFInst_1_n14 ,
         SubCellInst_LFInst_4_LFInst_1_n13 ,
         SubCellInst_LFInst_4_LFInst_1_n12 ,
         SubCellInst_LFInst_4_LFInst_1_n11 ,
         SubCellInst_LFInst_4_LFInst_1_n10 ,
         SubCellInst_LFInst_4_LFInst_0_n6 ,
         SubCellInst_LFInst_4_LFInst_0_n5 ,
         SubCellInst_LFInst_4_LFInst_0_n4 ,
         SubCellInst_LFInst_5_LFInst_3_n16 ,
         SubCellInst_LFInst_5_LFInst_3_n15 ,
         SubCellInst_LFInst_5_LFInst_3_n14 ,
         SubCellInst_LFInst_5_LFInst_3_n13 ,
         SubCellInst_LFInst_5_LFInst_3_n12 ,
         SubCellInst_LFInst_5_LFInst_3_n11 ,
         SubCellInst_LFInst_5_LFInst_2_n22 ,
         SubCellInst_LFInst_5_LFInst_2_n21 ,
         SubCellInst_LFInst_5_LFInst_2_n20 ,
         SubCellInst_LFInst_5_LFInst_2_n19 ,
         SubCellInst_LFInst_5_LFInst_2_n18 ,
         SubCellInst_LFInst_5_LFInst_2_n17 ,
         SubCellInst_LFInst_5_LFInst_2_n16 ,
         SubCellInst_LFInst_5_LFInst_2_n15 ,
         SubCellInst_LFInst_5_LFInst_1_n18 ,
         SubCellInst_LFInst_5_LFInst_1_n17 ,
         SubCellInst_LFInst_5_LFInst_1_n16 ,
         SubCellInst_LFInst_5_LFInst_1_n15 ,
         SubCellInst_LFInst_5_LFInst_1_n14 ,
         SubCellInst_LFInst_5_LFInst_1_n13 ,
         SubCellInst_LFInst_5_LFInst_1_n12 ,
         SubCellInst_LFInst_5_LFInst_1_n11 ,
         SubCellInst_LFInst_5_LFInst_1_n10 ,
         SubCellInst_LFInst_5_LFInst_0_n6 ,
         SubCellInst_LFInst_5_LFInst_0_n5 ,
         SubCellInst_LFInst_5_LFInst_0_n4 ,
         SubCellInst_LFInst_6_LFInst_3_n16 ,
         SubCellInst_LFInst_6_LFInst_3_n15 ,
         SubCellInst_LFInst_6_LFInst_3_n14 ,
         SubCellInst_LFInst_6_LFInst_3_n13 ,
         SubCellInst_LFInst_6_LFInst_3_n12 ,
         SubCellInst_LFInst_6_LFInst_3_n11 ,
         SubCellInst_LFInst_6_LFInst_2_n22 ,
         SubCellInst_LFInst_6_LFInst_2_n21 ,
         SubCellInst_LFInst_6_LFInst_2_n20 ,
         SubCellInst_LFInst_6_LFInst_2_n19 ,
         SubCellInst_LFInst_6_LFInst_2_n18 ,
         SubCellInst_LFInst_6_LFInst_2_n17 ,
         SubCellInst_LFInst_6_LFInst_2_n16 ,
         SubCellInst_LFInst_6_LFInst_2_n15 ,
         SubCellInst_LFInst_6_LFInst_1_n18 ,
         SubCellInst_LFInst_6_LFInst_1_n17 ,
         SubCellInst_LFInst_6_LFInst_1_n16 ,
         SubCellInst_LFInst_6_LFInst_1_n15 ,
         SubCellInst_LFInst_6_LFInst_1_n14 ,
         SubCellInst_LFInst_6_LFInst_1_n13 ,
         SubCellInst_LFInst_6_LFInst_1_n12 ,
         SubCellInst_LFInst_6_LFInst_1_n11 ,
         SubCellInst_LFInst_6_LFInst_1_n10 ,
         SubCellInst_LFInst_6_LFInst_0_n6 ,
         SubCellInst_LFInst_6_LFInst_0_n5 ,
         SubCellInst_LFInst_6_LFInst_0_n4 ,
         SubCellInst_LFInst_7_LFInst_3_n16 ,
         SubCellInst_LFInst_7_LFInst_3_n15 ,
         SubCellInst_LFInst_7_LFInst_3_n14 ,
         SubCellInst_LFInst_7_LFInst_3_n13 ,
         SubCellInst_LFInst_7_LFInst_3_n12 ,
         SubCellInst_LFInst_7_LFInst_3_n11 ,
         SubCellInst_LFInst_7_LFInst_2_n22 ,
         SubCellInst_LFInst_7_LFInst_2_n21 ,
         SubCellInst_LFInst_7_LFInst_2_n20 ,
         SubCellInst_LFInst_7_LFInst_2_n19 ,
         SubCellInst_LFInst_7_LFInst_2_n18 ,
         SubCellInst_LFInst_7_LFInst_2_n17 ,
         SubCellInst_LFInst_7_LFInst_2_n16 ,
         SubCellInst_LFInst_7_LFInst_2_n15 ,
         SubCellInst_LFInst_7_LFInst_1_n18 ,
         SubCellInst_LFInst_7_LFInst_1_n17 ,
         SubCellInst_LFInst_7_LFInst_1_n16 ,
         SubCellInst_LFInst_7_LFInst_1_n15 ,
         SubCellInst_LFInst_7_LFInst_1_n14 ,
         SubCellInst_LFInst_7_LFInst_1_n13 ,
         SubCellInst_LFInst_7_LFInst_1_n12 ,
         SubCellInst_LFInst_7_LFInst_1_n11 ,
         SubCellInst_LFInst_7_LFInst_1_n10 ,
         SubCellInst_LFInst_7_LFInst_0_n6 ,
         SubCellInst_LFInst_7_LFInst_0_n5 ,
         SubCellInst_LFInst_7_LFInst_0_n4 ,
         SubCellInst_LFInst_8_LFInst_3_n16 ,
         SubCellInst_LFInst_8_LFInst_3_n15 ,
         SubCellInst_LFInst_8_LFInst_3_n14 ,
         SubCellInst_LFInst_8_LFInst_3_n13 ,
         SubCellInst_LFInst_8_LFInst_3_n12 ,
         SubCellInst_LFInst_8_LFInst_3_n11 ,
         SubCellInst_LFInst_8_LFInst_2_n22 ,
         SubCellInst_LFInst_8_LFInst_2_n21 ,
         SubCellInst_LFInst_8_LFInst_2_n20 ,
         SubCellInst_LFInst_8_LFInst_2_n19 ,
         SubCellInst_LFInst_8_LFInst_2_n18 ,
         SubCellInst_LFInst_8_LFInst_2_n17 ,
         SubCellInst_LFInst_8_LFInst_2_n16 ,
         SubCellInst_LFInst_8_LFInst_2_n15 ,
         SubCellInst_LFInst_8_LFInst_1_n18 ,
         SubCellInst_LFInst_8_LFInst_1_n17 ,
         SubCellInst_LFInst_8_LFInst_1_n16 ,
         SubCellInst_LFInst_8_LFInst_1_n15 ,
         SubCellInst_LFInst_8_LFInst_1_n14 ,
         SubCellInst_LFInst_8_LFInst_1_n13 ,
         SubCellInst_LFInst_8_LFInst_1_n12 ,
         SubCellInst_LFInst_8_LFInst_1_n11 ,
         SubCellInst_LFInst_8_LFInst_1_n10 ,
         SubCellInst_LFInst_8_LFInst_0_n6 ,
         SubCellInst_LFInst_8_LFInst_0_n5 ,
         SubCellInst_LFInst_8_LFInst_0_n4 ,
         SubCellInst_LFInst_9_LFInst_3_n16 ,
         SubCellInst_LFInst_9_LFInst_3_n15 ,
         SubCellInst_LFInst_9_LFInst_3_n14 ,
         SubCellInst_LFInst_9_LFInst_3_n13 ,
         SubCellInst_LFInst_9_LFInst_3_n12 ,
         SubCellInst_LFInst_9_LFInst_3_n11 ,
         SubCellInst_LFInst_9_LFInst_2_n22 ,
         SubCellInst_LFInst_9_LFInst_2_n21 ,
         SubCellInst_LFInst_9_LFInst_2_n20 ,
         SubCellInst_LFInst_9_LFInst_2_n19 ,
         SubCellInst_LFInst_9_LFInst_2_n18 ,
         SubCellInst_LFInst_9_LFInst_2_n17 ,
         SubCellInst_LFInst_9_LFInst_2_n16 ,
         SubCellInst_LFInst_9_LFInst_2_n15 ,
         SubCellInst_LFInst_9_LFInst_1_n18 ,
         SubCellInst_LFInst_9_LFInst_1_n17 ,
         SubCellInst_LFInst_9_LFInst_1_n16 ,
         SubCellInst_LFInst_9_LFInst_1_n15 ,
         SubCellInst_LFInst_9_LFInst_1_n14 ,
         SubCellInst_LFInst_9_LFInst_1_n13 ,
         SubCellInst_LFInst_9_LFInst_1_n12 ,
         SubCellInst_LFInst_9_LFInst_1_n11 ,
         SubCellInst_LFInst_9_LFInst_1_n10 ,
         SubCellInst_LFInst_9_LFInst_0_n6 ,
         SubCellInst_LFInst_9_LFInst_0_n5 ,
         SubCellInst_LFInst_9_LFInst_0_n4 ,
         SubCellInst_LFInst_10_LFInst_3_n16 ,
         SubCellInst_LFInst_10_LFInst_3_n15 ,
         SubCellInst_LFInst_10_LFInst_3_n14 ,
         SubCellInst_LFInst_10_LFInst_3_n13 ,
         SubCellInst_LFInst_10_LFInst_3_n12 ,
         SubCellInst_LFInst_10_LFInst_3_n11 ,
         SubCellInst_LFInst_10_LFInst_2_n22 ,
         SubCellInst_LFInst_10_LFInst_2_n21 ,
         SubCellInst_LFInst_10_LFInst_2_n20 ,
         SubCellInst_LFInst_10_LFInst_2_n19 ,
         SubCellInst_LFInst_10_LFInst_2_n18 ,
         SubCellInst_LFInst_10_LFInst_2_n17 ,
         SubCellInst_LFInst_10_LFInst_2_n16 ,
         SubCellInst_LFInst_10_LFInst_2_n15 ,
         SubCellInst_LFInst_10_LFInst_1_n18 ,
         SubCellInst_LFInst_10_LFInst_1_n17 ,
         SubCellInst_LFInst_10_LFInst_1_n16 ,
         SubCellInst_LFInst_10_LFInst_1_n15 ,
         SubCellInst_LFInst_10_LFInst_1_n14 ,
         SubCellInst_LFInst_10_LFInst_1_n13 ,
         SubCellInst_LFInst_10_LFInst_1_n12 ,
         SubCellInst_LFInst_10_LFInst_1_n11 ,
         SubCellInst_LFInst_10_LFInst_1_n10 ,
         SubCellInst_LFInst_10_LFInst_0_n6 ,
         SubCellInst_LFInst_10_LFInst_0_n5 ,
         SubCellInst_LFInst_10_LFInst_0_n4 ,
         SubCellInst_LFInst_11_LFInst_3_n16 ,
         SubCellInst_LFInst_11_LFInst_3_n15 ,
         SubCellInst_LFInst_11_LFInst_3_n14 ,
         SubCellInst_LFInst_11_LFInst_3_n13 ,
         SubCellInst_LFInst_11_LFInst_3_n12 ,
         SubCellInst_LFInst_11_LFInst_3_n11 ,
         SubCellInst_LFInst_11_LFInst_2_n22 ,
         SubCellInst_LFInst_11_LFInst_2_n21 ,
         SubCellInst_LFInst_11_LFInst_2_n20 ,
         SubCellInst_LFInst_11_LFInst_2_n19 ,
         SubCellInst_LFInst_11_LFInst_2_n18 ,
         SubCellInst_LFInst_11_LFInst_2_n17 ,
         SubCellInst_LFInst_11_LFInst_2_n16 ,
         SubCellInst_LFInst_11_LFInst_2_n15 ,
         SubCellInst_LFInst_11_LFInst_1_n18 ,
         SubCellInst_LFInst_11_LFInst_1_n17 ,
         SubCellInst_LFInst_11_LFInst_1_n16 ,
         SubCellInst_LFInst_11_LFInst_1_n15 ,
         SubCellInst_LFInst_11_LFInst_1_n14 ,
         SubCellInst_LFInst_11_LFInst_1_n13 ,
         SubCellInst_LFInst_11_LFInst_1_n12 ,
         SubCellInst_LFInst_11_LFInst_1_n11 ,
         SubCellInst_LFInst_11_LFInst_1_n10 ,
         SubCellInst_LFInst_11_LFInst_0_n6 ,
         SubCellInst_LFInst_11_LFInst_0_n5 ,
         SubCellInst_LFInst_11_LFInst_0_n4 ,
         SubCellInst_LFInst_12_LFInst_3_n16 ,
         SubCellInst_LFInst_12_LFInst_3_n15 ,
         SubCellInst_LFInst_12_LFInst_3_n14 ,
         SubCellInst_LFInst_12_LFInst_3_n13 ,
         SubCellInst_LFInst_12_LFInst_3_n12 ,
         SubCellInst_LFInst_12_LFInst_3_n11 ,
         SubCellInst_LFInst_12_LFInst_2_n22 ,
         SubCellInst_LFInst_12_LFInst_2_n21 ,
         SubCellInst_LFInst_12_LFInst_2_n20 ,
         SubCellInst_LFInst_12_LFInst_2_n19 ,
         SubCellInst_LFInst_12_LFInst_2_n18 ,
         SubCellInst_LFInst_12_LFInst_2_n17 ,
         SubCellInst_LFInst_12_LFInst_2_n16 ,
         SubCellInst_LFInst_12_LFInst_2_n15 ,
         SubCellInst_LFInst_12_LFInst_1_n18 ,
         SubCellInst_LFInst_12_LFInst_1_n17 ,
         SubCellInst_LFInst_12_LFInst_1_n16 ,
         SubCellInst_LFInst_12_LFInst_1_n15 ,
         SubCellInst_LFInst_12_LFInst_1_n14 ,
         SubCellInst_LFInst_12_LFInst_1_n13 ,
         SubCellInst_LFInst_12_LFInst_1_n12 ,
         SubCellInst_LFInst_12_LFInst_1_n11 ,
         SubCellInst_LFInst_12_LFInst_1_n10 ,
         SubCellInst_LFInst_12_LFInst_0_n6 ,
         SubCellInst_LFInst_12_LFInst_0_n5 ,
         SubCellInst_LFInst_12_LFInst_0_n4 ,
         SubCellInst_LFInst_13_LFInst_3_n16 ,
         SubCellInst_LFInst_13_LFInst_3_n15 ,
         SubCellInst_LFInst_13_LFInst_3_n14 ,
         SubCellInst_LFInst_13_LFInst_3_n13 ,
         SubCellInst_LFInst_13_LFInst_3_n12 ,
         SubCellInst_LFInst_13_LFInst_3_n11 ,
         SubCellInst_LFInst_13_LFInst_2_n22 ,
         SubCellInst_LFInst_13_LFInst_2_n21 ,
         SubCellInst_LFInst_13_LFInst_2_n20 ,
         SubCellInst_LFInst_13_LFInst_2_n19 ,
         SubCellInst_LFInst_13_LFInst_2_n18 ,
         SubCellInst_LFInst_13_LFInst_2_n17 ,
         SubCellInst_LFInst_13_LFInst_2_n16 ,
         SubCellInst_LFInst_13_LFInst_2_n15 ,
         SubCellInst_LFInst_13_LFInst_1_n18 ,
         SubCellInst_LFInst_13_LFInst_1_n17 ,
         SubCellInst_LFInst_13_LFInst_1_n16 ,
         SubCellInst_LFInst_13_LFInst_1_n15 ,
         SubCellInst_LFInst_13_LFInst_1_n14 ,
         SubCellInst_LFInst_13_LFInst_1_n13 ,
         SubCellInst_LFInst_13_LFInst_1_n12 ,
         SubCellInst_LFInst_13_LFInst_1_n11 ,
         SubCellInst_LFInst_13_LFInst_1_n10 ,
         SubCellInst_LFInst_13_LFInst_0_n6 ,
         SubCellInst_LFInst_13_LFInst_0_n5 ,
         SubCellInst_LFInst_13_LFInst_0_n4 ,
         SubCellInst_LFInst_14_LFInst_3_n16 ,
         SubCellInst_LFInst_14_LFInst_3_n15 ,
         SubCellInst_LFInst_14_LFInst_3_n14 ,
         SubCellInst_LFInst_14_LFInst_3_n13 ,
         SubCellInst_LFInst_14_LFInst_3_n12 ,
         SubCellInst_LFInst_14_LFInst_3_n11 ,
         SubCellInst_LFInst_14_LFInst_2_n22 ,
         SubCellInst_LFInst_14_LFInst_2_n21 ,
         SubCellInst_LFInst_14_LFInst_2_n20 ,
         SubCellInst_LFInst_14_LFInst_2_n19 ,
         SubCellInst_LFInst_14_LFInst_2_n18 ,
         SubCellInst_LFInst_14_LFInst_2_n17 ,
         SubCellInst_LFInst_14_LFInst_2_n16 ,
         SubCellInst_LFInst_14_LFInst_2_n15 ,
         SubCellInst_LFInst_14_LFInst_1_n18 ,
         SubCellInst_LFInst_14_LFInst_1_n17 ,
         SubCellInst_LFInst_14_LFInst_1_n16 ,
         SubCellInst_LFInst_14_LFInst_1_n15 ,
         SubCellInst_LFInst_14_LFInst_1_n14 ,
         SubCellInst_LFInst_14_LFInst_1_n13 ,
         SubCellInst_LFInst_14_LFInst_1_n12 ,
         SubCellInst_LFInst_14_LFInst_1_n11 ,
         SubCellInst_LFInst_14_LFInst_1_n10 ,
         SubCellInst_LFInst_14_LFInst_0_n6 ,
         SubCellInst_LFInst_14_LFInst_0_n5 ,
         SubCellInst_LFInst_14_LFInst_0_n4 ,
         SubCellInst_LFInst_15_LFInst_3_n16 ,
         SubCellInst_LFInst_15_LFInst_3_n15 ,
         SubCellInst_LFInst_15_LFInst_3_n14 ,
         SubCellInst_LFInst_15_LFInst_3_n13 ,
         SubCellInst_LFInst_15_LFInst_3_n12 ,
         SubCellInst_LFInst_15_LFInst_3_n11 ,
         SubCellInst_LFInst_15_LFInst_2_n22 ,
         SubCellInst_LFInst_15_LFInst_2_n21 ,
         SubCellInst_LFInst_15_LFInst_2_n20 ,
         SubCellInst_LFInst_15_LFInst_2_n19 ,
         SubCellInst_LFInst_15_LFInst_2_n18 ,
         SubCellInst_LFInst_15_LFInst_2_n17 ,
         SubCellInst_LFInst_15_LFInst_2_n16 ,
         SubCellInst_LFInst_15_LFInst_2_n15 ,
         SubCellInst_LFInst_15_LFInst_1_n18 ,
         SubCellInst_LFInst_15_LFInst_1_n17 ,
         SubCellInst_LFInst_15_LFInst_1_n16 ,
         SubCellInst_LFInst_15_LFInst_1_n15 ,
         SubCellInst_LFInst_15_LFInst_1_n14 ,
         SubCellInst_LFInst_15_LFInst_1_n13 ,
         SubCellInst_LFInst_15_LFInst_1_n12 ,
         SubCellInst_LFInst_15_LFInst_1_n11 ,
         SubCellInst_LFInst_15_LFInst_1_n10 ,
         SubCellInst_LFInst_15_LFInst_0_n6 ,
         SubCellInst_LFInst_15_LFInst_0_n5 ,
         SubCellInst_LFInst_15_LFInst_0_n4 , MCInst1_MC0_v0_2Inst_0_n2 ,
         MCInst1_MC0_v1_2Inst_0_n2 , MCInst1_MC0_v2_3Inst_0_n4 ,
         MCInst1_MC0_v2_3Inst_0_n3 , MCInst1_MC0_v3_3Inst_0_n2 ,
         MCInst1_MC0_v0_2Inst_1_n2 , MCInst1_MC0_v2_1Inst_1_n2 ,
         MCInst1_MC0_v2_2Inst_1_n4 , MCInst1_MC0_v2_2Inst_1_n3 ,
         MCInst1_MC0_v3_3Inst_1_n2 , MCInst1_MC0_v1_1Inst_2_n2 ,
         MCInst1_MC0_v1_2Inst_2_n2 , MCInst1_MC0_v2_1Inst_2_n2 ,
         MCInst1_MC0_v2_2Inst_2_n2 , MCInst1_MC0_v3_1Inst_2_n2 ,
         MCInst1_MC0_v1_2Inst_3_n4 , MCInst1_MC0_v1_2Inst_3_n3 ,
         MCInst1_MC0_v2_2Inst_3_n2 , MCInst1_MC0_v2_3Inst_3_n2 ,
         MCInst1_MC0_r0Inst_XORInst_0_0_n5 ,
         MCInst1_MC0_r0Inst_XORInst_0_0_n4 ,
         MCInst1_MC0_r0Inst_XORInst_0_1_n5 ,
         MCInst1_MC0_r0Inst_XORInst_0_1_n4 ,
         MCInst1_MC0_r0Inst_XORInst_0_2_n5 ,
         MCInst1_MC0_r0Inst_XORInst_0_2_n4 ,
         MCInst1_MC0_r0Inst_XORInst_0_3_n5 ,
         MCInst1_MC0_r0Inst_XORInst_0_3_n4 ,
         MCInst1_MC0_r1Inst_XORInst_0_0_n5 ,
         MCInst1_MC0_r1Inst_XORInst_0_0_n4 ,
         MCInst1_MC0_r1Inst_XORInst_0_1_n5 ,
         MCInst1_MC0_r1Inst_XORInst_0_1_n4 ,
         MCInst1_MC0_r1Inst_XORInst_0_2_n5 ,
         MCInst1_MC0_r1Inst_XORInst_0_2_n4 ,
         MCInst1_MC0_r1Inst_XORInst_0_3_n5 ,
         MCInst1_MC0_r1Inst_XORInst_0_3_n4 ,
         MCInst1_MC0_r2Inst_XORInst_0_0_n5 ,
         MCInst1_MC0_r2Inst_XORInst_0_0_n4 ,
         MCInst1_MC0_r2Inst_XORInst_0_1_n5 ,
         MCInst1_MC0_r2Inst_XORInst_0_1_n4 ,
         MCInst1_MC0_r2Inst_XORInst_0_2_n5 ,
         MCInst1_MC0_r2Inst_XORInst_0_2_n4 ,
         MCInst1_MC0_r2Inst_XORInst_0_3_n5 ,
         MCInst1_MC0_r2Inst_XORInst_0_3_n4 ,
         MCInst1_MC0_r3Inst_XORInst_0_0_n5 ,
         MCInst1_MC0_r3Inst_XORInst_0_0_n4 ,
         MCInst1_MC0_r3Inst_XORInst_0_1_n5 ,
         MCInst1_MC0_r3Inst_XORInst_0_1_n4 ,
         MCInst1_MC0_r3Inst_XORInst_0_2_n5 ,
         MCInst1_MC0_r3Inst_XORInst_0_2_n4 ,
         MCInst1_MC0_r3Inst_XORInst_0_3_n5 ,
         MCInst1_MC0_r3Inst_XORInst_0_3_n4 , MCInst1_MC1_v0_2Inst_0_n2 ,
         MCInst1_MC1_v1_2Inst_0_n2 , MCInst1_MC1_v2_3Inst_0_n4 ,
         MCInst1_MC1_v2_3Inst_0_n3 , MCInst1_MC1_v3_3Inst_0_n2 ,
         MCInst1_MC1_v0_2Inst_1_n2 , MCInst1_MC1_v2_1Inst_1_n2 ,
         MCInst1_MC1_v2_2Inst_1_n4 , MCInst1_MC1_v2_2Inst_1_n3 ,
         MCInst1_MC1_v3_3Inst_1_n2 , MCInst1_MC1_v1_1Inst_2_n2 ,
         MCInst1_MC1_v1_2Inst_2_n2 , MCInst1_MC1_v2_1Inst_2_n2 ,
         MCInst1_MC1_v2_2Inst_2_n2 , MCInst1_MC1_v3_1Inst_2_n2 ,
         MCInst1_MC1_v1_2Inst_3_n4 , MCInst1_MC1_v1_2Inst_3_n3 ,
         MCInst1_MC1_v2_2Inst_3_n2 , MCInst1_MC1_v2_3Inst_3_n2 ,
         MCInst1_MC1_r0Inst_XORInst_0_0_n5 ,
         MCInst1_MC1_r0Inst_XORInst_0_0_n4 ,
         MCInst1_MC1_r0Inst_XORInst_0_1_n5 ,
         MCInst1_MC1_r0Inst_XORInst_0_1_n4 ,
         MCInst1_MC1_r0Inst_XORInst_0_2_n5 ,
         MCInst1_MC1_r0Inst_XORInst_0_2_n4 ,
         MCInst1_MC1_r0Inst_XORInst_0_3_n5 ,
         MCInst1_MC1_r0Inst_XORInst_0_3_n4 ,
         MCInst1_MC1_r1Inst_XORInst_0_0_n5 ,
         MCInst1_MC1_r1Inst_XORInst_0_0_n4 ,
         MCInst1_MC1_r1Inst_XORInst_0_1_n5 ,
         MCInst1_MC1_r1Inst_XORInst_0_1_n4 ,
         MCInst1_MC1_r1Inst_XORInst_0_2_n5 ,
         MCInst1_MC1_r1Inst_XORInst_0_2_n4 ,
         MCInst1_MC1_r1Inst_XORInst_0_3_n5 ,
         MCInst1_MC1_r1Inst_XORInst_0_3_n4 ,
         MCInst1_MC1_r2Inst_XORInst_0_0_n5 ,
         MCInst1_MC1_r2Inst_XORInst_0_0_n4 ,
         MCInst1_MC1_r2Inst_XORInst_0_1_n5 ,
         MCInst1_MC1_r2Inst_XORInst_0_1_n4 ,
         MCInst1_MC1_r2Inst_XORInst_0_2_n5 ,
         MCInst1_MC1_r2Inst_XORInst_0_2_n4 ,
         MCInst1_MC1_r2Inst_XORInst_0_3_n5 ,
         MCInst1_MC1_r2Inst_XORInst_0_3_n4 ,
         MCInst1_MC1_r3Inst_XORInst_0_0_n5 ,
         MCInst1_MC1_r3Inst_XORInst_0_0_n4 ,
         MCInst1_MC1_r3Inst_XORInst_0_1_n5 ,
         MCInst1_MC1_r3Inst_XORInst_0_1_n4 ,
         MCInst1_MC1_r3Inst_XORInst_0_2_n5 ,
         MCInst1_MC1_r3Inst_XORInst_0_2_n4 ,
         MCInst1_MC1_r3Inst_XORInst_0_3_n5 ,
         MCInst1_MC1_r3Inst_XORInst_0_3_n4 , MCInst1_MC2_v0_2Inst_0_n2 ,
         MCInst1_MC2_v1_2Inst_0_n2 , MCInst1_MC2_v2_3Inst_0_n4 ,
         MCInst1_MC2_v2_3Inst_0_n3 , MCInst1_MC2_v3_3Inst_0_n2 ,
         MCInst1_MC2_v0_2Inst_1_n2 , MCInst1_MC2_v2_1Inst_1_n2 ,
         MCInst1_MC2_v2_2Inst_1_n4 , MCInst1_MC2_v2_2Inst_1_n3 ,
         MCInst1_MC2_v3_3Inst_1_n2 , MCInst1_MC2_v1_1Inst_2_n2 ,
         MCInst1_MC2_v1_2Inst_2_n2 , MCInst1_MC2_v2_1Inst_2_n2 ,
         MCInst1_MC2_v2_2Inst_2_n2 , MCInst1_MC2_v3_1Inst_2_n2 ,
         MCInst1_MC2_v1_2Inst_3_n4 , MCInst1_MC2_v1_2Inst_3_n3 ,
         MCInst1_MC2_v2_2Inst_3_n2 , MCInst1_MC2_v2_3Inst_3_n2 ,
         MCInst1_MC2_r0Inst_XORInst_0_0_n5 ,
         MCInst1_MC2_r0Inst_XORInst_0_0_n4 ,
         MCInst1_MC2_r0Inst_XORInst_0_1_n5 ,
         MCInst1_MC2_r0Inst_XORInst_0_1_n4 ,
         MCInst1_MC2_r0Inst_XORInst_0_2_n5 ,
         MCInst1_MC2_r0Inst_XORInst_0_2_n4 ,
         MCInst1_MC2_r0Inst_XORInst_0_3_n5 ,
         MCInst1_MC2_r0Inst_XORInst_0_3_n4 ,
         MCInst1_MC2_r1Inst_XORInst_0_0_n5 ,
         MCInst1_MC2_r1Inst_XORInst_0_0_n4 ,
         MCInst1_MC2_r1Inst_XORInst_0_1_n5 ,
         MCInst1_MC2_r1Inst_XORInst_0_1_n4 ,
         MCInst1_MC2_r1Inst_XORInst_0_2_n5 ,
         MCInst1_MC2_r1Inst_XORInst_0_2_n4 ,
         MCInst1_MC2_r1Inst_XORInst_0_3_n5 ,
         MCInst1_MC2_r1Inst_XORInst_0_3_n4 ,
         MCInst1_MC2_r2Inst_XORInst_0_0_n5 ,
         MCInst1_MC2_r2Inst_XORInst_0_0_n4 ,
         MCInst1_MC2_r2Inst_XORInst_0_1_n5 ,
         MCInst1_MC2_r2Inst_XORInst_0_1_n4 ,
         MCInst1_MC2_r2Inst_XORInst_0_2_n5 ,
         MCInst1_MC2_r2Inst_XORInst_0_2_n4 ,
         MCInst1_MC2_r2Inst_XORInst_0_3_n5 ,
         MCInst1_MC2_r2Inst_XORInst_0_3_n4 ,
         MCInst1_MC2_r3Inst_XORInst_0_0_n5 ,
         MCInst1_MC2_r3Inst_XORInst_0_0_n4 ,
         MCInst1_MC2_r3Inst_XORInst_0_1_n5 ,
         MCInst1_MC2_r3Inst_XORInst_0_1_n4 ,
         MCInst1_MC2_r3Inst_XORInst_0_2_n5 ,
         MCInst1_MC2_r3Inst_XORInst_0_2_n4 ,
         MCInst1_MC2_r3Inst_XORInst_0_3_n5 ,
         MCInst1_MC2_r3Inst_XORInst_0_3_n4 , MCInst1_MC3_v0_2Inst_0_n2 ,
         MCInst1_MC3_v1_2Inst_0_n2 , MCInst1_MC3_v2_3Inst_0_n4 ,
         MCInst1_MC3_v2_3Inst_0_n3 , MCInst1_MC3_v3_3Inst_0_n2 ,
         MCInst1_MC3_v0_2Inst_1_n2 , MCInst1_MC3_v2_1Inst_1_n2 ,
         MCInst1_MC3_v2_2Inst_1_n4 , MCInst1_MC3_v2_2Inst_1_n3 ,
         MCInst1_MC3_v3_3Inst_1_n2 , MCInst1_MC3_v1_1Inst_2_n2 ,
         MCInst1_MC3_v1_2Inst_2_n2 , MCInst1_MC3_v2_1Inst_2_n2 ,
         MCInst1_MC3_v2_2Inst_2_n2 , MCInst1_MC3_v3_1Inst_2_n2 ,
         MCInst1_MC3_v1_2Inst_3_n4 , MCInst1_MC3_v1_2Inst_3_n3 ,
         MCInst1_MC3_v2_2Inst_3_n2 , MCInst1_MC3_v2_3Inst_3_n2 ,
         MCInst1_MC3_r0Inst_XORInst_0_0_n5 ,
         MCInst1_MC3_r0Inst_XORInst_0_0_n4 ,
         MCInst1_MC3_r0Inst_XORInst_0_1_n5 ,
         MCInst1_MC3_r0Inst_XORInst_0_1_n4 ,
         MCInst1_MC3_r0Inst_XORInst_0_2_n5 ,
         MCInst1_MC3_r0Inst_XORInst_0_2_n4 ,
         MCInst1_MC3_r0Inst_XORInst_0_3_n5 ,
         MCInst1_MC3_r0Inst_XORInst_0_3_n4 ,
         MCInst1_MC3_r1Inst_XORInst_0_0_n5 ,
         MCInst1_MC3_r1Inst_XORInst_0_0_n4 ,
         MCInst1_MC3_r1Inst_XORInst_0_1_n5 ,
         MCInst1_MC3_r1Inst_XORInst_0_1_n4 ,
         MCInst1_MC3_r1Inst_XORInst_0_2_n5 ,
         MCInst1_MC3_r1Inst_XORInst_0_2_n4 ,
         MCInst1_MC3_r1Inst_XORInst_0_3_n5 ,
         MCInst1_MC3_r1Inst_XORInst_0_3_n4 ,
         MCInst1_MC3_r2Inst_XORInst_0_0_n5 ,
         MCInst1_MC3_r2Inst_XORInst_0_0_n4 ,
         MCInst1_MC3_r2Inst_XORInst_0_1_n5 ,
         MCInst1_MC3_r2Inst_XORInst_0_1_n4 ,
         MCInst1_MC3_r2Inst_XORInst_0_2_n5 ,
         MCInst1_MC3_r2Inst_XORInst_0_2_n4 ,
         MCInst1_MC3_r2Inst_XORInst_0_3_n5 ,
         MCInst1_MC3_r2Inst_XORInst_0_3_n4 ,
         MCInst1_MC3_r3Inst_XORInst_0_0_n5 ,
         MCInst1_MC3_r3Inst_XORInst_0_0_n4 ,
         MCInst1_MC3_r3Inst_XORInst_0_1_n5 ,
         MCInst1_MC3_r3Inst_XORInst_0_1_n4 ,
         MCInst1_MC3_r3Inst_XORInst_0_2_n5 ,
         MCInst1_MC3_r3Inst_XORInst_0_2_n4 ,
         MCInst1_MC3_r3Inst_XORInst_0_3_n5 ,
         MCInst1_MC3_r3Inst_XORInst_0_3_n4 ;
  wire   [63:0] AddRoundKeyOutput;
  wire   [63:0] ShiftRowsOutput;
  wire   [3:0] MCInst1_MC0_v3_3 ;
  wire   [3:0] MCInst1_MC0_v3_2 ;
  wire   [3:0] MCInst1_MC0_v3_1 ;
  wire   [3:0] MCInst1_MC0_v3_0 ;
  wire   [3:0] MCInst1_MC0_v2_3 ;
  wire   [3:0] MCInst1_MC0_v2_2 ;
  wire   [3:0] MCInst1_MC0_v2_1 ;
  wire   [3:0] MCInst1_MC0_v2_0 ;
  wire   [3:0] MCInst1_MC0_v1_3 ;
  wire   [3:0] MCInst1_MC0_v1_2 ;
  wire   [3:0] MCInst1_MC0_v1_1 ;
  wire   [3:0] MCInst1_MC0_v0_3 ;
  wire   [3:0] MCInst1_MC0_v0_2 ;
  wire   [3:0] MCInst1_MC0_v0_1 ;
  wire   [3:0] MCInst1_MC0_v0_0 ;
  wire   [3:0] MCInst1_MC1_v3_3 ;
  wire   [3:0] MCInst1_MC1_v3_2 ;
  wire   [3:0] MCInst1_MC1_v3_1 ;
  wire   [3:0] MCInst1_MC1_v3_0 ;
  wire   [3:0] MCInst1_MC1_v2_3 ;
  wire   [3:0] MCInst1_MC1_v2_2 ;
  wire   [3:0] MCInst1_MC1_v2_1 ;
  wire   [3:0] MCInst1_MC1_v2_0 ;
  wire   [3:0] MCInst1_MC1_v1_3 ;
  wire   [3:0] MCInst1_MC1_v1_2 ;
  wire   [3:0] MCInst1_MC1_v1_1 ;
  wire   [3:0] MCInst1_MC1_v0_3 ;
  wire   [3:0] MCInst1_MC1_v0_2 ;
  wire   [3:0] MCInst1_MC1_v0_1 ;
  wire   [3:0] MCInst1_MC1_v0_0 ;
  wire   [3:0] MCInst1_MC2_v3_3 ;
  wire   [3:0] MCInst1_MC2_v3_2 ;
  wire   [3:0] MCInst1_MC2_v3_1 ;
  wire   [3:0] MCInst1_MC2_v3_0 ;
  wire   [3:0] MCInst1_MC2_v2_3 ;
  wire   [3:0] MCInst1_MC2_v2_2 ;
  wire   [3:0] MCInst1_MC2_v2_1 ;
  wire   [3:0] MCInst1_MC2_v2_0 ;
  wire   [3:0] MCInst1_MC2_v1_3 ;
  wire   [3:0] MCInst1_MC2_v1_2 ;
  wire   [3:0] MCInst1_MC2_v1_1 ;
  wire   [3:0] MCInst1_MC2_v0_3 ;
  wire   [3:0] MCInst1_MC2_v0_2 ;
  wire   [3:0] MCInst1_MC2_v0_1 ;
  wire   [3:0] MCInst1_MC2_v0_0 ;
  wire   [3:0] MCInst1_MC3_v3_3 ;
  wire   [3:0] MCInst1_MC3_v3_2 ;
  wire   [3:0] MCInst1_MC3_v3_1 ;
  wire   [3:0] MCInst1_MC3_v3_0 ;
  wire   [3:0] MCInst1_MC3_v2_3 ;
  wire   [3:0] MCInst1_MC3_v2_2 ;
  wire   [3:0] MCInst1_MC3_v2_1 ;
  wire   [3:0] MCInst1_MC3_v2_0 ;
  wire   [3:0] MCInst1_MC3_v1_3 ;
  wire   [3:0] MCInst1_MC3_v1_2 ;
  wire   [3:0] MCInst1_MC3_v1_1 ;
  wire   [3:0] MCInst1_MC3_v0_3 ;
  wire   [3:0] MCInst1_MC3_v0_2 ;
  wire   [3:0] MCInst1_MC3_v0_1 ;
  wire   [3:0] MCInst1_MC3_v0_0 ;

  XOR2_X1 AddKeyXOR_XORInst_0_0_U1  ( .A(Plaintext[0]), .B(Key[0]), .Z(
        AddRoundKeyOutput[0]) );
  XOR2_X1 AddKeyXOR_XORInst_0_1_U1  ( .A(Plaintext[1]), .B(Key[1]), .Z(
        AddRoundKeyOutput[1]) );
  XOR2_X1 AddKeyXOR_XORInst_0_2_U1  ( .A(Plaintext[2]), .B(Key[2]), .Z(
        AddRoundKeyOutput[2]) );
  XOR2_X1 AddKeyXOR_XORInst_0_3_U1  ( .A(Plaintext[3]), .B(Key[3]), .Z(
        AddRoundKeyOutput[3]) );
  XOR2_X1 AddKeyXOR_XORInst_1_0_U1  ( .A(Plaintext[4]), .B(Key[4]), .Z(
        AddRoundKeyOutput[4]) );
  XOR2_X1 AddKeyXOR_XORInst_1_1_U1  ( .A(Plaintext[5]), .B(Key[5]), .Z(
        AddRoundKeyOutput[5]) );
  XOR2_X1 AddKeyXOR_XORInst_1_2_U1  ( .A(Plaintext[6]), .B(Key[6]), .Z(
        AddRoundKeyOutput[6]) );
  XOR2_X1 AddKeyXOR_XORInst_1_3_U1  ( .A(Plaintext[7]), .B(Key[7]), .Z(
        AddRoundKeyOutput[7]) );
  XOR2_X1 AddKeyXOR_XORInst_2_0_U1  ( .A(Plaintext[8]), .B(Key[8]), .Z(
        AddRoundKeyOutput[8]) );
  XOR2_X1 AddKeyXOR_XORInst_2_1_U1  ( .A(Plaintext[9]), .B(Key[9]), .Z(
        AddRoundKeyOutput[9]) );
  XOR2_X1 AddKeyXOR_XORInst_2_2_U1  ( .A(Plaintext[10]), .B(Key[10]), .Z(
        AddRoundKeyOutput[10]) );
  XOR2_X1 AddKeyXOR_XORInst_2_3_U1  ( .A(Plaintext[11]), .B(Key[11]), .Z(
        AddRoundKeyOutput[11]) );
  XOR2_X1 AddKeyXOR_XORInst_3_0_U1  ( .A(Plaintext[12]), .B(Key[12]), .Z(
        AddRoundKeyOutput[12]) );
  XOR2_X1 AddKeyXOR_XORInst_3_1_U1  ( .A(Plaintext[13]), .B(Key[13]), .Z(
        AddRoundKeyOutput[13]) );
  XOR2_X1 AddKeyXOR_XORInst_3_2_U1  ( .A(Plaintext[14]), .B(Key[14]), .Z(
        AddRoundKeyOutput[14]) );
  XOR2_X1 AddKeyXOR_XORInst_3_3_U1  ( .A(Plaintext[15]), .B(Key[15]), .Z(
        AddRoundKeyOutput[15]) );
  XOR2_X1 AddKeyXOR_XORInst_4_0_U1  ( .A(Plaintext[16]), .B(Key[16]), .Z(
        AddRoundKeyOutput[16]) );
  XOR2_X1 AddKeyXOR_XORInst_4_1_U1  ( .A(Plaintext[17]), .B(Key[17]), .Z(
        AddRoundKeyOutput[17]) );
  XOR2_X1 AddKeyXOR_XORInst_4_2_U1  ( .A(Plaintext[18]), .B(Key[18]), .Z(
        AddRoundKeyOutput[18]) );
  XOR2_X1 AddKeyXOR_XORInst_4_3_U1  ( .A(Plaintext[19]), .B(Key[19]), .Z(
        AddRoundKeyOutput[19]) );
  XOR2_X1 AddKeyXOR_XORInst_5_0_U1  ( .A(Plaintext[20]), .B(Key[20]), .Z(
        AddRoundKeyOutput[20]) );
  XOR2_X1 AddKeyXOR_XORInst_5_1_U1  ( .A(Plaintext[21]), .B(Key[21]), .Z(
        AddRoundKeyOutput[21]) );
  XOR2_X1 AddKeyXOR_XORInst_5_2_U1  ( .A(Plaintext[22]), .B(Key[22]), .Z(
        AddRoundKeyOutput[22]) );
  XOR2_X1 AddKeyXOR_XORInst_5_3_U1  ( .A(Plaintext[23]), .B(Key[23]), .Z(
        AddRoundKeyOutput[23]) );
  XOR2_X1 AddKeyXOR_XORInst_6_0_U1  ( .A(Plaintext[24]), .B(Key[24]), .Z(
        AddRoundKeyOutput[24]) );
  XOR2_X1 AddKeyXOR_XORInst_6_1_U1  ( .A(Plaintext[25]), .B(Key[25]), .Z(
        AddRoundKeyOutput[25]) );
  XOR2_X1 AddKeyXOR_XORInst_6_2_U1  ( .A(Plaintext[26]), .B(Key[26]), .Z(
        AddRoundKeyOutput[26]) );
  XOR2_X1 AddKeyXOR_XORInst_6_3_U1  ( .A(Plaintext[27]), .B(Key[27]), .Z(
        AddRoundKeyOutput[27]) );
  XOR2_X1 AddKeyXOR_XORInst_7_0_U1  ( .A(Plaintext[28]), .B(Key[28]), .Z(
        AddRoundKeyOutput[28]) );
  XOR2_X1 AddKeyXOR_XORInst_7_1_U1  ( .A(Plaintext[29]), .B(Key[29]), .Z(
        AddRoundKeyOutput[29]) );
  XOR2_X1 AddKeyXOR_XORInst_7_2_U1  ( .A(Plaintext[30]), .B(Key[30]), .Z(
        AddRoundKeyOutput[30]) );
  XOR2_X1 AddKeyXOR_XORInst_7_3_U1  ( .A(Plaintext[31]), .B(Key[31]), .Z(
        AddRoundKeyOutput[31]) );
  XOR2_X1 AddKeyXOR_XORInst_8_0_U1  ( .A(Plaintext[32]), .B(Key[32]), .Z(
        AddRoundKeyOutput[32]) );
  XOR2_X1 AddKeyXOR_XORInst_8_1_U1  ( .A(Plaintext[33]), .B(Key[33]), .Z(
        AddRoundKeyOutput[33]) );
  XOR2_X1 AddKeyXOR_XORInst_8_2_U1  ( .A(Plaintext[34]), .B(Key[34]), .Z(
        AddRoundKeyOutput[34]) );
  XOR2_X1 AddKeyXOR_XORInst_8_3_U1  ( .A(Plaintext[35]), .B(Key[35]), .Z(
        AddRoundKeyOutput[35]) );
  XOR2_X1 AddKeyXOR_XORInst_9_0_U1  ( .A(Plaintext[36]), .B(Key[36]), .Z(
        AddRoundKeyOutput[36]) );
  XOR2_X1 AddKeyXOR_XORInst_9_1_U1  ( .A(Plaintext[37]), .B(Key[37]), .Z(
        AddRoundKeyOutput[37]) );
  XOR2_X1 AddKeyXOR_XORInst_9_2_U1  ( .A(Plaintext[38]), .B(Key[38]), .Z(
        AddRoundKeyOutput[38]) );
  XOR2_X1 AddKeyXOR_XORInst_9_3_U1  ( .A(Plaintext[39]), .B(Key[39]), .Z(
        AddRoundKeyOutput[39]) );
  XOR2_X1 AddKeyXOR_XORInst_10_0_U1  ( .A(Plaintext[40]), .B(Key[40]), .Z(
        AddRoundKeyOutput[40]) );
  XOR2_X1 AddKeyXOR_XORInst_10_1_U1  ( .A(Plaintext[41]), .B(Key[41]), .Z(
        AddRoundKeyOutput[41]) );
  XOR2_X1 AddKeyXOR_XORInst_10_2_U1  ( .A(Plaintext[42]), .B(Key[42]), .Z(
        AddRoundKeyOutput[42]) );
  XOR2_X1 AddKeyXOR_XORInst_10_3_U1  ( .A(Plaintext[43]), .B(Key[43]), .Z(
        AddRoundKeyOutput[43]) );
  XOR2_X1 AddKeyXOR_XORInst_11_0_U1  ( .A(Plaintext[44]), .B(Key[44]), .Z(
        AddRoundKeyOutput[44]) );
  XOR2_X1 AddKeyXOR_XORInst_11_1_U1  ( .A(Plaintext[45]), .B(Key[45]), .Z(
        AddRoundKeyOutput[45]) );
  XOR2_X1 AddKeyXOR_XORInst_11_2_U1  ( .A(Plaintext[46]), .B(Key[46]), .Z(
        AddRoundKeyOutput[46]) );
  XOR2_X1 AddKeyXOR_XORInst_11_3_U1  ( .A(Plaintext[47]), .B(Key[47]), .Z(
        AddRoundKeyOutput[47]) );
  XOR2_X1 AddKeyXOR_XORInst_12_0_U1  ( .A(Plaintext[48]), .B(Key[48]), .Z(
        AddRoundKeyOutput[48]) );
  XOR2_X1 AddKeyXOR_XORInst_12_1_U1  ( .A(Plaintext[49]), .B(Key[49]), .Z(
        AddRoundKeyOutput[49]) );
  XOR2_X1 AddKeyXOR_XORInst_12_2_U1  ( .A(Plaintext[50]), .B(Key[50]), .Z(
        AddRoundKeyOutput[50]) );
  XOR2_X1 AddKeyXOR_XORInst_12_3_U1  ( .A(Plaintext[51]), .B(Key[51]), .Z(
        AddRoundKeyOutput[51]) );
  XOR2_X1 AddKeyXOR_XORInst_13_0_U1  ( .A(Plaintext[52]), .B(Key[52]), .Z(
        AddRoundKeyOutput[52]) );
  XOR2_X1 AddKeyXOR_XORInst_13_1_U1  ( .A(Plaintext[53]), .B(Key[53]), .Z(
        AddRoundKeyOutput[53]) );
  XOR2_X1 AddKeyXOR_XORInst_13_2_U1  ( .A(Plaintext[54]), .B(Key[54]), .Z(
        AddRoundKeyOutput[54]) );
  XOR2_X1 AddKeyXOR_XORInst_13_3_U1  ( .A(Plaintext[55]), .B(Key[55]), .Z(
        AddRoundKeyOutput[55]) );
  XOR2_X1 AddKeyXOR_XORInst_14_0_U1  ( .A(Plaintext[56]), .B(Key[56]), .Z(
        AddRoundKeyOutput[56]) );
  XOR2_X1 AddKeyXOR_XORInst_14_1_U1  ( .A(Plaintext[57]), .B(Key[57]), .Z(
        AddRoundKeyOutput[57]) );
  XOR2_X1 AddKeyXOR_XORInst_14_2_U1  ( .A(Plaintext[58]), .B(Key[58]), .Z(
        AddRoundKeyOutput[58]) );
  XOR2_X1 AddKeyXOR_XORInst_14_3_U1  ( .A(Plaintext[59]), .B(Key[59]), .Z(
        AddRoundKeyOutput[59]) );
  XOR2_X1 AddKeyXOR_XORInst_15_0_U1  ( .A(Plaintext[60]), .B(Key[60]), .Z(
        AddRoundKeyOutput[60]) );
  XOR2_X1 AddKeyXOR_XORInst_15_1_U1  ( .A(Plaintext[61]), .B(Key[61]), .Z(
        AddRoundKeyOutput[61]) );
  XOR2_X1 AddKeyXOR_XORInst_15_2_U1  ( .A(Plaintext[62]), .B(Key[62]), .Z(
        AddRoundKeyOutput[62]) );
  XOR2_X1 AddKeyXOR_XORInst_15_3_U1  ( .A(Plaintext[63]), .B(Key[63]), .Z(
        AddRoundKeyOutput[63]) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_3_U9  ( .A1(
        SubCellInst_LFInst_0_LFInst_3_n16 ), .A2(
        SubCellInst_LFInst_0_LFInst_3_n15 ), .ZN(MCInst1_MC0_v3_2 [2]) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_3_U8  ( .A1(AddRoundKeyOutput[1]), 
        .A2(SubCellInst_LFInst_0_LFInst_3_n14 ), .ZN(
        SubCellInst_LFInst_0_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst_LFInst_0_LFInst_3_U7  ( .A(AddRoundKeyOutput[3]), .B(
        AddRoundKeyOutput[2]), .Z(SubCellInst_LFInst_0_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_3_U6  ( .A1(
        SubCellInst_LFInst_0_LFInst_3_n13 ), .A2(
        SubCellInst_LFInst_0_LFInst_3_n12 ), .ZN(
        SubCellInst_LFInst_0_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_3_U5  ( .A1(AddRoundKeyOutput[0]), 
        .A2(AddRoundKeyOutput[2]), .ZN(SubCellInst_LFInst_0_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst_LFInst_0_LFInst_3_U4  ( .A(AddRoundKeyOutput[0]), .B(
        SubCellInst_LFInst_0_LFInst_3_n11 ), .ZN(
        SubCellInst_LFInst_0_LFInst_3_n13 ) );
  OR2_X1 SubCellInst_LFInst_0_LFInst_3_U3  ( .A1(AddRoundKeyOutput[3]), .A2(
        AddRoundKeyOutput[1]), .ZN(SubCellInst_LFInst_0_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_2_U11  ( .A1(
        SubCellInst_LFInst_0_LFInst_2_n22 ), .A2(
        SubCellInst_LFInst_0_LFInst_2_n21 ), .ZN(MCInst1_MC0_v3_0 [3]) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_2_U10  ( .A1(AddRoundKeyOutput[2]), 
        .A2(SubCellInst_LFInst_0_LFInst_2_n20 ), .ZN(
        SubCellInst_LFInst_0_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst_LFInst_0_LFInst_2_U9  ( .A1(AddRoundKeyOutput[1]), .A2(
        SubCellInst_LFInst_0_LFInst_2_n19 ), .ZN(
        SubCellInst_LFInst_0_LFInst_2_n20 ) );
  INV_X1 SubCellInst_LFInst_0_LFInst_2_U8  ( .A(AddRoundKeyOutput[3]), .ZN(
        SubCellInst_LFInst_0_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_2_U7  ( .A1(
        SubCellInst_LFInst_0_LFInst_2_n18 ), .A2(
        SubCellInst_LFInst_0_LFInst_2_n17 ), .ZN(
        SubCellInst_LFInst_0_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst_LFInst_0_LFInst_2_U6  ( .A(
        SubCellInst_LFInst_0_LFInst_2_n16 ), .B(AddRoundKeyOutput[2]), .Z(
        SubCellInst_LFInst_0_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_2_U5  ( .A1(AddRoundKeyOutput[0]), 
        .A2(AddRoundKeyOutput[1]), .ZN(SubCellInst_LFInst_0_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_2_U4  ( .A1(
        SubCellInst_LFInst_0_LFInst_2_n15 ), .A2(AddRoundKeyOutput[3]), .ZN(
        SubCellInst_LFInst_0_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst_LFInst_0_LFInst_2_U3  ( .A(AddRoundKeyOutput[0]), .B(
        AddRoundKeyOutput[1]), .ZN(SubCellInst_LFInst_0_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_1_U12  ( .A1(
        SubCellInst_LFInst_0_LFInst_1_n18 ), .A2(
        SubCellInst_LFInst_0_LFInst_1_n17 ), .ZN(MCInst1_MC0_v3_0 [2]) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_1_U11  ( .A1(AddRoundKeyOutput[1]), 
        .A2(SubCellInst_LFInst_0_LFInst_1_n16 ), .ZN(
        SubCellInst_LFInst_0_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst_LFInst_0_LFInst_1_U10  ( .A1(AddRoundKeyOutput[3]), 
        .A2(SubCellInst_LFInst_0_LFInst_1_n15 ), .ZN(
        SubCellInst_LFInst_0_LFInst_1_n16 ) );
  AND2_X1 SubCellInst_LFInst_0_LFInst_1_U9  ( .A1(AddRoundKeyOutput[0]), .A2(
        AddRoundKeyOutput[2]), .ZN(SubCellInst_LFInst_0_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_1_U8  ( .A1(AddRoundKeyOutput[3]), 
        .A2(SubCellInst_LFInst_0_LFInst_1_n14 ), .ZN(
        SubCellInst_LFInst_0_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_1_U7  ( .A1(
        SubCellInst_LFInst_0_LFInst_1_n13 ), .A2(
        SubCellInst_LFInst_0_LFInst_1_n12 ), .ZN(
        SubCellInst_LFInst_0_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_1_U6  ( .A1(AddRoundKeyOutput[0]), 
        .A2(AddRoundKeyOutput[2]), .ZN(SubCellInst_LFInst_0_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_1_U5  ( .A1(
        SubCellInst_LFInst_0_LFInst_1_n11 ), .A2(
        SubCellInst_LFInst_0_LFInst_1_n10 ), .ZN(
        SubCellInst_LFInst_0_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_1_U4  ( .A1(AddRoundKeyOutput[0]), 
        .A2(AddRoundKeyOutput[1]), .ZN(SubCellInst_LFInst_0_LFInst_1_n10 ) );
  INV_X1 SubCellInst_LFInst_0_LFInst_1_U3  ( .A(AddRoundKeyOutput[2]), .ZN(
        SubCellInst_LFInst_0_LFInst_1_n11 ) );
  XNOR2_X1 SubCellInst_LFInst_0_LFInst_0_U6  ( .A(
        SubCellInst_LFInst_0_LFInst_0_n6 ), .B(
        SubCellInst_LFInst_0_LFInst_0_n5 ), .ZN(MCInst1_MC0_v3_2 [3]) );
  NAND2_X1 SubCellInst_LFInst_0_LFInst_0_U5  ( .A1(AddRoundKeyOutput[2]), 
        .A2(SubCellInst_LFInst_0_LFInst_0_n4 ), .ZN(
        SubCellInst_LFInst_0_LFInst_0_n5 ) );
  INV_X1 SubCellInst_LFInst_0_LFInst_0_U4  ( .A(AddRoundKeyOutput[1]), .ZN(
        SubCellInst_LFInst_0_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst_LFInst_0_LFInst_0_U3  ( .A(AddRoundKeyOutput[0]), .B(
        AddRoundKeyOutput[3]), .Z(SubCellInst_LFInst_0_LFInst_0_n6 ) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_3_U9  ( .A1(
        SubCellInst_LFInst_1_LFInst_3_n16 ), .A2(
        SubCellInst_LFInst_1_LFInst_3_n15 ), .ZN(MCInst1_MC3_v3_2 [2]) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_3_U8  ( .A1(AddRoundKeyOutput[5]), 
        .A2(SubCellInst_LFInst_1_LFInst_3_n14 ), .ZN(
        SubCellInst_LFInst_1_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst_LFInst_1_LFInst_3_U7  ( .A(AddRoundKeyOutput[7]), .B(
        AddRoundKeyOutput[6]), .Z(SubCellInst_LFInst_1_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_3_U6  ( .A1(
        SubCellInst_LFInst_1_LFInst_3_n13 ), .A2(
        SubCellInst_LFInst_1_LFInst_3_n12 ), .ZN(
        SubCellInst_LFInst_1_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_3_U5  ( .A1(AddRoundKeyOutput[4]), 
        .A2(AddRoundKeyOutput[6]), .ZN(SubCellInst_LFInst_1_LFInst_3_n12 ) );
  XNOR2_X1 SubCellInst_LFInst_1_LFInst_3_U4  ( .A(AddRoundKeyOutput[4]), .B(
        SubCellInst_LFInst_1_LFInst_3_n11 ), .ZN(
        SubCellInst_LFInst_1_LFInst_3_n13 ) );
  OR2_X1 SubCellInst_LFInst_1_LFInst_3_U3  ( .A1(AddRoundKeyOutput[7]), .A2(
        AddRoundKeyOutput[5]), .ZN(SubCellInst_LFInst_1_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_2_U11  ( .A1(
        SubCellInst_LFInst_1_LFInst_2_n22 ), .A2(
        SubCellInst_LFInst_1_LFInst_2_n21 ), .ZN(MCInst1_MC3_v3_0 [3]) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_2_U10  ( .A1(AddRoundKeyOutput[6]), 
        .A2(SubCellInst_LFInst_1_LFInst_2_n20 ), .ZN(
        SubCellInst_LFInst_1_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst_LFInst_1_LFInst_2_U9  ( .A1(AddRoundKeyOutput[5]), .A2(
        SubCellInst_LFInst_1_LFInst_2_n19 ), .ZN(
        SubCellInst_LFInst_1_LFInst_2_n20 ) );
  INV_X1 SubCellInst_LFInst_1_LFInst_2_U8  ( .A(AddRoundKeyOutput[7]), .ZN(
        SubCellInst_LFInst_1_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_2_U7  ( .A1(
        SubCellInst_LFInst_1_LFInst_2_n18 ), .A2(
        SubCellInst_LFInst_1_LFInst_2_n17 ), .ZN(
        SubCellInst_LFInst_1_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst_LFInst_1_LFInst_2_U6  ( .A(
        SubCellInst_LFInst_1_LFInst_2_n16 ), .B(AddRoundKeyOutput[6]), .Z(
        SubCellInst_LFInst_1_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_2_U5  ( .A1(AddRoundKeyOutput[4]), 
        .A2(AddRoundKeyOutput[5]), .ZN(SubCellInst_LFInst_1_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_2_U4  ( .A1(
        SubCellInst_LFInst_1_LFInst_2_n15 ), .A2(AddRoundKeyOutput[7]), .ZN(
        SubCellInst_LFInst_1_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst_LFInst_1_LFInst_2_U3  ( .A(AddRoundKeyOutput[4]), .B(
        AddRoundKeyOutput[5]), .ZN(SubCellInst_LFInst_1_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_1_U12  ( .A1(
        SubCellInst_LFInst_1_LFInst_1_n18 ), .A2(
        SubCellInst_LFInst_1_LFInst_1_n17 ), .ZN(MCInst1_MC3_v3_0 [2]) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_1_U11  ( .A1(AddRoundKeyOutput[5]), 
        .A2(SubCellInst_LFInst_1_LFInst_1_n16 ), .ZN(
        SubCellInst_LFInst_1_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst_LFInst_1_LFInst_1_U10  ( .A1(AddRoundKeyOutput[7]), 
        .A2(SubCellInst_LFInst_1_LFInst_1_n15 ), .ZN(
        SubCellInst_LFInst_1_LFInst_1_n16 ) );
  AND2_X1 SubCellInst_LFInst_1_LFInst_1_U9  ( .A1(AddRoundKeyOutput[4]), .A2(
        AddRoundKeyOutput[6]), .ZN(SubCellInst_LFInst_1_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_1_U8  ( .A1(AddRoundKeyOutput[7]), 
        .A2(SubCellInst_LFInst_1_LFInst_1_n14 ), .ZN(
        SubCellInst_LFInst_1_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_1_U7  ( .A1(
        SubCellInst_LFInst_1_LFInst_1_n13 ), .A2(
        SubCellInst_LFInst_1_LFInst_1_n12 ), .ZN(
        SubCellInst_LFInst_1_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_1_U6  ( .A1(AddRoundKeyOutput[4]), 
        .A2(AddRoundKeyOutput[6]), .ZN(SubCellInst_LFInst_1_LFInst_1_n12 ) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_1_U5  ( .A1(
        SubCellInst_LFInst_1_LFInst_1_n11 ), .A2(
        SubCellInst_LFInst_1_LFInst_1_n10 ), .ZN(
        SubCellInst_LFInst_1_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_1_U4  ( .A1(AddRoundKeyOutput[4]), 
        .A2(AddRoundKeyOutput[5]), .ZN(SubCellInst_LFInst_1_LFInst_1_n10 ) );
  INV_X1 SubCellInst_LFInst_1_LFInst_1_U3  ( .A(AddRoundKeyOutput[6]), .ZN(
        SubCellInst_LFInst_1_LFInst_1_n11 ) );
  XNOR2_X1 SubCellInst_LFInst_1_LFInst_0_U6  ( .A(
        SubCellInst_LFInst_1_LFInst_0_n6 ), .B(
        SubCellInst_LFInst_1_LFInst_0_n5 ), .ZN(MCInst1_MC3_v3_2 [3]) );
  NAND2_X1 SubCellInst_LFInst_1_LFInst_0_U5  ( .A1(AddRoundKeyOutput[6]), 
        .A2(SubCellInst_LFInst_1_LFInst_0_n4 ), .ZN(
        SubCellInst_LFInst_1_LFInst_0_n5 ) );
  INV_X1 SubCellInst_LFInst_1_LFInst_0_U4  ( .A(AddRoundKeyOutput[5]), .ZN(
        SubCellInst_LFInst_1_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst_LFInst_1_LFInst_0_U3  ( .A(AddRoundKeyOutput[4]), .B(
        AddRoundKeyOutput[7]), .Z(SubCellInst_LFInst_1_LFInst_0_n6 ) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_3_U9  ( .A1(
        SubCellInst_LFInst_2_LFInst_3_n16 ), .A2(
        SubCellInst_LFInst_2_LFInst_3_n15 ), .ZN(MCInst1_MC2_v3_2 [2]) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_3_U8  ( .A1(AddRoundKeyOutput[9]), 
        .A2(SubCellInst_LFInst_2_LFInst_3_n14 ), .ZN(
        SubCellInst_LFInst_2_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst_LFInst_2_LFInst_3_U7  ( .A(AddRoundKeyOutput[11]), .B(
        AddRoundKeyOutput[10]), .Z(SubCellInst_LFInst_2_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_3_U6  ( .A1(
        SubCellInst_LFInst_2_LFInst_3_n13 ), .A2(
        SubCellInst_LFInst_2_LFInst_3_n12 ), .ZN(
        SubCellInst_LFInst_2_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_3_U5  ( .A1(AddRoundKeyOutput[8]), 
        .A2(AddRoundKeyOutput[10]), .ZN(SubCellInst_LFInst_2_LFInst_3_n12 )
         );
  XNOR2_X1 SubCellInst_LFInst_2_LFInst_3_U4  ( .A(AddRoundKeyOutput[8]), .B(
        SubCellInst_LFInst_2_LFInst_3_n11 ), .ZN(
        SubCellInst_LFInst_2_LFInst_3_n13 ) );
  OR2_X1 SubCellInst_LFInst_2_LFInst_3_U3  ( .A1(AddRoundKeyOutput[11]), .A2(
        AddRoundKeyOutput[9]), .ZN(SubCellInst_LFInst_2_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_2_U11  ( .A1(
        SubCellInst_LFInst_2_LFInst_2_n22 ), .A2(
        SubCellInst_LFInst_2_LFInst_2_n21 ), .ZN(MCInst1_MC2_v3_0 [3]) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_2_U10  ( .A1(AddRoundKeyOutput[10]), 
        .A2(SubCellInst_LFInst_2_LFInst_2_n20 ), .ZN(
        SubCellInst_LFInst_2_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst_LFInst_2_LFInst_2_U9  ( .A1(AddRoundKeyOutput[9]), .A2(
        SubCellInst_LFInst_2_LFInst_2_n19 ), .ZN(
        SubCellInst_LFInst_2_LFInst_2_n20 ) );
  INV_X1 SubCellInst_LFInst_2_LFInst_2_U8  ( .A(AddRoundKeyOutput[11]), .ZN(
        SubCellInst_LFInst_2_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_2_U7  ( .A1(
        SubCellInst_LFInst_2_LFInst_2_n18 ), .A2(
        SubCellInst_LFInst_2_LFInst_2_n17 ), .ZN(
        SubCellInst_LFInst_2_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst_LFInst_2_LFInst_2_U6  ( .A(
        SubCellInst_LFInst_2_LFInst_2_n16 ), .B(AddRoundKeyOutput[10]), .Z(
        SubCellInst_LFInst_2_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_2_U5  ( .A1(AddRoundKeyOutput[8]), 
        .A2(AddRoundKeyOutput[9]), .ZN(SubCellInst_LFInst_2_LFInst_2_n16 ) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_2_U4  ( .A1(
        SubCellInst_LFInst_2_LFInst_2_n15 ), .A2(AddRoundKeyOutput[11]), .ZN(
        SubCellInst_LFInst_2_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst_LFInst_2_LFInst_2_U3  ( .A(AddRoundKeyOutput[8]), .B(
        AddRoundKeyOutput[9]), .ZN(SubCellInst_LFInst_2_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_1_U12  ( .A1(
        SubCellInst_LFInst_2_LFInst_1_n18 ), .A2(
        SubCellInst_LFInst_2_LFInst_1_n17 ), .ZN(MCInst1_MC2_v3_0 [2]) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_1_U11  ( .A1(AddRoundKeyOutput[9]), 
        .A2(SubCellInst_LFInst_2_LFInst_1_n16 ), .ZN(
        SubCellInst_LFInst_2_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst_LFInst_2_LFInst_1_U10  ( .A1(AddRoundKeyOutput[11]), 
        .A2(SubCellInst_LFInst_2_LFInst_1_n15 ), .ZN(
        SubCellInst_LFInst_2_LFInst_1_n16 ) );
  AND2_X1 SubCellInst_LFInst_2_LFInst_1_U9  ( .A1(AddRoundKeyOutput[8]), .A2(
        AddRoundKeyOutput[10]), .ZN(SubCellInst_LFInst_2_LFInst_1_n15 ) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_1_U8  ( .A1(AddRoundKeyOutput[11]), 
        .A2(SubCellInst_LFInst_2_LFInst_1_n14 ), .ZN(
        SubCellInst_LFInst_2_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_1_U7  ( .A1(
        SubCellInst_LFInst_2_LFInst_1_n13 ), .A2(
        SubCellInst_LFInst_2_LFInst_1_n12 ), .ZN(
        SubCellInst_LFInst_2_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_1_U6  ( .A1(AddRoundKeyOutput[8]), 
        .A2(AddRoundKeyOutput[10]), .ZN(SubCellInst_LFInst_2_LFInst_1_n12 )
         );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_1_U5  ( .A1(
        SubCellInst_LFInst_2_LFInst_1_n11 ), .A2(
        SubCellInst_LFInst_2_LFInst_1_n10 ), .ZN(
        SubCellInst_LFInst_2_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_1_U4  ( .A1(AddRoundKeyOutput[8]), 
        .A2(AddRoundKeyOutput[9]), .ZN(SubCellInst_LFInst_2_LFInst_1_n10 ) );
  INV_X1 SubCellInst_LFInst_2_LFInst_1_U3  ( .A(AddRoundKeyOutput[10]), .ZN(
        SubCellInst_LFInst_2_LFInst_1_n11 ) );
  XNOR2_X1 SubCellInst_LFInst_2_LFInst_0_U6  ( .A(
        SubCellInst_LFInst_2_LFInst_0_n6 ), .B(
        SubCellInst_LFInst_2_LFInst_0_n5 ), .ZN(MCInst1_MC2_v3_2 [3]) );
  NAND2_X1 SubCellInst_LFInst_2_LFInst_0_U5  ( .A1(AddRoundKeyOutput[10]), 
        .A2(SubCellInst_LFInst_2_LFInst_0_n4 ), .ZN(
        SubCellInst_LFInst_2_LFInst_0_n5 ) );
  INV_X1 SubCellInst_LFInst_2_LFInst_0_U4  ( .A(AddRoundKeyOutput[9]), .ZN(
        SubCellInst_LFInst_2_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst_LFInst_2_LFInst_0_U3  ( .A(AddRoundKeyOutput[8]), .B(
        AddRoundKeyOutput[11]), .Z(SubCellInst_LFInst_2_LFInst_0_n6 ) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_3_U9  ( .A1(
        SubCellInst_LFInst_3_LFInst_3_n16 ), .A2(
        SubCellInst_LFInst_3_LFInst_3_n15 ), .ZN(MCInst1_MC1_v3_2 [2]) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_3_U8  ( .A1(AddRoundKeyOutput[13]), 
        .A2(SubCellInst_LFInst_3_LFInst_3_n14 ), .ZN(
        SubCellInst_LFInst_3_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst_LFInst_3_LFInst_3_U7  ( .A(AddRoundKeyOutput[15]), .B(
        AddRoundKeyOutput[14]), .Z(SubCellInst_LFInst_3_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_3_U6  ( .A1(
        SubCellInst_LFInst_3_LFInst_3_n13 ), .A2(
        SubCellInst_LFInst_3_LFInst_3_n12 ), .ZN(
        SubCellInst_LFInst_3_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_3_U5  ( .A1(AddRoundKeyOutput[12]), 
        .A2(AddRoundKeyOutput[14]), .ZN(SubCellInst_LFInst_3_LFInst_3_n12 )
         );
  XNOR2_X1 SubCellInst_LFInst_3_LFInst_3_U4  ( .A(AddRoundKeyOutput[12]), .B(
        SubCellInst_LFInst_3_LFInst_3_n11 ), .ZN(
        SubCellInst_LFInst_3_LFInst_3_n13 ) );
  OR2_X1 SubCellInst_LFInst_3_LFInst_3_U3  ( .A1(AddRoundKeyOutput[15]), .A2(
        AddRoundKeyOutput[13]), .ZN(SubCellInst_LFInst_3_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_2_U11  ( .A1(
        SubCellInst_LFInst_3_LFInst_2_n22 ), .A2(
        SubCellInst_LFInst_3_LFInst_2_n21 ), .ZN(MCInst1_MC1_v3_0 [3]) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_2_U10  ( .A1(AddRoundKeyOutput[14]), 
        .A2(SubCellInst_LFInst_3_LFInst_2_n20 ), .ZN(
        SubCellInst_LFInst_3_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst_LFInst_3_LFInst_2_U9  ( .A1(AddRoundKeyOutput[13]), 
        .A2(SubCellInst_LFInst_3_LFInst_2_n19 ), .ZN(
        SubCellInst_LFInst_3_LFInst_2_n20 ) );
  INV_X1 SubCellInst_LFInst_3_LFInst_2_U8  ( .A(AddRoundKeyOutput[15]), .ZN(
        SubCellInst_LFInst_3_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_2_U7  ( .A1(
        SubCellInst_LFInst_3_LFInst_2_n18 ), .A2(
        SubCellInst_LFInst_3_LFInst_2_n17 ), .ZN(
        SubCellInst_LFInst_3_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst_LFInst_3_LFInst_2_U6  ( .A(
        SubCellInst_LFInst_3_LFInst_2_n16 ), .B(AddRoundKeyOutput[14]), .Z(
        SubCellInst_LFInst_3_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_2_U5  ( .A1(AddRoundKeyOutput[12]), 
        .A2(AddRoundKeyOutput[13]), .ZN(SubCellInst_LFInst_3_LFInst_2_n16 )
         );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_2_U4  ( .A1(
        SubCellInst_LFInst_3_LFInst_2_n15 ), .A2(AddRoundKeyOutput[15]), .ZN(
        SubCellInst_LFInst_3_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst_LFInst_3_LFInst_2_U3  ( .A(AddRoundKeyOutput[12]), .B(
        AddRoundKeyOutput[13]), .ZN(SubCellInst_LFInst_3_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_1_U12  ( .A1(
        SubCellInst_LFInst_3_LFInst_1_n18 ), .A2(
        SubCellInst_LFInst_3_LFInst_1_n17 ), .ZN(MCInst1_MC1_v3_0 [2]) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_1_U11  ( .A1(AddRoundKeyOutput[13]), 
        .A2(SubCellInst_LFInst_3_LFInst_1_n16 ), .ZN(
        SubCellInst_LFInst_3_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst_LFInst_3_LFInst_1_U10  ( .A1(AddRoundKeyOutput[15]), 
        .A2(SubCellInst_LFInst_3_LFInst_1_n15 ), .ZN(
        SubCellInst_LFInst_3_LFInst_1_n16 ) );
  AND2_X1 SubCellInst_LFInst_3_LFInst_1_U9  ( .A1(AddRoundKeyOutput[12]), 
        .A2(AddRoundKeyOutput[14]), .ZN(SubCellInst_LFInst_3_LFInst_1_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_1_U8  ( .A1(AddRoundKeyOutput[15]), 
        .A2(SubCellInst_LFInst_3_LFInst_1_n14 ), .ZN(
        SubCellInst_LFInst_3_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_1_U7  ( .A1(
        SubCellInst_LFInst_3_LFInst_1_n13 ), .A2(
        SubCellInst_LFInst_3_LFInst_1_n12 ), .ZN(
        SubCellInst_LFInst_3_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_1_U6  ( .A1(AddRoundKeyOutput[12]), 
        .A2(AddRoundKeyOutput[14]), .ZN(SubCellInst_LFInst_3_LFInst_1_n12 )
         );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_1_U5  ( .A1(
        SubCellInst_LFInst_3_LFInst_1_n11 ), .A2(
        SubCellInst_LFInst_3_LFInst_1_n10 ), .ZN(
        SubCellInst_LFInst_3_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_1_U4  ( .A1(AddRoundKeyOutput[12]), 
        .A2(AddRoundKeyOutput[13]), .ZN(SubCellInst_LFInst_3_LFInst_1_n10 )
         );
  INV_X1 SubCellInst_LFInst_3_LFInst_1_U3  ( .A(AddRoundKeyOutput[14]), .ZN(
        SubCellInst_LFInst_3_LFInst_1_n11 ) );
  XNOR2_X1 SubCellInst_LFInst_3_LFInst_0_U6  ( .A(
        SubCellInst_LFInst_3_LFInst_0_n6 ), .B(
        SubCellInst_LFInst_3_LFInst_0_n5 ), .ZN(MCInst1_MC1_v3_2 [3]) );
  NAND2_X1 SubCellInst_LFInst_3_LFInst_0_U5  ( .A1(AddRoundKeyOutput[14]), 
        .A2(SubCellInst_LFInst_3_LFInst_0_n4 ), .ZN(
        SubCellInst_LFInst_3_LFInst_0_n5 ) );
  INV_X1 SubCellInst_LFInst_3_LFInst_0_U4  ( .A(AddRoundKeyOutput[13]), .ZN(
        SubCellInst_LFInst_3_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst_LFInst_3_LFInst_0_U3  ( .A(AddRoundKeyOutput[12]), .B(
        AddRoundKeyOutput[15]), .Z(SubCellInst_LFInst_3_LFInst_0_n6 ) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_3_U9  ( .A1(
        SubCellInst_LFInst_4_LFInst_3_n16 ), .A2(
        SubCellInst_LFInst_4_LFInst_3_n15 ), .ZN(MCInst1_MC1_v2_0 [0]) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_3_U8  ( .A1(AddRoundKeyOutput[17]), 
        .A2(SubCellInst_LFInst_4_LFInst_3_n14 ), .ZN(
        SubCellInst_LFInst_4_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst_LFInst_4_LFInst_3_U7  ( .A(AddRoundKeyOutput[19]), .B(
        AddRoundKeyOutput[18]), .Z(SubCellInst_LFInst_4_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_3_U6  ( .A1(
        SubCellInst_LFInst_4_LFInst_3_n13 ), .A2(
        SubCellInst_LFInst_4_LFInst_3_n12 ), .ZN(
        SubCellInst_LFInst_4_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_3_U5  ( .A1(AddRoundKeyOutput[16]), 
        .A2(AddRoundKeyOutput[18]), .ZN(SubCellInst_LFInst_4_LFInst_3_n12 )
         );
  XNOR2_X1 SubCellInst_LFInst_4_LFInst_3_U4  ( .A(AddRoundKeyOutput[16]), .B(
        SubCellInst_LFInst_4_LFInst_3_n11 ), .ZN(
        SubCellInst_LFInst_4_LFInst_3_n13 ) );
  OR2_X1 SubCellInst_LFInst_4_LFInst_3_U3  ( .A1(AddRoundKeyOutput[19]), .A2(
        AddRoundKeyOutput[17]), .ZN(SubCellInst_LFInst_4_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_2_U11  ( .A1(
        SubCellInst_LFInst_4_LFInst_2_n22 ), .A2(
        SubCellInst_LFInst_4_LFInst_2_n21 ), .ZN(MCInst1_MC1_v2_0 [3]) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_2_U10  ( .A1(AddRoundKeyOutput[18]), 
        .A2(SubCellInst_LFInst_4_LFInst_2_n20 ), .ZN(
        SubCellInst_LFInst_4_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst_LFInst_4_LFInst_2_U9  ( .A1(AddRoundKeyOutput[17]), 
        .A2(SubCellInst_LFInst_4_LFInst_2_n19 ), .ZN(
        SubCellInst_LFInst_4_LFInst_2_n20 ) );
  INV_X1 SubCellInst_LFInst_4_LFInst_2_U8  ( .A(AddRoundKeyOutput[19]), .ZN(
        SubCellInst_LFInst_4_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_2_U7  ( .A1(
        SubCellInst_LFInst_4_LFInst_2_n18 ), .A2(
        SubCellInst_LFInst_4_LFInst_2_n17 ), .ZN(
        SubCellInst_LFInst_4_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst_LFInst_4_LFInst_2_U6  ( .A(
        SubCellInst_LFInst_4_LFInst_2_n16 ), .B(AddRoundKeyOutput[18]), .Z(
        SubCellInst_LFInst_4_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_2_U5  ( .A1(AddRoundKeyOutput[16]), 
        .A2(AddRoundKeyOutput[17]), .ZN(SubCellInst_LFInst_4_LFInst_2_n16 )
         );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_2_U4  ( .A1(
        SubCellInst_LFInst_4_LFInst_2_n15 ), .A2(AddRoundKeyOutput[19]), .ZN(
        SubCellInst_LFInst_4_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst_LFInst_4_LFInst_2_U3  ( .A(AddRoundKeyOutput[16]), .B(
        AddRoundKeyOutput[17]), .ZN(SubCellInst_LFInst_4_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_1_U12  ( .A1(
        SubCellInst_LFInst_4_LFInst_1_n18 ), .A2(
        SubCellInst_LFInst_4_LFInst_1_n17 ), .ZN(MCInst1_MC1_v2_0 [2]) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_1_U11  ( .A1(AddRoundKeyOutput[17]), 
        .A2(SubCellInst_LFInst_4_LFInst_1_n16 ), .ZN(
        SubCellInst_LFInst_4_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst_LFInst_4_LFInst_1_U10  ( .A1(AddRoundKeyOutput[19]), 
        .A2(SubCellInst_LFInst_4_LFInst_1_n15 ), .ZN(
        SubCellInst_LFInst_4_LFInst_1_n16 ) );
  AND2_X1 SubCellInst_LFInst_4_LFInst_1_U9  ( .A1(AddRoundKeyOutput[16]), 
        .A2(AddRoundKeyOutput[18]), .ZN(SubCellInst_LFInst_4_LFInst_1_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_1_U8  ( .A1(AddRoundKeyOutput[19]), 
        .A2(SubCellInst_LFInst_4_LFInst_1_n14 ), .ZN(
        SubCellInst_LFInst_4_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_1_U7  ( .A1(
        SubCellInst_LFInst_4_LFInst_1_n13 ), .A2(
        SubCellInst_LFInst_4_LFInst_1_n12 ), .ZN(
        SubCellInst_LFInst_4_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_1_U6  ( .A1(AddRoundKeyOutput[16]), 
        .A2(AddRoundKeyOutput[18]), .ZN(SubCellInst_LFInst_4_LFInst_1_n12 )
         );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_1_U5  ( .A1(
        SubCellInst_LFInst_4_LFInst_1_n11 ), .A2(
        SubCellInst_LFInst_4_LFInst_1_n10 ), .ZN(
        SubCellInst_LFInst_4_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_1_U4  ( .A1(AddRoundKeyOutput[16]), 
        .A2(AddRoundKeyOutput[17]), .ZN(SubCellInst_LFInst_4_LFInst_1_n10 )
         );
  INV_X1 SubCellInst_LFInst_4_LFInst_1_U3  ( .A(AddRoundKeyOutput[18]), .ZN(
        SubCellInst_LFInst_4_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst_LFInst_4_LFInst_0_U6  ( .A1(AddRoundKeyOutput[18]), 
        .A2(SubCellInst_LFInst_4_LFInst_0_n4 ), .ZN(
        SubCellInst_LFInst_4_LFInst_0_n5 ) );
  INV_X1 SubCellInst_LFInst_4_LFInst_0_U5  ( .A(AddRoundKeyOutput[17]), .ZN(
        SubCellInst_LFInst_4_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst_LFInst_4_LFInst_0_U4  ( .A(AddRoundKeyOutput[16]), .B(
        AddRoundKeyOutput[19]), .Z(SubCellInst_LFInst_4_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst_LFInst_4_LFInst_0_U3  ( .A(
        SubCellInst_LFInst_4_LFInst_0_n6 ), .B(
        SubCellInst_LFInst_4_LFInst_0_n5 ), .ZN(MCInst1_MC1_v2_3 [1]) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_3_U9  ( .A1(
        SubCellInst_LFInst_5_LFInst_3_n16 ), .A2(
        SubCellInst_LFInst_5_LFInst_3_n15 ), .ZN(MCInst1_MC0_v2_0 [0]) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_3_U8  ( .A1(AddRoundKeyOutput[21]), 
        .A2(SubCellInst_LFInst_5_LFInst_3_n14 ), .ZN(
        SubCellInst_LFInst_5_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst_LFInst_5_LFInst_3_U7  ( .A(AddRoundKeyOutput[23]), .B(
        AddRoundKeyOutput[22]), .Z(SubCellInst_LFInst_5_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_3_U6  ( .A1(
        SubCellInst_LFInst_5_LFInst_3_n13 ), .A2(
        SubCellInst_LFInst_5_LFInst_3_n12 ), .ZN(
        SubCellInst_LFInst_5_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_3_U5  ( .A1(AddRoundKeyOutput[20]), 
        .A2(AddRoundKeyOutput[22]), .ZN(SubCellInst_LFInst_5_LFInst_3_n12 )
         );
  XNOR2_X1 SubCellInst_LFInst_5_LFInst_3_U4  ( .A(AddRoundKeyOutput[20]), .B(
        SubCellInst_LFInst_5_LFInst_3_n11 ), .ZN(
        SubCellInst_LFInst_5_LFInst_3_n13 ) );
  OR2_X1 SubCellInst_LFInst_5_LFInst_3_U3  ( .A1(AddRoundKeyOutput[23]), .A2(
        AddRoundKeyOutput[21]), .ZN(SubCellInst_LFInst_5_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_2_U11  ( .A1(
        SubCellInst_LFInst_5_LFInst_2_n22 ), .A2(
        SubCellInst_LFInst_5_LFInst_2_n21 ), .ZN(MCInst1_MC0_v2_0 [3]) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_2_U10  ( .A1(AddRoundKeyOutput[22]), 
        .A2(SubCellInst_LFInst_5_LFInst_2_n20 ), .ZN(
        SubCellInst_LFInst_5_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst_LFInst_5_LFInst_2_U9  ( .A1(AddRoundKeyOutput[21]), 
        .A2(SubCellInst_LFInst_5_LFInst_2_n19 ), .ZN(
        SubCellInst_LFInst_5_LFInst_2_n20 ) );
  INV_X1 SubCellInst_LFInst_5_LFInst_2_U8  ( .A(AddRoundKeyOutput[23]), .ZN(
        SubCellInst_LFInst_5_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_2_U7  ( .A1(
        SubCellInst_LFInst_5_LFInst_2_n18 ), .A2(
        SubCellInst_LFInst_5_LFInst_2_n17 ), .ZN(
        SubCellInst_LFInst_5_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst_LFInst_5_LFInst_2_U6  ( .A(
        SubCellInst_LFInst_5_LFInst_2_n16 ), .B(AddRoundKeyOutput[22]), .Z(
        SubCellInst_LFInst_5_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_2_U5  ( .A1(AddRoundKeyOutput[20]), 
        .A2(AddRoundKeyOutput[21]), .ZN(SubCellInst_LFInst_5_LFInst_2_n16 )
         );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_2_U4  ( .A1(
        SubCellInst_LFInst_5_LFInst_2_n15 ), .A2(AddRoundKeyOutput[23]), .ZN(
        SubCellInst_LFInst_5_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst_LFInst_5_LFInst_2_U3  ( .A(AddRoundKeyOutput[20]), .B(
        AddRoundKeyOutput[21]), .ZN(SubCellInst_LFInst_5_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_1_U12  ( .A1(
        SubCellInst_LFInst_5_LFInst_1_n18 ), .A2(
        SubCellInst_LFInst_5_LFInst_1_n17 ), .ZN(MCInst1_MC0_v2_0 [2]) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_1_U11  ( .A1(AddRoundKeyOutput[21]), 
        .A2(SubCellInst_LFInst_5_LFInst_1_n16 ), .ZN(
        SubCellInst_LFInst_5_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst_LFInst_5_LFInst_1_U10  ( .A1(AddRoundKeyOutput[23]), 
        .A2(SubCellInst_LFInst_5_LFInst_1_n15 ), .ZN(
        SubCellInst_LFInst_5_LFInst_1_n16 ) );
  AND2_X1 SubCellInst_LFInst_5_LFInst_1_U9  ( .A1(AddRoundKeyOutput[20]), 
        .A2(AddRoundKeyOutput[22]), .ZN(SubCellInst_LFInst_5_LFInst_1_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_1_U8  ( .A1(AddRoundKeyOutput[23]), 
        .A2(SubCellInst_LFInst_5_LFInst_1_n14 ), .ZN(
        SubCellInst_LFInst_5_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_1_U7  ( .A1(
        SubCellInst_LFInst_5_LFInst_1_n13 ), .A2(
        SubCellInst_LFInst_5_LFInst_1_n12 ), .ZN(
        SubCellInst_LFInst_5_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_1_U6  ( .A1(AddRoundKeyOutput[20]), 
        .A2(AddRoundKeyOutput[22]), .ZN(SubCellInst_LFInst_5_LFInst_1_n12 )
         );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_1_U5  ( .A1(
        SubCellInst_LFInst_5_LFInst_1_n11 ), .A2(
        SubCellInst_LFInst_5_LFInst_1_n10 ), .ZN(
        SubCellInst_LFInst_5_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_1_U4  ( .A1(AddRoundKeyOutput[20]), 
        .A2(AddRoundKeyOutput[21]), .ZN(SubCellInst_LFInst_5_LFInst_1_n10 )
         );
  INV_X1 SubCellInst_LFInst_5_LFInst_1_U3  ( .A(AddRoundKeyOutput[22]), .ZN(
        SubCellInst_LFInst_5_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst_LFInst_5_LFInst_0_U6  ( .A1(AddRoundKeyOutput[22]), 
        .A2(SubCellInst_LFInst_5_LFInst_0_n4 ), .ZN(
        SubCellInst_LFInst_5_LFInst_0_n5 ) );
  INV_X1 SubCellInst_LFInst_5_LFInst_0_U5  ( .A(AddRoundKeyOutput[21]), .ZN(
        SubCellInst_LFInst_5_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst_LFInst_5_LFInst_0_U4  ( .A(AddRoundKeyOutput[20]), .B(
        AddRoundKeyOutput[23]), .Z(SubCellInst_LFInst_5_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst_LFInst_5_LFInst_0_U3  ( .A(
        SubCellInst_LFInst_5_LFInst_0_n6 ), .B(
        SubCellInst_LFInst_5_LFInst_0_n5 ), .ZN(MCInst1_MC0_v2_3 [1]) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_3_U9  ( .A1(
        SubCellInst_LFInst_6_LFInst_3_n16 ), .A2(
        SubCellInst_LFInst_6_LFInst_3_n15 ), .ZN(MCInst1_MC3_v2_0 [0]) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_3_U8  ( .A1(AddRoundKeyOutput[25]), 
        .A2(SubCellInst_LFInst_6_LFInst_3_n14 ), .ZN(
        SubCellInst_LFInst_6_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst_LFInst_6_LFInst_3_U7  ( .A(AddRoundKeyOutput[27]), .B(
        AddRoundKeyOutput[26]), .Z(SubCellInst_LFInst_6_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_3_U6  ( .A1(
        SubCellInst_LFInst_6_LFInst_3_n13 ), .A2(
        SubCellInst_LFInst_6_LFInst_3_n12 ), .ZN(
        SubCellInst_LFInst_6_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_3_U5  ( .A1(AddRoundKeyOutput[24]), 
        .A2(AddRoundKeyOutput[26]), .ZN(SubCellInst_LFInst_6_LFInst_3_n12 )
         );
  XNOR2_X1 SubCellInst_LFInst_6_LFInst_3_U4  ( .A(AddRoundKeyOutput[24]), .B(
        SubCellInst_LFInst_6_LFInst_3_n11 ), .ZN(
        SubCellInst_LFInst_6_LFInst_3_n13 ) );
  OR2_X1 SubCellInst_LFInst_6_LFInst_3_U3  ( .A1(AddRoundKeyOutput[27]), .A2(
        AddRoundKeyOutput[25]), .ZN(SubCellInst_LFInst_6_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_2_U11  ( .A1(
        SubCellInst_LFInst_6_LFInst_2_n22 ), .A2(
        SubCellInst_LFInst_6_LFInst_2_n21 ), .ZN(MCInst1_MC3_v2_0 [3]) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_2_U10  ( .A1(AddRoundKeyOutput[26]), 
        .A2(SubCellInst_LFInst_6_LFInst_2_n20 ), .ZN(
        SubCellInst_LFInst_6_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst_LFInst_6_LFInst_2_U9  ( .A1(AddRoundKeyOutput[25]), 
        .A2(SubCellInst_LFInst_6_LFInst_2_n19 ), .ZN(
        SubCellInst_LFInst_6_LFInst_2_n20 ) );
  INV_X1 SubCellInst_LFInst_6_LFInst_2_U8  ( .A(AddRoundKeyOutput[27]), .ZN(
        SubCellInst_LFInst_6_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_2_U7  ( .A1(
        SubCellInst_LFInst_6_LFInst_2_n18 ), .A2(
        SubCellInst_LFInst_6_LFInst_2_n17 ), .ZN(
        SubCellInst_LFInst_6_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst_LFInst_6_LFInst_2_U6  ( .A(
        SubCellInst_LFInst_6_LFInst_2_n16 ), .B(AddRoundKeyOutput[26]), .Z(
        SubCellInst_LFInst_6_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_2_U5  ( .A1(AddRoundKeyOutput[24]), 
        .A2(AddRoundKeyOutput[25]), .ZN(SubCellInst_LFInst_6_LFInst_2_n16 )
         );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_2_U4  ( .A1(
        SubCellInst_LFInst_6_LFInst_2_n15 ), .A2(AddRoundKeyOutput[27]), .ZN(
        SubCellInst_LFInst_6_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst_LFInst_6_LFInst_2_U3  ( .A(AddRoundKeyOutput[24]), .B(
        AddRoundKeyOutput[25]), .ZN(SubCellInst_LFInst_6_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_1_U12  ( .A1(
        SubCellInst_LFInst_6_LFInst_1_n18 ), .A2(
        SubCellInst_LFInst_6_LFInst_1_n17 ), .ZN(MCInst1_MC3_v2_0 [2]) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_1_U11  ( .A1(AddRoundKeyOutput[25]), 
        .A2(SubCellInst_LFInst_6_LFInst_1_n16 ), .ZN(
        SubCellInst_LFInst_6_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst_LFInst_6_LFInst_1_U10  ( .A1(AddRoundKeyOutput[27]), 
        .A2(SubCellInst_LFInst_6_LFInst_1_n15 ), .ZN(
        SubCellInst_LFInst_6_LFInst_1_n16 ) );
  AND2_X1 SubCellInst_LFInst_6_LFInst_1_U9  ( .A1(AddRoundKeyOutput[24]), 
        .A2(AddRoundKeyOutput[26]), .ZN(SubCellInst_LFInst_6_LFInst_1_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_1_U8  ( .A1(AddRoundKeyOutput[27]), 
        .A2(SubCellInst_LFInst_6_LFInst_1_n14 ), .ZN(
        SubCellInst_LFInst_6_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_1_U7  ( .A1(
        SubCellInst_LFInst_6_LFInst_1_n13 ), .A2(
        SubCellInst_LFInst_6_LFInst_1_n12 ), .ZN(
        SubCellInst_LFInst_6_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_1_U6  ( .A1(AddRoundKeyOutput[24]), 
        .A2(AddRoundKeyOutput[26]), .ZN(SubCellInst_LFInst_6_LFInst_1_n12 )
         );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_1_U5  ( .A1(
        SubCellInst_LFInst_6_LFInst_1_n11 ), .A2(
        SubCellInst_LFInst_6_LFInst_1_n10 ), .ZN(
        SubCellInst_LFInst_6_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_1_U4  ( .A1(AddRoundKeyOutput[24]), 
        .A2(AddRoundKeyOutput[25]), .ZN(SubCellInst_LFInst_6_LFInst_1_n10 )
         );
  INV_X1 SubCellInst_LFInst_6_LFInst_1_U3  ( .A(AddRoundKeyOutput[26]), .ZN(
        SubCellInst_LFInst_6_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst_LFInst_6_LFInst_0_U6  ( .A1(AddRoundKeyOutput[26]), 
        .A2(SubCellInst_LFInst_6_LFInst_0_n4 ), .ZN(
        SubCellInst_LFInst_6_LFInst_0_n5 ) );
  INV_X1 SubCellInst_LFInst_6_LFInst_0_U5  ( .A(AddRoundKeyOutput[25]), .ZN(
        SubCellInst_LFInst_6_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst_LFInst_6_LFInst_0_U4  ( .A(AddRoundKeyOutput[24]), .B(
        AddRoundKeyOutput[27]), .Z(SubCellInst_LFInst_6_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst_LFInst_6_LFInst_0_U3  ( .A(
        SubCellInst_LFInst_6_LFInst_0_n6 ), .B(
        SubCellInst_LFInst_6_LFInst_0_n5 ), .ZN(MCInst1_MC3_v2_3 [1]) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_3_U9  ( .A1(
        SubCellInst_LFInst_7_LFInst_3_n16 ), .A2(
        SubCellInst_LFInst_7_LFInst_3_n15 ), .ZN(MCInst1_MC2_v2_0 [0]) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_3_U8  ( .A1(AddRoundKeyOutput[29]), 
        .A2(SubCellInst_LFInst_7_LFInst_3_n14 ), .ZN(
        SubCellInst_LFInst_7_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst_LFInst_7_LFInst_3_U7  ( .A(AddRoundKeyOutput[31]), .B(
        AddRoundKeyOutput[30]), .Z(SubCellInst_LFInst_7_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_3_U6  ( .A1(
        SubCellInst_LFInst_7_LFInst_3_n13 ), .A2(
        SubCellInst_LFInst_7_LFInst_3_n12 ), .ZN(
        SubCellInst_LFInst_7_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_3_U5  ( .A1(AddRoundKeyOutput[28]), 
        .A2(AddRoundKeyOutput[30]), .ZN(SubCellInst_LFInst_7_LFInst_3_n12 )
         );
  XNOR2_X1 SubCellInst_LFInst_7_LFInst_3_U4  ( .A(AddRoundKeyOutput[28]), .B(
        SubCellInst_LFInst_7_LFInst_3_n11 ), .ZN(
        SubCellInst_LFInst_7_LFInst_3_n13 ) );
  OR2_X1 SubCellInst_LFInst_7_LFInst_3_U3  ( .A1(AddRoundKeyOutput[31]), .A2(
        AddRoundKeyOutput[29]), .ZN(SubCellInst_LFInst_7_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_2_U11  ( .A1(
        SubCellInst_LFInst_7_LFInst_2_n22 ), .A2(
        SubCellInst_LFInst_7_LFInst_2_n21 ), .ZN(MCInst1_MC2_v2_0 [3]) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_2_U10  ( .A1(AddRoundKeyOutput[30]), 
        .A2(SubCellInst_LFInst_7_LFInst_2_n20 ), .ZN(
        SubCellInst_LFInst_7_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst_LFInst_7_LFInst_2_U9  ( .A1(AddRoundKeyOutput[29]), 
        .A2(SubCellInst_LFInst_7_LFInst_2_n19 ), .ZN(
        SubCellInst_LFInst_7_LFInst_2_n20 ) );
  INV_X1 SubCellInst_LFInst_7_LFInst_2_U8  ( .A(AddRoundKeyOutput[31]), .ZN(
        SubCellInst_LFInst_7_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_2_U7  ( .A1(
        SubCellInst_LFInst_7_LFInst_2_n18 ), .A2(
        SubCellInst_LFInst_7_LFInst_2_n17 ), .ZN(
        SubCellInst_LFInst_7_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst_LFInst_7_LFInst_2_U6  ( .A(
        SubCellInst_LFInst_7_LFInst_2_n16 ), .B(AddRoundKeyOutput[30]), .Z(
        SubCellInst_LFInst_7_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_2_U5  ( .A1(AddRoundKeyOutput[28]), 
        .A2(AddRoundKeyOutput[29]), .ZN(SubCellInst_LFInst_7_LFInst_2_n16 )
         );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_2_U4  ( .A1(
        SubCellInst_LFInst_7_LFInst_2_n15 ), .A2(AddRoundKeyOutput[31]), .ZN(
        SubCellInst_LFInst_7_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst_LFInst_7_LFInst_2_U3  ( .A(AddRoundKeyOutput[28]), .B(
        AddRoundKeyOutput[29]), .ZN(SubCellInst_LFInst_7_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_1_U12  ( .A1(
        SubCellInst_LFInst_7_LFInst_1_n18 ), .A2(
        SubCellInst_LFInst_7_LFInst_1_n17 ), .ZN(MCInst1_MC2_v2_0 [2]) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_1_U11  ( .A1(AddRoundKeyOutput[29]), 
        .A2(SubCellInst_LFInst_7_LFInst_1_n16 ), .ZN(
        SubCellInst_LFInst_7_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst_LFInst_7_LFInst_1_U10  ( .A1(AddRoundKeyOutput[31]), 
        .A2(SubCellInst_LFInst_7_LFInst_1_n15 ), .ZN(
        SubCellInst_LFInst_7_LFInst_1_n16 ) );
  AND2_X1 SubCellInst_LFInst_7_LFInst_1_U9  ( .A1(AddRoundKeyOutput[28]), 
        .A2(AddRoundKeyOutput[30]), .ZN(SubCellInst_LFInst_7_LFInst_1_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_1_U8  ( .A1(AddRoundKeyOutput[31]), 
        .A2(SubCellInst_LFInst_7_LFInst_1_n14 ), .ZN(
        SubCellInst_LFInst_7_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_1_U7  ( .A1(
        SubCellInst_LFInst_7_LFInst_1_n13 ), .A2(
        SubCellInst_LFInst_7_LFInst_1_n12 ), .ZN(
        SubCellInst_LFInst_7_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_1_U6  ( .A1(AddRoundKeyOutput[28]), 
        .A2(AddRoundKeyOutput[30]), .ZN(SubCellInst_LFInst_7_LFInst_1_n12 )
         );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_1_U5  ( .A1(
        SubCellInst_LFInst_7_LFInst_1_n11 ), .A2(
        SubCellInst_LFInst_7_LFInst_1_n10 ), .ZN(
        SubCellInst_LFInst_7_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_1_U4  ( .A1(AddRoundKeyOutput[28]), 
        .A2(AddRoundKeyOutput[29]), .ZN(SubCellInst_LFInst_7_LFInst_1_n10 )
         );
  INV_X1 SubCellInst_LFInst_7_LFInst_1_U3  ( .A(AddRoundKeyOutput[30]), .ZN(
        SubCellInst_LFInst_7_LFInst_1_n11 ) );
  NAND2_X1 SubCellInst_LFInst_7_LFInst_0_U6  ( .A1(AddRoundKeyOutput[30]), 
        .A2(SubCellInst_LFInst_7_LFInst_0_n4 ), .ZN(
        SubCellInst_LFInst_7_LFInst_0_n5 ) );
  INV_X1 SubCellInst_LFInst_7_LFInst_0_U5  ( .A(AddRoundKeyOutput[29]), .ZN(
        SubCellInst_LFInst_7_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst_LFInst_7_LFInst_0_U4  ( .A(AddRoundKeyOutput[28]), .B(
        AddRoundKeyOutput[31]), .Z(SubCellInst_LFInst_7_LFInst_0_n6 ) );
  XNOR2_X2 SubCellInst_LFInst_7_LFInst_0_U3  ( .A(
        SubCellInst_LFInst_7_LFInst_0_n6 ), .B(
        SubCellInst_LFInst_7_LFInst_0_n5 ), .ZN(MCInst1_MC2_v2_3 [1]) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_3_U9  ( .A1(
        SubCellInst_LFInst_8_LFInst_3_n16 ), .A2(
        SubCellInst_LFInst_8_LFInst_3_n15 ), .ZN(MCInst1_MC2_v1_3 [0]) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_3_U8  ( .A1(AddRoundKeyOutput[33]), 
        .A2(SubCellInst_LFInst_8_LFInst_3_n14 ), .ZN(
        SubCellInst_LFInst_8_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst_LFInst_8_LFInst_3_U7  ( .A(AddRoundKeyOutput[35]), .B(
        AddRoundKeyOutput[34]), .Z(SubCellInst_LFInst_8_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_3_U6  ( .A1(
        SubCellInst_LFInst_8_LFInst_3_n13 ), .A2(
        SubCellInst_LFInst_8_LFInst_3_n12 ), .ZN(
        SubCellInst_LFInst_8_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_3_U5  ( .A1(AddRoundKeyOutput[32]), 
        .A2(AddRoundKeyOutput[34]), .ZN(SubCellInst_LFInst_8_LFInst_3_n12 )
         );
  XNOR2_X1 SubCellInst_LFInst_8_LFInst_3_U4  ( .A(AddRoundKeyOutput[32]), .B(
        SubCellInst_LFInst_8_LFInst_3_n11 ), .ZN(
        SubCellInst_LFInst_8_LFInst_3_n13 ) );
  OR2_X1 SubCellInst_LFInst_8_LFInst_3_U3  ( .A1(AddRoundKeyOutput[35]), .A2(
        AddRoundKeyOutput[33]), .ZN(SubCellInst_LFInst_8_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_2_U11  ( .A1(
        SubCellInst_LFInst_8_LFInst_2_n22 ), .A2(
        SubCellInst_LFInst_8_LFInst_2_n21 ), .ZN(MCInst1_MC2_v1_3 [3]) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_2_U10  ( .A1(AddRoundKeyOutput[34]), 
        .A2(SubCellInst_LFInst_8_LFInst_2_n20 ), .ZN(
        SubCellInst_LFInst_8_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst_LFInst_8_LFInst_2_U9  ( .A1(AddRoundKeyOutput[33]), 
        .A2(SubCellInst_LFInst_8_LFInst_2_n19 ), .ZN(
        SubCellInst_LFInst_8_LFInst_2_n20 ) );
  INV_X1 SubCellInst_LFInst_8_LFInst_2_U8  ( .A(AddRoundKeyOutput[35]), .ZN(
        SubCellInst_LFInst_8_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_2_U7  ( .A1(
        SubCellInst_LFInst_8_LFInst_2_n18 ), .A2(
        SubCellInst_LFInst_8_LFInst_2_n17 ), .ZN(
        SubCellInst_LFInst_8_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst_LFInst_8_LFInst_2_U6  ( .A(
        SubCellInst_LFInst_8_LFInst_2_n16 ), .B(AddRoundKeyOutput[34]), .Z(
        SubCellInst_LFInst_8_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_2_U5  ( .A1(AddRoundKeyOutput[32]), 
        .A2(AddRoundKeyOutput[33]), .ZN(SubCellInst_LFInst_8_LFInst_2_n16 )
         );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_2_U4  ( .A1(
        SubCellInst_LFInst_8_LFInst_2_n15 ), .A2(AddRoundKeyOutput[35]), .ZN(
        SubCellInst_LFInst_8_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst_LFInst_8_LFInst_2_U3  ( .A(AddRoundKeyOutput[32]), .B(
        AddRoundKeyOutput[33]), .ZN(SubCellInst_LFInst_8_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_1_U12  ( .A1(
        SubCellInst_LFInst_8_LFInst_1_n18 ), .A2(
        SubCellInst_LFInst_8_LFInst_1_n17 ), .ZN(MCInst1_MC2_v1_3 [2]) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_1_U11  ( .A1(AddRoundKeyOutput[33]), 
        .A2(SubCellInst_LFInst_8_LFInst_1_n16 ), .ZN(
        SubCellInst_LFInst_8_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst_LFInst_8_LFInst_1_U10  ( .A1(AddRoundKeyOutput[35]), 
        .A2(SubCellInst_LFInst_8_LFInst_1_n15 ), .ZN(
        SubCellInst_LFInst_8_LFInst_1_n16 ) );
  AND2_X1 SubCellInst_LFInst_8_LFInst_1_U9  ( .A1(AddRoundKeyOutput[32]), 
        .A2(AddRoundKeyOutput[34]), .ZN(SubCellInst_LFInst_8_LFInst_1_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_1_U8  ( .A1(AddRoundKeyOutput[35]), 
        .A2(SubCellInst_LFInst_8_LFInst_1_n14 ), .ZN(
        SubCellInst_LFInst_8_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_1_U7  ( .A1(
        SubCellInst_LFInst_8_LFInst_1_n13 ), .A2(
        SubCellInst_LFInst_8_LFInst_1_n12 ), .ZN(
        SubCellInst_LFInst_8_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_1_U6  ( .A1(AddRoundKeyOutput[32]), 
        .A2(AddRoundKeyOutput[34]), .ZN(SubCellInst_LFInst_8_LFInst_1_n12 )
         );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_1_U5  ( .A1(
        SubCellInst_LFInst_8_LFInst_1_n11 ), .A2(
        SubCellInst_LFInst_8_LFInst_1_n10 ), .ZN(
        SubCellInst_LFInst_8_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_1_U4  ( .A1(AddRoundKeyOutput[32]), 
        .A2(AddRoundKeyOutput[33]), .ZN(SubCellInst_LFInst_8_LFInst_1_n10 )
         );
  INV_X1 SubCellInst_LFInst_8_LFInst_1_U3  ( .A(AddRoundKeyOutput[34]), .ZN(
        SubCellInst_LFInst_8_LFInst_1_n11 ) );
  XNOR2_X1 SubCellInst_LFInst_8_LFInst_0_U6  ( .A(
        SubCellInst_LFInst_8_LFInst_0_n6 ), .B(
        SubCellInst_LFInst_8_LFInst_0_n5 ), .ZN(ShiftRowsOutput[36]) );
  NAND2_X1 SubCellInst_LFInst_8_LFInst_0_U5  ( .A1(AddRoundKeyOutput[34]), 
        .A2(SubCellInst_LFInst_8_LFInst_0_n4 ), .ZN(
        SubCellInst_LFInst_8_LFInst_0_n5 ) );
  INV_X1 SubCellInst_LFInst_8_LFInst_0_U4  ( .A(AddRoundKeyOutput[33]), .ZN(
        SubCellInst_LFInst_8_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst_LFInst_8_LFInst_0_U3  ( .A(AddRoundKeyOutput[32]), .B(
        AddRoundKeyOutput[35]), .Z(SubCellInst_LFInst_8_LFInst_0_n6 ) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_3_U9  ( .A1(
        SubCellInst_LFInst_9_LFInst_3_n16 ), .A2(
        SubCellInst_LFInst_9_LFInst_3_n15 ), .ZN(MCInst1_MC1_v1_3 [0]) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_3_U8  ( .A1(AddRoundKeyOutput[37]), 
        .A2(SubCellInst_LFInst_9_LFInst_3_n14 ), .ZN(
        SubCellInst_LFInst_9_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst_LFInst_9_LFInst_3_U7  ( .A(AddRoundKeyOutput[39]), .B(
        AddRoundKeyOutput[38]), .Z(SubCellInst_LFInst_9_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_3_U6  ( .A1(
        SubCellInst_LFInst_9_LFInst_3_n13 ), .A2(
        SubCellInst_LFInst_9_LFInst_3_n12 ), .ZN(
        SubCellInst_LFInst_9_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_3_U5  ( .A1(AddRoundKeyOutput[36]), 
        .A2(AddRoundKeyOutput[38]), .ZN(SubCellInst_LFInst_9_LFInst_3_n12 )
         );
  XNOR2_X1 SubCellInst_LFInst_9_LFInst_3_U4  ( .A(AddRoundKeyOutput[36]), .B(
        SubCellInst_LFInst_9_LFInst_3_n11 ), .ZN(
        SubCellInst_LFInst_9_LFInst_3_n13 ) );
  OR2_X1 SubCellInst_LFInst_9_LFInst_3_U3  ( .A1(AddRoundKeyOutput[39]), .A2(
        AddRoundKeyOutput[37]), .ZN(SubCellInst_LFInst_9_LFInst_3_n11 ) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_2_U11  ( .A1(
        SubCellInst_LFInst_9_LFInst_2_n22 ), .A2(
        SubCellInst_LFInst_9_LFInst_2_n21 ), .ZN(MCInst1_MC1_v1_3 [3]) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_2_U10  ( .A1(AddRoundKeyOutput[38]), 
        .A2(SubCellInst_LFInst_9_LFInst_2_n20 ), .ZN(
        SubCellInst_LFInst_9_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst_LFInst_9_LFInst_2_U9  ( .A1(AddRoundKeyOutput[37]), 
        .A2(SubCellInst_LFInst_9_LFInst_2_n19 ), .ZN(
        SubCellInst_LFInst_9_LFInst_2_n20 ) );
  INV_X1 SubCellInst_LFInst_9_LFInst_2_U8  ( .A(AddRoundKeyOutput[39]), .ZN(
        SubCellInst_LFInst_9_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_2_U7  ( .A1(
        SubCellInst_LFInst_9_LFInst_2_n18 ), .A2(
        SubCellInst_LFInst_9_LFInst_2_n17 ), .ZN(
        SubCellInst_LFInst_9_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst_LFInst_9_LFInst_2_U6  ( .A(
        SubCellInst_LFInst_9_LFInst_2_n16 ), .B(AddRoundKeyOutput[38]), .Z(
        SubCellInst_LFInst_9_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_2_U5  ( .A1(AddRoundKeyOutput[36]), 
        .A2(AddRoundKeyOutput[37]), .ZN(SubCellInst_LFInst_9_LFInst_2_n16 )
         );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_2_U4  ( .A1(
        SubCellInst_LFInst_9_LFInst_2_n15 ), .A2(AddRoundKeyOutput[39]), .ZN(
        SubCellInst_LFInst_9_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst_LFInst_9_LFInst_2_U3  ( .A(AddRoundKeyOutput[36]), .B(
        AddRoundKeyOutput[37]), .ZN(SubCellInst_LFInst_9_LFInst_2_n15 ) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_1_U12  ( .A1(
        SubCellInst_LFInst_9_LFInst_1_n18 ), .A2(
        SubCellInst_LFInst_9_LFInst_1_n17 ), .ZN(MCInst1_MC1_v1_3 [2]) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_1_U11  ( .A1(AddRoundKeyOutput[37]), 
        .A2(SubCellInst_LFInst_9_LFInst_1_n16 ), .ZN(
        SubCellInst_LFInst_9_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst_LFInst_9_LFInst_1_U10  ( .A1(AddRoundKeyOutput[39]), 
        .A2(SubCellInst_LFInst_9_LFInst_1_n15 ), .ZN(
        SubCellInst_LFInst_9_LFInst_1_n16 ) );
  AND2_X1 SubCellInst_LFInst_9_LFInst_1_U9  ( .A1(AddRoundKeyOutput[36]), 
        .A2(AddRoundKeyOutput[38]), .ZN(SubCellInst_LFInst_9_LFInst_1_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_1_U8  ( .A1(AddRoundKeyOutput[39]), 
        .A2(SubCellInst_LFInst_9_LFInst_1_n14 ), .ZN(
        SubCellInst_LFInst_9_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_1_U7  ( .A1(
        SubCellInst_LFInst_9_LFInst_1_n13 ), .A2(
        SubCellInst_LFInst_9_LFInst_1_n12 ), .ZN(
        SubCellInst_LFInst_9_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_1_U6  ( .A1(AddRoundKeyOutput[36]), 
        .A2(AddRoundKeyOutput[38]), .ZN(SubCellInst_LFInst_9_LFInst_1_n12 )
         );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_1_U5  ( .A1(
        SubCellInst_LFInst_9_LFInst_1_n11 ), .A2(
        SubCellInst_LFInst_9_LFInst_1_n10 ), .ZN(
        SubCellInst_LFInst_9_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_1_U4  ( .A1(AddRoundKeyOutput[36]), 
        .A2(AddRoundKeyOutput[37]), .ZN(SubCellInst_LFInst_9_LFInst_1_n10 )
         );
  INV_X1 SubCellInst_LFInst_9_LFInst_1_U3  ( .A(AddRoundKeyOutput[38]), .ZN(
        SubCellInst_LFInst_9_LFInst_1_n11 ) );
  XNOR2_X1 SubCellInst_LFInst_9_LFInst_0_U6  ( .A(
        SubCellInst_LFInst_9_LFInst_0_n6 ), .B(
        SubCellInst_LFInst_9_LFInst_0_n5 ), .ZN(ShiftRowsOutput[40]) );
  NAND2_X1 SubCellInst_LFInst_9_LFInst_0_U5  ( .A1(AddRoundKeyOutput[38]), 
        .A2(SubCellInst_LFInst_9_LFInst_0_n4 ), .ZN(
        SubCellInst_LFInst_9_LFInst_0_n5 ) );
  INV_X1 SubCellInst_LFInst_9_LFInst_0_U4  ( .A(AddRoundKeyOutput[37]), .ZN(
        SubCellInst_LFInst_9_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst_LFInst_9_LFInst_0_U3  ( .A(AddRoundKeyOutput[36]), .B(
        AddRoundKeyOutput[39]), .Z(SubCellInst_LFInst_9_LFInst_0_n6 ) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_3_U9  ( .A1(
        SubCellInst_LFInst_10_LFInst_3_n16 ), .A2(
        SubCellInst_LFInst_10_LFInst_3_n15 ), .ZN(MCInst1_MC0_v1_3 [0]) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_3_U8  ( .A1(AddRoundKeyOutput[41]), 
        .A2(SubCellInst_LFInst_10_LFInst_3_n14 ), .ZN(
        SubCellInst_LFInst_10_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst_LFInst_10_LFInst_3_U7  ( .A(AddRoundKeyOutput[43]), .B(
        AddRoundKeyOutput[42]), .Z(SubCellInst_LFInst_10_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_3_U6  ( .A1(
        SubCellInst_LFInst_10_LFInst_3_n13 ), .A2(
        SubCellInst_LFInst_10_LFInst_3_n12 ), .ZN(
        SubCellInst_LFInst_10_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_3_U5  ( .A1(AddRoundKeyOutput[40]), 
        .A2(AddRoundKeyOutput[42]), .ZN(SubCellInst_LFInst_10_LFInst_3_n12 )
         );
  XNOR2_X1 SubCellInst_LFInst_10_LFInst_3_U4  ( .A(AddRoundKeyOutput[40]), 
        .B(SubCellInst_LFInst_10_LFInst_3_n11 ), .ZN(
        SubCellInst_LFInst_10_LFInst_3_n13 ) );
  OR2_X1 SubCellInst_LFInst_10_LFInst_3_U3  ( .A1(AddRoundKeyOutput[43]), 
        .A2(AddRoundKeyOutput[41]), .ZN(SubCellInst_LFInst_10_LFInst_3_n11 )
         );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_2_U11  ( .A1(
        SubCellInst_LFInst_10_LFInst_2_n22 ), .A2(
        SubCellInst_LFInst_10_LFInst_2_n21 ), .ZN(MCInst1_MC0_v1_3 [3]) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_2_U10  ( .A1(AddRoundKeyOutput[42]), 
        .A2(SubCellInst_LFInst_10_LFInst_2_n20 ), .ZN(
        SubCellInst_LFInst_10_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst_LFInst_10_LFInst_2_U9  ( .A1(AddRoundKeyOutput[41]), 
        .A2(SubCellInst_LFInst_10_LFInst_2_n19 ), .ZN(
        SubCellInst_LFInst_10_LFInst_2_n20 ) );
  INV_X1 SubCellInst_LFInst_10_LFInst_2_U8  ( .A(AddRoundKeyOutput[43]), .ZN(
        SubCellInst_LFInst_10_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_2_U7  ( .A1(
        SubCellInst_LFInst_10_LFInst_2_n18 ), .A2(
        SubCellInst_LFInst_10_LFInst_2_n17 ), .ZN(
        SubCellInst_LFInst_10_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst_LFInst_10_LFInst_2_U6  ( .A(
        SubCellInst_LFInst_10_LFInst_2_n16 ), .B(AddRoundKeyOutput[42]), .Z(
        SubCellInst_LFInst_10_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_2_U5  ( .A1(AddRoundKeyOutput[40]), 
        .A2(AddRoundKeyOutput[41]), .ZN(SubCellInst_LFInst_10_LFInst_2_n16 )
         );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_2_U4  ( .A1(
        SubCellInst_LFInst_10_LFInst_2_n15 ), .A2(AddRoundKeyOutput[43]), 
        .ZN(SubCellInst_LFInst_10_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst_LFInst_10_LFInst_2_U3  ( .A(AddRoundKeyOutput[40]), 
        .B(AddRoundKeyOutput[41]), .ZN(SubCellInst_LFInst_10_LFInst_2_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_1_U12  ( .A1(
        SubCellInst_LFInst_10_LFInst_1_n18 ), .A2(
        SubCellInst_LFInst_10_LFInst_1_n17 ), .ZN(MCInst1_MC0_v1_3 [2]) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_1_U11  ( .A1(AddRoundKeyOutput[41]), 
        .A2(SubCellInst_LFInst_10_LFInst_1_n16 ), .ZN(
        SubCellInst_LFInst_10_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst_LFInst_10_LFInst_1_U10  ( .A1(AddRoundKeyOutput[43]), 
        .A2(SubCellInst_LFInst_10_LFInst_1_n15 ), .ZN(
        SubCellInst_LFInst_10_LFInst_1_n16 ) );
  AND2_X1 SubCellInst_LFInst_10_LFInst_1_U9  ( .A1(AddRoundKeyOutput[40]), 
        .A2(AddRoundKeyOutput[42]), .ZN(SubCellInst_LFInst_10_LFInst_1_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_1_U8  ( .A1(AddRoundKeyOutput[43]), 
        .A2(SubCellInst_LFInst_10_LFInst_1_n14 ), .ZN(
        SubCellInst_LFInst_10_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_1_U7  ( .A1(
        SubCellInst_LFInst_10_LFInst_1_n13 ), .A2(
        SubCellInst_LFInst_10_LFInst_1_n12 ), .ZN(
        SubCellInst_LFInst_10_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_1_U6  ( .A1(AddRoundKeyOutput[40]), 
        .A2(AddRoundKeyOutput[42]), .ZN(SubCellInst_LFInst_10_LFInst_1_n12 )
         );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_1_U5  ( .A1(
        SubCellInst_LFInst_10_LFInst_1_n11 ), .A2(
        SubCellInst_LFInst_10_LFInst_1_n10 ), .ZN(
        SubCellInst_LFInst_10_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_1_U4  ( .A1(AddRoundKeyOutput[40]), 
        .A2(AddRoundKeyOutput[41]), .ZN(SubCellInst_LFInst_10_LFInst_1_n10 )
         );
  INV_X1 SubCellInst_LFInst_10_LFInst_1_U3  ( .A(AddRoundKeyOutput[42]), .ZN(
        SubCellInst_LFInst_10_LFInst_1_n11 ) );
  XNOR2_X1 SubCellInst_LFInst_10_LFInst_0_U6  ( .A(
        SubCellInst_LFInst_10_LFInst_0_n6 ), .B(
        SubCellInst_LFInst_10_LFInst_0_n5 ), .ZN(ShiftRowsOutput[44]) );
  NAND2_X1 SubCellInst_LFInst_10_LFInst_0_U5  ( .A1(AddRoundKeyOutput[42]), 
        .A2(SubCellInst_LFInst_10_LFInst_0_n4 ), .ZN(
        SubCellInst_LFInst_10_LFInst_0_n5 ) );
  INV_X1 SubCellInst_LFInst_10_LFInst_0_U4  ( .A(AddRoundKeyOutput[41]), .ZN(
        SubCellInst_LFInst_10_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst_LFInst_10_LFInst_0_U3  ( .A(AddRoundKeyOutput[40]), .B(
        AddRoundKeyOutput[43]), .Z(SubCellInst_LFInst_10_LFInst_0_n6 ) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_3_U9  ( .A1(
        SubCellInst_LFInst_11_LFInst_3_n16 ), .A2(
        SubCellInst_LFInst_11_LFInst_3_n15 ), .ZN(MCInst1_MC3_v1_3 [0]) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_3_U8  ( .A1(AddRoundKeyOutput[45]), 
        .A2(SubCellInst_LFInst_11_LFInst_3_n14 ), .ZN(
        SubCellInst_LFInst_11_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst_LFInst_11_LFInst_3_U7  ( .A(AddRoundKeyOutput[47]), .B(
        AddRoundKeyOutput[46]), .Z(SubCellInst_LFInst_11_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_3_U6  ( .A1(
        SubCellInst_LFInst_11_LFInst_3_n13 ), .A2(
        SubCellInst_LFInst_11_LFInst_3_n12 ), .ZN(
        SubCellInst_LFInst_11_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_3_U5  ( .A1(AddRoundKeyOutput[44]), 
        .A2(AddRoundKeyOutput[46]), .ZN(SubCellInst_LFInst_11_LFInst_3_n12 )
         );
  XNOR2_X1 SubCellInst_LFInst_11_LFInst_3_U4  ( .A(AddRoundKeyOutput[44]), 
        .B(SubCellInst_LFInst_11_LFInst_3_n11 ), .ZN(
        SubCellInst_LFInst_11_LFInst_3_n13 ) );
  OR2_X1 SubCellInst_LFInst_11_LFInst_3_U3  ( .A1(AddRoundKeyOutput[47]), 
        .A2(AddRoundKeyOutput[45]), .ZN(SubCellInst_LFInst_11_LFInst_3_n11 )
         );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_2_U11  ( .A1(
        SubCellInst_LFInst_11_LFInst_2_n22 ), .A2(
        SubCellInst_LFInst_11_LFInst_2_n21 ), .ZN(MCInst1_MC3_v1_3 [3]) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_2_U10  ( .A1(AddRoundKeyOutput[46]), 
        .A2(SubCellInst_LFInst_11_LFInst_2_n20 ), .ZN(
        SubCellInst_LFInst_11_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst_LFInst_11_LFInst_2_U9  ( .A1(AddRoundKeyOutput[45]), 
        .A2(SubCellInst_LFInst_11_LFInst_2_n19 ), .ZN(
        SubCellInst_LFInst_11_LFInst_2_n20 ) );
  INV_X1 SubCellInst_LFInst_11_LFInst_2_U8  ( .A(AddRoundKeyOutput[47]), .ZN(
        SubCellInst_LFInst_11_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_2_U7  ( .A1(
        SubCellInst_LFInst_11_LFInst_2_n18 ), .A2(
        SubCellInst_LFInst_11_LFInst_2_n17 ), .ZN(
        SubCellInst_LFInst_11_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst_LFInst_11_LFInst_2_U6  ( .A(
        SubCellInst_LFInst_11_LFInst_2_n16 ), .B(AddRoundKeyOutput[46]), .Z(
        SubCellInst_LFInst_11_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_2_U5  ( .A1(AddRoundKeyOutput[44]), 
        .A2(AddRoundKeyOutput[45]), .ZN(SubCellInst_LFInst_11_LFInst_2_n16 )
         );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_2_U4  ( .A1(
        SubCellInst_LFInst_11_LFInst_2_n15 ), .A2(AddRoundKeyOutput[47]), 
        .ZN(SubCellInst_LFInst_11_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst_LFInst_11_LFInst_2_U3  ( .A(AddRoundKeyOutput[44]), 
        .B(AddRoundKeyOutput[45]), .ZN(SubCellInst_LFInst_11_LFInst_2_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_1_U12  ( .A1(
        SubCellInst_LFInst_11_LFInst_1_n18 ), .A2(
        SubCellInst_LFInst_11_LFInst_1_n17 ), .ZN(MCInst1_MC3_v1_3 [2]) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_1_U11  ( .A1(AddRoundKeyOutput[45]), 
        .A2(SubCellInst_LFInst_11_LFInst_1_n16 ), .ZN(
        SubCellInst_LFInst_11_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst_LFInst_11_LFInst_1_U10  ( .A1(AddRoundKeyOutput[47]), 
        .A2(SubCellInst_LFInst_11_LFInst_1_n15 ), .ZN(
        SubCellInst_LFInst_11_LFInst_1_n16 ) );
  AND2_X1 SubCellInst_LFInst_11_LFInst_1_U9  ( .A1(AddRoundKeyOutput[44]), 
        .A2(AddRoundKeyOutput[46]), .ZN(SubCellInst_LFInst_11_LFInst_1_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_1_U8  ( .A1(AddRoundKeyOutput[47]), 
        .A2(SubCellInst_LFInst_11_LFInst_1_n14 ), .ZN(
        SubCellInst_LFInst_11_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_1_U7  ( .A1(
        SubCellInst_LFInst_11_LFInst_1_n13 ), .A2(
        SubCellInst_LFInst_11_LFInst_1_n12 ), .ZN(
        SubCellInst_LFInst_11_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_1_U6  ( .A1(AddRoundKeyOutput[44]), 
        .A2(AddRoundKeyOutput[46]), .ZN(SubCellInst_LFInst_11_LFInst_1_n12 )
         );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_1_U5  ( .A1(
        SubCellInst_LFInst_11_LFInst_1_n11 ), .A2(
        SubCellInst_LFInst_11_LFInst_1_n10 ), .ZN(
        SubCellInst_LFInst_11_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_1_U4  ( .A1(AddRoundKeyOutput[44]), 
        .A2(AddRoundKeyOutput[45]), .ZN(SubCellInst_LFInst_11_LFInst_1_n10 )
         );
  INV_X1 SubCellInst_LFInst_11_LFInst_1_U3  ( .A(AddRoundKeyOutput[46]), .ZN(
        SubCellInst_LFInst_11_LFInst_1_n11 ) );
  XNOR2_X1 SubCellInst_LFInst_11_LFInst_0_U6  ( .A(
        SubCellInst_LFInst_11_LFInst_0_n6 ), .B(
        SubCellInst_LFInst_11_LFInst_0_n5 ), .ZN(ShiftRowsOutput[32]) );
  NAND2_X1 SubCellInst_LFInst_11_LFInst_0_U5  ( .A1(AddRoundKeyOutput[46]), 
        .A2(SubCellInst_LFInst_11_LFInst_0_n4 ), .ZN(
        SubCellInst_LFInst_11_LFInst_0_n5 ) );
  INV_X1 SubCellInst_LFInst_11_LFInst_0_U4  ( .A(AddRoundKeyOutput[45]), .ZN(
        SubCellInst_LFInst_11_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst_LFInst_11_LFInst_0_U3  ( .A(AddRoundKeyOutput[44]), .B(
        AddRoundKeyOutput[47]), .Z(SubCellInst_LFInst_11_LFInst_0_n6 ) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_3_U9  ( .A1(
        SubCellInst_LFInst_12_LFInst_3_n16 ), .A2(
        SubCellInst_LFInst_12_LFInst_3_n15 ), .ZN(MCInst1_MC3_v0_3 [0]) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_3_U8  ( .A1(AddRoundKeyOutput[49]), 
        .A2(SubCellInst_LFInst_12_LFInst_3_n14 ), .ZN(
        SubCellInst_LFInst_12_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst_LFInst_12_LFInst_3_U7  ( .A(AddRoundKeyOutput[51]), .B(
        AddRoundKeyOutput[50]), .Z(SubCellInst_LFInst_12_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_3_U6  ( .A1(
        SubCellInst_LFInst_12_LFInst_3_n13 ), .A2(
        SubCellInst_LFInst_12_LFInst_3_n12 ), .ZN(
        SubCellInst_LFInst_12_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_3_U5  ( .A1(AddRoundKeyOutput[48]), 
        .A2(AddRoundKeyOutput[50]), .ZN(SubCellInst_LFInst_12_LFInst_3_n12 )
         );
  XNOR2_X1 SubCellInst_LFInst_12_LFInst_3_U4  ( .A(AddRoundKeyOutput[48]), 
        .B(SubCellInst_LFInst_12_LFInst_3_n11 ), .ZN(
        SubCellInst_LFInst_12_LFInst_3_n13 ) );
  OR2_X1 SubCellInst_LFInst_12_LFInst_3_U3  ( .A1(AddRoundKeyOutput[51]), 
        .A2(AddRoundKeyOutput[49]), .ZN(SubCellInst_LFInst_12_LFInst_3_n11 )
         );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_2_U11  ( .A1(
        SubCellInst_LFInst_12_LFInst_2_n22 ), .A2(
        SubCellInst_LFInst_12_LFInst_2_n21 ), .ZN(MCInst1_MC3_v0_3 [3]) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_2_U10  ( .A1(AddRoundKeyOutput[50]), 
        .A2(SubCellInst_LFInst_12_LFInst_2_n20 ), .ZN(
        SubCellInst_LFInst_12_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst_LFInst_12_LFInst_2_U9  ( .A1(AddRoundKeyOutput[49]), 
        .A2(SubCellInst_LFInst_12_LFInst_2_n19 ), .ZN(
        SubCellInst_LFInst_12_LFInst_2_n20 ) );
  INV_X1 SubCellInst_LFInst_12_LFInst_2_U8  ( .A(AddRoundKeyOutput[51]), .ZN(
        SubCellInst_LFInst_12_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_2_U7  ( .A1(
        SubCellInst_LFInst_12_LFInst_2_n18 ), .A2(
        SubCellInst_LFInst_12_LFInst_2_n17 ), .ZN(
        SubCellInst_LFInst_12_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst_LFInst_12_LFInst_2_U6  ( .A(
        SubCellInst_LFInst_12_LFInst_2_n16 ), .B(AddRoundKeyOutput[50]), .Z(
        SubCellInst_LFInst_12_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_2_U5  ( .A1(AddRoundKeyOutput[48]), 
        .A2(AddRoundKeyOutput[49]), .ZN(SubCellInst_LFInst_12_LFInst_2_n16 )
         );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_2_U4  ( .A1(
        SubCellInst_LFInst_12_LFInst_2_n15 ), .A2(AddRoundKeyOutput[51]), 
        .ZN(SubCellInst_LFInst_12_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst_LFInst_12_LFInst_2_U3  ( .A(AddRoundKeyOutput[48]), 
        .B(AddRoundKeyOutput[49]), .ZN(SubCellInst_LFInst_12_LFInst_2_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_1_U12  ( .A1(
        SubCellInst_LFInst_12_LFInst_1_n18 ), .A2(
        SubCellInst_LFInst_12_LFInst_1_n17 ), .ZN(MCInst1_MC3_v0_0 [3]) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_1_U11  ( .A1(AddRoundKeyOutput[49]), 
        .A2(SubCellInst_LFInst_12_LFInst_1_n16 ), .ZN(
        SubCellInst_LFInst_12_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst_LFInst_12_LFInst_1_U10  ( .A1(AddRoundKeyOutput[51]), 
        .A2(SubCellInst_LFInst_12_LFInst_1_n15 ), .ZN(
        SubCellInst_LFInst_12_LFInst_1_n16 ) );
  AND2_X1 SubCellInst_LFInst_12_LFInst_1_U9  ( .A1(AddRoundKeyOutput[48]), 
        .A2(AddRoundKeyOutput[50]), .ZN(SubCellInst_LFInst_12_LFInst_1_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_1_U8  ( .A1(AddRoundKeyOutput[51]), 
        .A2(SubCellInst_LFInst_12_LFInst_1_n14 ), .ZN(
        SubCellInst_LFInst_12_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_1_U7  ( .A1(
        SubCellInst_LFInst_12_LFInst_1_n13 ), .A2(
        SubCellInst_LFInst_12_LFInst_1_n12 ), .ZN(
        SubCellInst_LFInst_12_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_1_U6  ( .A1(AddRoundKeyOutput[48]), 
        .A2(AddRoundKeyOutput[50]), .ZN(SubCellInst_LFInst_12_LFInst_1_n12 )
         );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_1_U5  ( .A1(
        SubCellInst_LFInst_12_LFInst_1_n11 ), .A2(
        SubCellInst_LFInst_12_LFInst_1_n10 ), .ZN(
        SubCellInst_LFInst_12_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_1_U4  ( .A1(AddRoundKeyOutput[48]), 
        .A2(AddRoundKeyOutput[49]), .ZN(SubCellInst_LFInst_12_LFInst_1_n10 )
         );
  INV_X1 SubCellInst_LFInst_12_LFInst_1_U3  ( .A(AddRoundKeyOutput[50]), .ZN(
        SubCellInst_LFInst_12_LFInst_1_n11 ) );
  XNOR2_X1 SubCellInst_LFInst_12_LFInst_0_U6  ( .A(
        SubCellInst_LFInst_12_LFInst_0_n6 ), .B(
        SubCellInst_LFInst_12_LFInst_0_n5 ), .ZN(ShiftRowsOutput[48]) );
  NAND2_X1 SubCellInst_LFInst_12_LFInst_0_U5  ( .A1(AddRoundKeyOutput[50]), 
        .A2(SubCellInst_LFInst_12_LFInst_0_n4 ), .ZN(
        SubCellInst_LFInst_12_LFInst_0_n5 ) );
  INV_X1 SubCellInst_LFInst_12_LFInst_0_U4  ( .A(AddRoundKeyOutput[49]), .ZN(
        SubCellInst_LFInst_12_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst_LFInst_12_LFInst_0_U3  ( .A(AddRoundKeyOutput[48]), .B(
        AddRoundKeyOutput[51]), .Z(SubCellInst_LFInst_12_LFInst_0_n6 ) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_3_U9  ( .A1(
        SubCellInst_LFInst_13_LFInst_3_n16 ), .A2(
        SubCellInst_LFInst_13_LFInst_3_n15 ), .ZN(MCInst1_MC2_v0_3 [0]) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_3_U8  ( .A1(AddRoundKeyOutput[53]), 
        .A2(SubCellInst_LFInst_13_LFInst_3_n14 ), .ZN(
        SubCellInst_LFInst_13_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst_LFInst_13_LFInst_3_U7  ( .A(AddRoundKeyOutput[55]), .B(
        AddRoundKeyOutput[54]), .Z(SubCellInst_LFInst_13_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_3_U6  ( .A1(
        SubCellInst_LFInst_13_LFInst_3_n13 ), .A2(
        SubCellInst_LFInst_13_LFInst_3_n12 ), .ZN(
        SubCellInst_LFInst_13_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_3_U5  ( .A1(AddRoundKeyOutput[52]), 
        .A2(AddRoundKeyOutput[54]), .ZN(SubCellInst_LFInst_13_LFInst_3_n12 )
         );
  XNOR2_X1 SubCellInst_LFInst_13_LFInst_3_U4  ( .A(AddRoundKeyOutput[52]), 
        .B(SubCellInst_LFInst_13_LFInst_3_n11 ), .ZN(
        SubCellInst_LFInst_13_LFInst_3_n13 ) );
  OR2_X1 SubCellInst_LFInst_13_LFInst_3_U3  ( .A1(AddRoundKeyOutput[55]), 
        .A2(AddRoundKeyOutput[53]), .ZN(SubCellInst_LFInst_13_LFInst_3_n11 )
         );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_2_U11  ( .A1(
        SubCellInst_LFInst_13_LFInst_2_n22 ), .A2(
        SubCellInst_LFInst_13_LFInst_2_n21 ), .ZN(MCInst1_MC2_v0_3 [3]) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_2_U10  ( .A1(AddRoundKeyOutput[54]), 
        .A2(SubCellInst_LFInst_13_LFInst_2_n20 ), .ZN(
        SubCellInst_LFInst_13_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst_LFInst_13_LFInst_2_U9  ( .A1(AddRoundKeyOutput[53]), 
        .A2(SubCellInst_LFInst_13_LFInst_2_n19 ), .ZN(
        SubCellInst_LFInst_13_LFInst_2_n20 ) );
  INV_X1 SubCellInst_LFInst_13_LFInst_2_U8  ( .A(AddRoundKeyOutput[55]), .ZN(
        SubCellInst_LFInst_13_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_2_U7  ( .A1(
        SubCellInst_LFInst_13_LFInst_2_n18 ), .A2(
        SubCellInst_LFInst_13_LFInst_2_n17 ), .ZN(
        SubCellInst_LFInst_13_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst_LFInst_13_LFInst_2_U6  ( .A(
        SubCellInst_LFInst_13_LFInst_2_n16 ), .B(AddRoundKeyOutput[54]), .Z(
        SubCellInst_LFInst_13_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_2_U5  ( .A1(AddRoundKeyOutput[52]), 
        .A2(AddRoundKeyOutput[53]), .ZN(SubCellInst_LFInst_13_LFInst_2_n16 )
         );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_2_U4  ( .A1(
        SubCellInst_LFInst_13_LFInst_2_n15 ), .A2(AddRoundKeyOutput[55]), 
        .ZN(SubCellInst_LFInst_13_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst_LFInst_13_LFInst_2_U3  ( .A(AddRoundKeyOutput[52]), 
        .B(AddRoundKeyOutput[53]), .ZN(SubCellInst_LFInst_13_LFInst_2_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_1_U12  ( .A1(
        SubCellInst_LFInst_13_LFInst_1_n18 ), .A2(
        SubCellInst_LFInst_13_LFInst_1_n17 ), .ZN(MCInst1_MC2_v0_0 [3]) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_1_U11  ( .A1(AddRoundKeyOutput[53]), 
        .A2(SubCellInst_LFInst_13_LFInst_1_n16 ), .ZN(
        SubCellInst_LFInst_13_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst_LFInst_13_LFInst_1_U10  ( .A1(AddRoundKeyOutput[55]), 
        .A2(SubCellInst_LFInst_13_LFInst_1_n15 ), .ZN(
        SubCellInst_LFInst_13_LFInst_1_n16 ) );
  AND2_X1 SubCellInst_LFInst_13_LFInst_1_U9  ( .A1(AddRoundKeyOutput[52]), 
        .A2(AddRoundKeyOutput[54]), .ZN(SubCellInst_LFInst_13_LFInst_1_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_1_U8  ( .A1(AddRoundKeyOutput[55]), 
        .A2(SubCellInst_LFInst_13_LFInst_1_n14 ), .ZN(
        SubCellInst_LFInst_13_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_1_U7  ( .A1(
        SubCellInst_LFInst_13_LFInst_1_n13 ), .A2(
        SubCellInst_LFInst_13_LFInst_1_n12 ), .ZN(
        SubCellInst_LFInst_13_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_1_U6  ( .A1(AddRoundKeyOutput[52]), 
        .A2(AddRoundKeyOutput[54]), .ZN(SubCellInst_LFInst_13_LFInst_1_n12 )
         );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_1_U5  ( .A1(
        SubCellInst_LFInst_13_LFInst_1_n11 ), .A2(
        SubCellInst_LFInst_13_LFInst_1_n10 ), .ZN(
        SubCellInst_LFInst_13_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_1_U4  ( .A1(AddRoundKeyOutput[52]), 
        .A2(AddRoundKeyOutput[53]), .ZN(SubCellInst_LFInst_13_LFInst_1_n10 )
         );
  INV_X1 SubCellInst_LFInst_13_LFInst_1_U3  ( .A(AddRoundKeyOutput[54]), .ZN(
        SubCellInst_LFInst_13_LFInst_1_n11 ) );
  XNOR2_X1 SubCellInst_LFInst_13_LFInst_0_U6  ( .A(
        SubCellInst_LFInst_13_LFInst_0_n6 ), .B(
        SubCellInst_LFInst_13_LFInst_0_n5 ), .ZN(ShiftRowsOutput[52]) );
  NAND2_X1 SubCellInst_LFInst_13_LFInst_0_U5  ( .A1(AddRoundKeyOutput[54]), 
        .A2(SubCellInst_LFInst_13_LFInst_0_n4 ), .ZN(
        SubCellInst_LFInst_13_LFInst_0_n5 ) );
  INV_X1 SubCellInst_LFInst_13_LFInst_0_U4  ( .A(AddRoundKeyOutput[53]), .ZN(
        SubCellInst_LFInst_13_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst_LFInst_13_LFInst_0_U3  ( .A(AddRoundKeyOutput[52]), .B(
        AddRoundKeyOutput[55]), .Z(SubCellInst_LFInst_13_LFInst_0_n6 ) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_3_U9  ( .A1(
        SubCellInst_LFInst_14_LFInst_3_n16 ), .A2(
        SubCellInst_LFInst_14_LFInst_3_n15 ), .ZN(MCInst1_MC1_v0_3 [0]) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_3_U8  ( .A1(AddRoundKeyOutput[57]), 
        .A2(SubCellInst_LFInst_14_LFInst_3_n14 ), .ZN(
        SubCellInst_LFInst_14_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst_LFInst_14_LFInst_3_U7  ( .A(AddRoundKeyOutput[59]), .B(
        AddRoundKeyOutput[58]), .Z(SubCellInst_LFInst_14_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_3_U6  ( .A1(
        SubCellInst_LFInst_14_LFInst_3_n13 ), .A2(
        SubCellInst_LFInst_14_LFInst_3_n12 ), .ZN(
        SubCellInst_LFInst_14_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_3_U5  ( .A1(AddRoundKeyOutput[56]), 
        .A2(AddRoundKeyOutput[58]), .ZN(SubCellInst_LFInst_14_LFInst_3_n12 )
         );
  XNOR2_X1 SubCellInst_LFInst_14_LFInst_3_U4  ( .A(AddRoundKeyOutput[56]), 
        .B(SubCellInst_LFInst_14_LFInst_3_n11 ), .ZN(
        SubCellInst_LFInst_14_LFInst_3_n13 ) );
  OR2_X1 SubCellInst_LFInst_14_LFInst_3_U3  ( .A1(AddRoundKeyOutput[59]), 
        .A2(AddRoundKeyOutput[57]), .ZN(SubCellInst_LFInst_14_LFInst_3_n11 )
         );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_2_U11  ( .A1(
        SubCellInst_LFInst_14_LFInst_2_n22 ), .A2(
        SubCellInst_LFInst_14_LFInst_2_n21 ), .ZN(MCInst1_MC1_v0_3 [3]) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_2_U10  ( .A1(AddRoundKeyOutput[58]), 
        .A2(SubCellInst_LFInst_14_LFInst_2_n20 ), .ZN(
        SubCellInst_LFInst_14_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst_LFInst_14_LFInst_2_U9  ( .A1(AddRoundKeyOutput[57]), 
        .A2(SubCellInst_LFInst_14_LFInst_2_n19 ), .ZN(
        SubCellInst_LFInst_14_LFInst_2_n20 ) );
  INV_X1 SubCellInst_LFInst_14_LFInst_2_U8  ( .A(AddRoundKeyOutput[59]), .ZN(
        SubCellInst_LFInst_14_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_2_U7  ( .A1(
        SubCellInst_LFInst_14_LFInst_2_n18 ), .A2(
        SubCellInst_LFInst_14_LFInst_2_n17 ), .ZN(
        SubCellInst_LFInst_14_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst_LFInst_14_LFInst_2_U6  ( .A(
        SubCellInst_LFInst_14_LFInst_2_n16 ), .B(AddRoundKeyOutput[58]), .Z(
        SubCellInst_LFInst_14_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_2_U5  ( .A1(AddRoundKeyOutput[56]), 
        .A2(AddRoundKeyOutput[57]), .ZN(SubCellInst_LFInst_14_LFInst_2_n16 )
         );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_2_U4  ( .A1(
        SubCellInst_LFInst_14_LFInst_2_n15 ), .A2(AddRoundKeyOutput[59]), 
        .ZN(SubCellInst_LFInst_14_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst_LFInst_14_LFInst_2_U3  ( .A(AddRoundKeyOutput[56]), 
        .B(AddRoundKeyOutput[57]), .ZN(SubCellInst_LFInst_14_LFInst_2_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_1_U12  ( .A1(
        SubCellInst_LFInst_14_LFInst_1_n18 ), .A2(
        SubCellInst_LFInst_14_LFInst_1_n17 ), .ZN(MCInst1_MC1_v0_0 [3]) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_1_U11  ( .A1(AddRoundKeyOutput[57]), 
        .A2(SubCellInst_LFInst_14_LFInst_1_n16 ), .ZN(
        SubCellInst_LFInst_14_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst_LFInst_14_LFInst_1_U10  ( .A1(AddRoundKeyOutput[59]), 
        .A2(SubCellInst_LFInst_14_LFInst_1_n15 ), .ZN(
        SubCellInst_LFInst_14_LFInst_1_n16 ) );
  AND2_X1 SubCellInst_LFInst_14_LFInst_1_U9  ( .A1(AddRoundKeyOutput[56]), 
        .A2(AddRoundKeyOutput[58]), .ZN(SubCellInst_LFInst_14_LFInst_1_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_1_U8  ( .A1(AddRoundKeyOutput[59]), 
        .A2(SubCellInst_LFInst_14_LFInst_1_n14 ), .ZN(
        SubCellInst_LFInst_14_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_1_U7  ( .A1(
        SubCellInst_LFInst_14_LFInst_1_n13 ), .A2(
        SubCellInst_LFInst_14_LFInst_1_n12 ), .ZN(
        SubCellInst_LFInst_14_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_1_U6  ( .A1(AddRoundKeyOutput[56]), 
        .A2(AddRoundKeyOutput[58]), .ZN(SubCellInst_LFInst_14_LFInst_1_n12 )
         );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_1_U5  ( .A1(
        SubCellInst_LFInst_14_LFInst_1_n11 ), .A2(
        SubCellInst_LFInst_14_LFInst_1_n10 ), .ZN(
        SubCellInst_LFInst_14_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_1_U4  ( .A1(AddRoundKeyOutput[56]), 
        .A2(AddRoundKeyOutput[57]), .ZN(SubCellInst_LFInst_14_LFInst_1_n10 )
         );
  INV_X1 SubCellInst_LFInst_14_LFInst_1_U3  ( .A(AddRoundKeyOutput[58]), .ZN(
        SubCellInst_LFInst_14_LFInst_1_n11 ) );
  XNOR2_X1 SubCellInst_LFInst_14_LFInst_0_U6  ( .A(
        SubCellInst_LFInst_14_LFInst_0_n6 ), .B(
        SubCellInst_LFInst_14_LFInst_0_n5 ), .ZN(ShiftRowsOutput[56]) );
  NAND2_X1 SubCellInst_LFInst_14_LFInst_0_U5  ( .A1(AddRoundKeyOutput[58]), 
        .A2(SubCellInst_LFInst_14_LFInst_0_n4 ), .ZN(
        SubCellInst_LFInst_14_LFInst_0_n5 ) );
  INV_X1 SubCellInst_LFInst_14_LFInst_0_U4  ( .A(AddRoundKeyOutput[57]), .ZN(
        SubCellInst_LFInst_14_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst_LFInst_14_LFInst_0_U3  ( .A(AddRoundKeyOutput[56]), .B(
        AddRoundKeyOutput[59]), .Z(SubCellInst_LFInst_14_LFInst_0_n6 ) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_3_U9  ( .A1(
        SubCellInst_LFInst_15_LFInst_3_n16 ), .A2(
        SubCellInst_LFInst_15_LFInst_3_n15 ), .ZN(MCInst1_MC0_v0_3 [0]) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_3_U8  ( .A1(AddRoundKeyOutput[61]), 
        .A2(SubCellInst_LFInst_15_LFInst_3_n14 ), .ZN(
        SubCellInst_LFInst_15_LFInst_3_n15 ) );
  XOR2_X1 SubCellInst_LFInst_15_LFInst_3_U7  ( .A(AddRoundKeyOutput[63]), .B(
        AddRoundKeyOutput[62]), .Z(SubCellInst_LFInst_15_LFInst_3_n14 ) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_3_U6  ( .A1(
        SubCellInst_LFInst_15_LFInst_3_n13 ), .A2(
        SubCellInst_LFInst_15_LFInst_3_n12 ), .ZN(
        SubCellInst_LFInst_15_LFInst_3_n16 ) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_3_U5  ( .A1(AddRoundKeyOutput[60]), 
        .A2(AddRoundKeyOutput[62]), .ZN(SubCellInst_LFInst_15_LFInst_3_n12 )
         );
  XNOR2_X1 SubCellInst_LFInst_15_LFInst_3_U4  ( .A(AddRoundKeyOutput[60]), 
        .B(SubCellInst_LFInst_15_LFInst_3_n11 ), .ZN(
        SubCellInst_LFInst_15_LFInst_3_n13 ) );
  OR2_X1 SubCellInst_LFInst_15_LFInst_3_U3  ( .A1(AddRoundKeyOutput[63]), 
        .A2(AddRoundKeyOutput[61]), .ZN(SubCellInst_LFInst_15_LFInst_3_n11 )
         );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_2_U11  ( .A1(
        SubCellInst_LFInst_15_LFInst_2_n22 ), .A2(
        SubCellInst_LFInst_15_LFInst_2_n21 ), .ZN(MCInst1_MC0_v0_3 [3]) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_2_U10  ( .A1(AddRoundKeyOutput[62]), 
        .A2(SubCellInst_LFInst_15_LFInst_2_n20 ), .ZN(
        SubCellInst_LFInst_15_LFInst_2_n21 ) );
  NOR2_X1 SubCellInst_LFInst_15_LFInst_2_U9  ( .A1(AddRoundKeyOutput[61]), 
        .A2(SubCellInst_LFInst_15_LFInst_2_n19 ), .ZN(
        SubCellInst_LFInst_15_LFInst_2_n20 ) );
  INV_X1 SubCellInst_LFInst_15_LFInst_2_U8  ( .A(AddRoundKeyOutput[63]), .ZN(
        SubCellInst_LFInst_15_LFInst_2_n19 ) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_2_U7  ( .A1(
        SubCellInst_LFInst_15_LFInst_2_n18 ), .A2(
        SubCellInst_LFInst_15_LFInst_2_n17 ), .ZN(
        SubCellInst_LFInst_15_LFInst_2_n22 ) );
  XOR2_X1 SubCellInst_LFInst_15_LFInst_2_U6  ( .A(
        SubCellInst_LFInst_15_LFInst_2_n16 ), .B(AddRoundKeyOutput[62]), .Z(
        SubCellInst_LFInst_15_LFInst_2_n17 ) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_2_U5  ( .A1(AddRoundKeyOutput[60]), 
        .A2(AddRoundKeyOutput[61]), .ZN(SubCellInst_LFInst_15_LFInst_2_n16 )
         );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_2_U4  ( .A1(
        SubCellInst_LFInst_15_LFInst_2_n15 ), .A2(AddRoundKeyOutput[63]), 
        .ZN(SubCellInst_LFInst_15_LFInst_2_n18 ) );
  XNOR2_X1 SubCellInst_LFInst_15_LFInst_2_U3  ( .A(AddRoundKeyOutput[60]), 
        .B(AddRoundKeyOutput[61]), .ZN(SubCellInst_LFInst_15_LFInst_2_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_1_U12  ( .A1(
        SubCellInst_LFInst_15_LFInst_1_n18 ), .A2(
        SubCellInst_LFInst_15_LFInst_1_n17 ), .ZN(MCInst1_MC0_v0_0 [3]) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_1_U11  ( .A1(AddRoundKeyOutput[61]), 
        .A2(SubCellInst_LFInst_15_LFInst_1_n16 ), .ZN(
        SubCellInst_LFInst_15_LFInst_1_n17 ) );
  NOR2_X1 SubCellInst_LFInst_15_LFInst_1_U10  ( .A1(AddRoundKeyOutput[63]), 
        .A2(SubCellInst_LFInst_15_LFInst_1_n15 ), .ZN(
        SubCellInst_LFInst_15_LFInst_1_n16 ) );
  AND2_X1 SubCellInst_LFInst_15_LFInst_1_U9  ( .A1(AddRoundKeyOutput[60]), 
        .A2(AddRoundKeyOutput[62]), .ZN(SubCellInst_LFInst_15_LFInst_1_n15 )
         );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_1_U8  ( .A1(AddRoundKeyOutput[63]), 
        .A2(SubCellInst_LFInst_15_LFInst_1_n14 ), .ZN(
        SubCellInst_LFInst_15_LFInst_1_n18 ) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_1_U7  ( .A1(
        SubCellInst_LFInst_15_LFInst_1_n13 ), .A2(
        SubCellInst_LFInst_15_LFInst_1_n12 ), .ZN(
        SubCellInst_LFInst_15_LFInst_1_n14 ) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_1_U6  ( .A1(AddRoundKeyOutput[60]), 
        .A2(AddRoundKeyOutput[62]), .ZN(SubCellInst_LFInst_15_LFInst_1_n12 )
         );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_1_U5  ( .A1(
        SubCellInst_LFInst_15_LFInst_1_n11 ), .A2(
        SubCellInst_LFInst_15_LFInst_1_n10 ), .ZN(
        SubCellInst_LFInst_15_LFInst_1_n13 ) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_1_U4  ( .A1(AddRoundKeyOutput[60]), 
        .A2(AddRoundKeyOutput[61]), .ZN(SubCellInst_LFInst_15_LFInst_1_n10 )
         );
  INV_X1 SubCellInst_LFInst_15_LFInst_1_U3  ( .A(AddRoundKeyOutput[62]), .ZN(
        SubCellInst_LFInst_15_LFInst_1_n11 ) );
  XNOR2_X1 SubCellInst_LFInst_15_LFInst_0_U6  ( .A(
        SubCellInst_LFInst_15_LFInst_0_n6 ), .B(
        SubCellInst_LFInst_15_LFInst_0_n5 ), .ZN(ShiftRowsOutput[60]) );
  NAND2_X1 SubCellInst_LFInst_15_LFInst_0_U5  ( .A1(AddRoundKeyOutput[62]), 
        .A2(SubCellInst_LFInst_15_LFInst_0_n4 ), .ZN(
        SubCellInst_LFInst_15_LFInst_0_n5 ) );
  INV_X1 SubCellInst_LFInst_15_LFInst_0_U4  ( .A(AddRoundKeyOutput[61]), .ZN(
        SubCellInst_LFInst_15_LFInst_0_n4 ) );
  XOR2_X1 SubCellInst_LFInst_15_LFInst_0_U3  ( .A(AddRoundKeyOutput[60]), .B(
        AddRoundKeyOutput[63]), .Z(SubCellInst_LFInst_15_LFInst_0_n6 ) );
  XNOR2_X1 MCInst1_MC0_v0_2Inst_0_U4  ( .A(MCInst1_MC0_v0_2Inst_0_n2 ), .B(
        MCInst1_MC0_v0_0 [3]), .ZN(MCInst1_MC0_v0_2 [0]) );
  XNOR2_X1 MCInst1_MC0_v0_2Inst_0_U3  ( .A(MCInst1_MC0_v0_3 [0]), .B(
        ShiftRowsOutput[60]), .ZN(MCInst1_MC0_v0_2Inst_0_n2 ) );
  XOR2_X1 MCInst1_MC0_v1_1Inst_0_U3  ( .A(MCInst1_MC0_v1_3 [3]), .B(
        MCInst1_MC0_v1_3 [0]), .Z(MCInst1_MC0_v1_1 [0]) );
  XNOR2_X1 MCInst1_MC0_v1_2Inst_0_U4  ( .A(MCInst1_MC0_v1_2Inst_0_n2 ), .B(
        MCInst1_MC0_v1_3 [3]), .ZN(MCInst1_MC0_v1_2 [0]) );
  XNOR2_X1 MCInst1_MC0_v1_2Inst_0_U3  ( .A(MCInst1_MC0_v1_3 [0]), .B(
        MCInst1_MC0_v1_3 [2]), .ZN(MCInst1_MC0_v1_2Inst_0_n2 ) );
  XOR2_X1 MCInst1_MC0_v2_1Inst_0_U3  ( .A(MCInst1_MC0_v2_3 [1]), .B(
        MCInst1_MC0_v2_0 [3]), .Z(MCInst1_MC0_v2_1 [0]) );
  XOR2_X1 MCInst1_MC0_v2_2Inst_0_U3  ( .A(MCInst1_MC0_v2_0 [2]), .B(
        MCInst1_MC0_v2_0 [0]), .Z(MCInst1_MC0_v2_2 [0]) );
  XNOR2_X1 MCInst1_MC0_v2_3Inst_0_U5  ( .A(MCInst1_MC0_v2_3Inst_0_n4 ), .B(
        MCInst1_MC0_v2_3Inst_0_n3 ), .ZN(MCInst1_MC0_v2_3 [0]) );
  XNOR2_X1 MCInst1_MC0_v2_3Inst_0_U4  ( .A(MCInst1_MC0_v2_0 [2]), .B(
        MCInst1_MC0_v2_3 [1]), .ZN(MCInst1_MC0_v2_3Inst_0_n3 ) );
  XOR2_X1 MCInst1_MC0_v2_3Inst_0_U3  ( .A(MCInst1_MC0_v2_0 [3]), .B(
        MCInst1_MC0_v2_0 [0]), .Z(MCInst1_MC0_v2_3Inst_0_n4 ) );
  XOR2_X1 MCInst1_MC0_v3_1Inst_0_U3  ( .A(MCInst1_MC0_v3_0 [3]), .B(
        MCInst1_MC0_v3_2 [2]), .Z(MCInst1_MC0_v3_1 [0]) );
  XOR2_X1 MCInst1_MC0_v3_2Inst_0_U3  ( .A(MCInst1_MC0_v3_2 [3]), .B(
        MCInst1_MC0_v3_0 [2]), .Z(MCInst1_MC0_v3_2 [0]) );
  XNOR2_X1 MCInst1_MC0_v3_3Inst_0_U4  ( .A(MCInst1_MC0_v3_3Inst_0_n2 ), .B(
        MCInst1_MC0_v3_0 [2]), .ZN(MCInst1_MC0_v3_3 [0]) );
  XNOR2_X1 MCInst1_MC0_v3_3Inst_0_U3  ( .A(MCInst1_MC0_v3_2 [2]), .B(
        MCInst1_MC0_v3_2 [3]), .ZN(MCInst1_MC0_v3_3Inst_0_n2 ) );
  XOR2_X1 MCInst1_MC0_v0_0Inst_1_U3  ( .A(MCInst1_MC0_v0_3 [3]), .B(
        MCInst1_MC0_v0_3 [0]), .Z(MCInst1_MC0_v0_0 [1]) );
  XOR2_X1 MCInst1_MC0_v0_1Inst_1_U3  ( .A(MCInst1_MC0_v0_0 [3]), .B(
        MCInst1_MC0_v0_3 [3]), .Z(MCInst1_MC0_v0_1 [1]) );
  XNOR2_X1 MCInst1_MC0_v0_2Inst_1_U4  ( .A(MCInst1_MC0_v0_2Inst_1_n2 ), .B(
        MCInst1_MC0_v0_3 [3]), .ZN(MCInst1_MC0_v0_2 [1]) );
  XNOR2_X1 MCInst1_MC0_v0_2Inst_1_U3  ( .A(MCInst1_MC0_v0_3 [0]), .B(
        ShiftRowsOutput[60]), .ZN(MCInst1_MC0_v0_2Inst_1_n2 ) );
  XOR2_X1 MCInst1_MC0_v0_3Inst_1_U3  ( .A(ShiftRowsOutput[60]), .B(
        MCInst1_MC0_v0_3 [0]), .Z(MCInst1_MC0_v0_3 [1]) );
  XOR2_X1 MCInst1_MC0_v1_1Inst_1_U3  ( .A(ShiftRowsOutput[44]), .B(
        MCInst1_MC0_v1_3 [3]), .Z(MCInst1_MC0_v1_1 [1]) );
  XOR2_X1 MCInst1_MC0_v1_2Inst_1_U3  ( .A(ShiftRowsOutput[44]), .B(
        MCInst1_MC0_v1_3 [2]), .Z(MCInst1_MC0_v1_2 [1]) );
  XOR2_X1 MCInst1_MC0_v1_3Inst_1_U3  ( .A(ShiftRowsOutput[44]), .B(
        MCInst1_MC0_v1_3 [0]), .Z(MCInst1_MC0_v1_3 [1]) );
  XOR2_X1 MCInst1_MC0_v2_0Inst_1_U3  ( .A(MCInst1_MC0_v2_3 [1]), .B(
        MCInst1_MC0_v2_0 [0]), .Z(MCInst1_MC0_v2_0 [1]) );
  XNOR2_X1 MCInst1_MC0_v2_1Inst_1_U4  ( .A(MCInst1_MC0_v2_1Inst_1_n2 ), .B(
        MCInst1_MC0_v2_0 [3]), .ZN(MCInst1_MC0_v2_1 [1]) );
  XNOR2_X1 MCInst1_MC0_v2_1Inst_1_U3  ( .A(MCInst1_MC0_v2_0 [0]), .B(
        MCInst1_MC0_v2_0 [2]), .ZN(MCInst1_MC0_v2_1Inst_1_n2 ) );
  XNOR2_X1 MCInst1_MC0_v2_2Inst_1_U5  ( .A(MCInst1_MC0_v2_2Inst_1_n4 ), .B(
        MCInst1_MC0_v2_2Inst_1_n3 ), .ZN(MCInst1_MC0_v2_2 [1]) );
  XNOR2_X1 MCInst1_MC0_v2_2Inst_1_U4  ( .A(MCInst1_MC0_v2_0 [2]), .B(
        MCInst1_MC0_v2_3 [1]), .ZN(MCInst1_MC0_v2_2Inst_1_n3 ) );
  XOR2_X1 MCInst1_MC0_v2_2Inst_1_U3  ( .A(MCInst1_MC0_v2_0 [3]), .B(
        MCInst1_MC0_v2_0 [0]), .Z(MCInst1_MC0_v2_2Inst_1_n4 ) );
  XOR2_X1 MCInst1_MC0_v3_0Inst_1_U3  ( .A(MCInst1_MC0_v3_2 [3]), .B(
        MCInst1_MC0_v3_2 [2]), .Z(MCInst1_MC0_v3_0 [1]) );
  XOR2_X1 MCInst1_MC0_v3_1Inst_1_U3  ( .A(MCInst1_MC0_v3_2 [3]), .B(
        MCInst1_MC0_v3_0 [3]), .Z(MCInst1_MC0_v3_1 [1]) );
  XNOR2_X1 MCInst1_MC0_v3_3Inst_1_U4  ( .A(MCInst1_MC0_v3_3Inst_1_n2 ), .B(
        MCInst1_MC0_v3_0 [3]), .ZN(MCInst1_MC0_v3_3 [1]) );
  XNOR2_X1 MCInst1_MC0_v3_3Inst_1_U3  ( .A(MCInst1_MC0_v3_2 [2]), .B(
        MCInst1_MC0_v3_2 [3]), .ZN(MCInst1_MC0_v3_3Inst_1_n2 ) );
  XOR2_X1 MCInst1_MC0_v0_0Inst_2_U3  ( .A(ShiftRowsOutput[60]), .B(
        MCInst1_MC0_v0_3 [0]), .Z(MCInst1_MC0_v0_0 [2]) );
  XOR2_X1 MCInst1_MC0_v0_1Inst_2_U3  ( .A(MCInst1_MC0_v0_3 [3]), .B(
        MCInst1_MC0_v0_3 [0]), .Z(MCInst1_MC0_v0_1 [2]) );
  XOR2_X1 MCInst1_MC0_v0_2Inst_2_U3  ( .A(MCInst1_MC0_v0_0 [3]), .B(
        MCInst1_MC0_v0_3 [0]), .Z(MCInst1_MC0_v0_2 [2]) );
  XNOR2_X1 MCInst1_MC0_v1_1Inst_2_U4  ( .A(MCInst1_MC0_v1_1Inst_2_n2 ), .B(
        MCInst1_MC0_v1_3 [2]), .ZN(MCInst1_MC0_v1_1 [2]) );
  XNOR2_X1 MCInst1_MC0_v1_1Inst_2_U3  ( .A(MCInst1_MC0_v1_3 [0]), .B(
        ShiftRowsOutput[44]), .ZN(MCInst1_MC0_v1_1Inst_2_n2 ) );
  XNOR2_X1 MCInst1_MC0_v1_2Inst_2_U4  ( .A(MCInst1_MC0_v1_2Inst_2_n2 ), .B(
        MCInst1_MC0_v1_3 [2]), .ZN(MCInst1_MC0_v1_2 [2]) );
  XNOR2_X1 MCInst1_MC0_v1_2Inst_2_U3  ( .A(MCInst1_MC0_v1_3 [3]), .B(
        ShiftRowsOutput[44]), .ZN(MCInst1_MC0_v1_2Inst_2_n2 ) );
  XNOR2_X1 MCInst1_MC0_v2_1Inst_2_U4  ( .A(MCInst1_MC0_v2_1Inst_2_n2 ), .B(
        MCInst1_MC0_v2_0 [3]), .ZN(MCInst1_MC0_v2_1 [2]) );
  XNOR2_X1 MCInst1_MC0_v2_1Inst_2_U3  ( .A(MCInst1_MC0_v2_0 [0]), .B(
        MCInst1_MC0_v2_3 [1]), .ZN(MCInst1_MC0_v2_1Inst_2_n2 ) );
  XNOR2_X1 MCInst1_MC0_v2_2Inst_2_U4  ( .A(MCInst1_MC0_v2_2Inst_2_n2 ), .B(
        MCInst1_MC0_v2_0 [3]), .ZN(MCInst1_MC0_v2_2 [2]) );
  XNOR2_X1 MCInst1_MC0_v2_2Inst_2_U3  ( .A(MCInst1_MC0_v2_0 [0]), .B(
        MCInst1_MC0_v2_0 [2]), .ZN(MCInst1_MC0_v2_2Inst_2_n2 ) );
  XOR2_X1 MCInst1_MC0_v2_3Inst_2_U3  ( .A(MCInst1_MC0_v2_3 [1]), .B(
        MCInst1_MC0_v2_0 [2]), .Z(MCInst1_MC0_v2_3 [2]) );
  XNOR2_X1 MCInst1_MC0_v3_1Inst_2_U4  ( .A(MCInst1_MC0_v3_1Inst_2_n2 ), .B(
        MCInst1_MC0_v3_0 [2]), .ZN(MCInst1_MC0_v3_1 [2]) );
  XNOR2_X1 MCInst1_MC0_v3_1Inst_2_U3  ( .A(MCInst1_MC0_v3_2 [2]), .B(
        MCInst1_MC0_v3_2 [3]), .ZN(MCInst1_MC0_v3_1Inst_2_n2 ) );
  XOR2_X1 MCInst1_MC0_v3_3Inst_2_U3  ( .A(MCInst1_MC0_v3_0 [2]), .B(
        MCInst1_MC0_v3_2 [2]), .Z(MCInst1_MC0_v3_3 [2]) );
  XOR2_X1 MCInst1_MC0_v0_1Inst_3_U3  ( .A(ShiftRowsOutput[60]), .B(
        MCInst1_MC0_v0_3 [0]), .Z(MCInst1_MC0_v0_1 [3]) );
  XOR2_X1 MCInst1_MC0_v0_2Inst_3_U3  ( .A(ShiftRowsOutput[60]), .B(
        MCInst1_MC0_v0_3 [3]), .Z(MCInst1_MC0_v0_2 [3]) );
  XOR2_X1 MCInst1_MC0_v1_1Inst_3_U3  ( .A(MCInst1_MC0_v1_3 [2]), .B(
        MCInst1_MC0_v1_3 [3]), .Z(MCInst1_MC0_v1_1 [3]) );
  XNOR2_X1 MCInst1_MC0_v1_2Inst_3_U5  ( .A(MCInst1_MC0_v1_2Inst_3_n4 ), .B(
        MCInst1_MC0_v1_2Inst_3_n3 ), .ZN(MCInst1_MC0_v1_2 [3]) );
  XNOR2_X1 MCInst1_MC0_v1_2Inst_3_U4  ( .A(MCInst1_MC0_v1_3 [2]), .B(
        ShiftRowsOutput[44]), .ZN(MCInst1_MC0_v1_2Inst_3_n3 ) );
  XOR2_X1 MCInst1_MC0_v1_2Inst_3_U3  ( .A(MCInst1_MC0_v1_3 [3]), .B(
        MCInst1_MC0_v1_3 [0]), .Z(MCInst1_MC0_v1_2Inst_3_n4 ) );
  XOR2_X1 MCInst1_MC0_v2_1Inst_3_U3  ( .A(MCInst1_MC0_v2_0 [2]), .B(
        MCInst1_MC0_v2_0 [0]), .Z(MCInst1_MC0_v2_1 [3]) );
  XNOR2_X1 MCInst1_MC0_v2_2Inst_3_U4  ( .A(MCInst1_MC0_v2_2Inst_3_n2 ), .B(
        MCInst1_MC0_v2_0 [3]), .ZN(MCInst1_MC0_v2_2 [3]) );
  XNOR2_X1 MCInst1_MC0_v2_2Inst_3_U3  ( .A(MCInst1_MC0_v2_0 [0]), .B(
        MCInst1_MC0_v2_3 [1]), .ZN(MCInst1_MC0_v2_2Inst_3_n2 ) );
  XNOR2_X1 MCInst1_MC0_v2_3Inst_3_U4  ( .A(MCInst1_MC0_v2_3Inst_3_n2 ), .B(
        MCInst1_MC0_v2_0 [2]), .ZN(MCInst1_MC0_v2_3 [3]) );
  XNOR2_X1 MCInst1_MC0_v2_3Inst_3_U3  ( .A(MCInst1_MC0_v2_0 [3]), .B(
        MCInst1_MC0_v2_3 [1]), .ZN(MCInst1_MC0_v2_3Inst_3_n2 ) );
  XOR2_X1 MCInst1_MC0_v3_1Inst_3_U3  ( .A(MCInst1_MC0_v3_0 [2]), .B(
        MCInst1_MC0_v3_0 [3]), .Z(MCInst1_MC0_v3_1 [3]) );
  XOR2_X1 MCInst1_MC0_v3_3Inst_3_U3  ( .A(MCInst1_MC0_v3_2 [3]), .B(
        MCInst1_MC0_v3_0 [3]), .Z(MCInst1_MC0_v3_3 [3]) );
  XNOR2_X1 MCInst1_MC0_r0Inst_XORInst_0_0_U3  ( .A(
        MCInst1_MC0_r0Inst_XORInst_0_0_n5 ), .B(
        MCInst1_MC0_r0Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[60]) );
  XNOR2_X1 MCInst1_MC0_r0Inst_XORInst_0_0_U2  ( .A(MCInst1_MC0_v3_2 [2]), 
        .B(MCInst1_MC0_v2_0 [0]), .ZN(MCInst1_MC0_r0Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst1_MC0_r0Inst_XORInst_0_0_U1  ( .A(MCInst1_MC0_v0_3 [3]), .B(
        ShiftRowsOutput[44]), .Z(MCInst1_MC0_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst1_MC0_r0Inst_XORInst_0_1_U3  ( .A(
        MCInst1_MC0_r0Inst_XORInst_0_1_n5 ), .B(
        MCInst1_MC0_r0Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[61]) );
  XNOR2_X1 MCInst1_MC0_r0Inst_XORInst_0_1_U2  ( .A(MCInst1_MC0_v3_0 [1]), 
        .B(MCInst1_MC0_v2_0 [1]), .ZN(MCInst1_MC0_r0Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst1_MC0_r0Inst_XORInst_0_1_U1  ( .A(MCInst1_MC0_v0_0 [1]), .B(
        MCInst1_MC0_v1_3 [2]), .Z(MCInst1_MC0_r0Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst1_MC0_r0Inst_XORInst_0_2_U3  ( .A(
        MCInst1_MC0_r0Inst_XORInst_0_2_n5 ), .B(
        MCInst1_MC0_r0Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[62]) );
  XNOR2_X1 MCInst1_MC0_r0Inst_XORInst_0_2_U2  ( .A(MCInst1_MC0_v3_0 [2]), 
        .B(MCInst1_MC0_v2_0 [2]), .ZN(MCInst1_MC0_r0Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst1_MC0_r0Inst_XORInst_0_2_U1  ( .A(MCInst1_MC0_v0_0 [2]), .B(
        MCInst1_MC0_v1_3 [3]), .Z(MCInst1_MC0_r0Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst1_MC0_r0Inst_XORInst_0_3_U3  ( .A(
        MCInst1_MC0_r0Inst_XORInst_0_3_n5 ), .B(
        MCInst1_MC0_r0Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[63]) );
  XNOR2_X1 MCInst1_MC0_r0Inst_XORInst_0_3_U2  ( .A(MCInst1_MC0_v3_0 [3]), 
        .B(MCInst1_MC0_v2_0 [3]), .ZN(MCInst1_MC0_r0Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst1_MC0_r0Inst_XORInst_0_3_U1  ( .A(MCInst1_MC0_v0_0 [3]), .B(
        MCInst1_MC0_v1_3 [0]), .Z(MCInst1_MC0_r0Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst1_MC0_r1Inst_XORInst_0_0_U3  ( .A(
        MCInst1_MC0_r1Inst_XORInst_0_0_n5 ), .B(
        MCInst1_MC0_r1Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[44]) );
  XNOR2_X1 MCInst1_MC0_r1Inst_XORInst_0_0_U2  ( .A(MCInst1_MC0_v3_1 [0]), 
        .B(MCInst1_MC0_v2_1 [0]), .ZN(MCInst1_MC0_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst1_MC0_r1Inst_XORInst_0_0_U1  ( .A(MCInst1_MC0_v0_0 [3]), .B(
        MCInst1_MC0_v1_1 [0]), .Z(MCInst1_MC0_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst1_MC0_r1Inst_XORInst_0_1_U3  ( .A(
        MCInst1_MC0_r1Inst_XORInst_0_1_n5 ), .B(
        MCInst1_MC0_r1Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[45]) );
  XNOR2_X1 MCInst1_MC0_r1Inst_XORInst_0_1_U2  ( .A(MCInst1_MC0_v3_1 [1]), 
        .B(MCInst1_MC0_v2_1 [1]), .ZN(MCInst1_MC0_r1Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst1_MC0_r1Inst_XORInst_0_1_U1  ( .A(MCInst1_MC0_v0_1 [1]), .B(
        MCInst1_MC0_v1_1 [1]), .Z(MCInst1_MC0_r1Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst1_MC0_r1Inst_XORInst_0_2_U3  ( .A(
        MCInst1_MC0_r1Inst_XORInst_0_2_n5 ), .B(
        MCInst1_MC0_r1Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[46]) );
  XNOR2_X1 MCInst1_MC0_r1Inst_XORInst_0_2_U2  ( .A(MCInst1_MC0_v3_1 [2]), 
        .B(MCInst1_MC0_v2_1 [2]), .ZN(MCInst1_MC0_r1Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst1_MC0_r1Inst_XORInst_0_2_U1  ( .A(MCInst1_MC0_v0_1 [2]), .B(
        MCInst1_MC0_v1_1 [2]), .Z(MCInst1_MC0_r1Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst1_MC0_r1Inst_XORInst_0_3_U3  ( .A(
        MCInst1_MC0_r1Inst_XORInst_0_3_n5 ), .B(
        MCInst1_MC0_r1Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[47]) );
  XNOR2_X1 MCInst1_MC0_r1Inst_XORInst_0_3_U2  ( .A(MCInst1_MC0_v3_1 [3]), 
        .B(MCInst1_MC0_v2_1 [3]), .ZN(MCInst1_MC0_r1Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst1_MC0_r1Inst_XORInst_0_3_U1  ( .A(MCInst1_MC0_v0_1 [3]), .B(
        MCInst1_MC0_v1_1 [3]), .Z(MCInst1_MC0_r1Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst1_MC0_r2Inst_XORInst_0_0_U3  ( .A(
        MCInst1_MC0_r2Inst_XORInst_0_0_n5 ), .B(
        MCInst1_MC0_r2Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[28]) );
  XNOR2_X1 MCInst1_MC0_r2Inst_XORInst_0_0_U2  ( .A(MCInst1_MC0_v3_2 [0]), 
        .B(MCInst1_MC0_v2_2 [0]), .ZN(MCInst1_MC0_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst1_MC0_r2Inst_XORInst_0_0_U1  ( .A(MCInst1_MC0_v0_2 [0]), .B(
        MCInst1_MC0_v1_2 [0]), .Z(MCInst1_MC0_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst1_MC0_r2Inst_XORInst_0_1_U3  ( .A(
        MCInst1_MC0_r2Inst_XORInst_0_1_n5 ), .B(
        MCInst1_MC0_r2Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[29]) );
  XNOR2_X1 MCInst1_MC0_r2Inst_XORInst_0_1_U2  ( .A(MCInst1_MC0_v3_0 [3]), 
        .B(MCInst1_MC0_v2_2 [1]), .ZN(MCInst1_MC0_r2Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst1_MC0_r2Inst_XORInst_0_1_U1  ( .A(MCInst1_MC0_v0_2 [1]), .B(
        MCInst1_MC0_v1_2 [1]), .Z(MCInst1_MC0_r2Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst1_MC0_r2Inst_XORInst_0_2_U3  ( .A(
        MCInst1_MC0_r2Inst_XORInst_0_2_n5 ), .B(
        MCInst1_MC0_r2Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[30]) );
  XNOR2_X1 MCInst1_MC0_r2Inst_XORInst_0_2_U2  ( .A(MCInst1_MC0_v3_2 [2]), 
        .B(MCInst1_MC0_v2_2 [2]), .ZN(MCInst1_MC0_r2Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst1_MC0_r2Inst_XORInst_0_2_U1  ( .A(MCInst1_MC0_v0_2 [2]), .B(
        MCInst1_MC0_v1_2 [2]), .Z(MCInst1_MC0_r2Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst1_MC0_r2Inst_XORInst_0_3_U3  ( .A(
        MCInst1_MC0_r2Inst_XORInst_0_3_n5 ), .B(
        MCInst1_MC0_r2Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[31]) );
  XNOR2_X1 MCInst1_MC0_r2Inst_XORInst_0_3_U2  ( .A(MCInst1_MC0_v3_2 [3]), 
        .B(MCInst1_MC0_v2_2 [3]), .ZN(MCInst1_MC0_r2Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst1_MC0_r2Inst_XORInst_0_3_U1  ( .A(MCInst1_MC0_v0_2 [3]), .B(
        MCInst1_MC0_v1_2 [3]), .Z(MCInst1_MC0_r2Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst1_MC0_r3Inst_XORInst_0_0_U3  ( .A(
        MCInst1_MC0_r3Inst_XORInst_0_0_n5 ), .B(
        MCInst1_MC0_r3Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[12]) );
  XNOR2_X1 MCInst1_MC0_r3Inst_XORInst_0_0_U2  ( .A(MCInst1_MC0_v3_3 [0]), 
        .B(MCInst1_MC0_v2_3 [0]), .ZN(MCInst1_MC0_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst1_MC0_r3Inst_XORInst_0_0_U1  ( .A(MCInst1_MC0_v0_3 [0]), .B(
        MCInst1_MC0_v1_3 [0]), .Z(MCInst1_MC0_r3Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst1_MC0_r3Inst_XORInst_0_1_U3  ( .A(
        MCInst1_MC0_r3Inst_XORInst_0_1_n5 ), .B(
        MCInst1_MC0_r3Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[13]) );
  XNOR2_X1 MCInst1_MC0_r3Inst_XORInst_0_1_U2  ( .A(MCInst1_MC0_v3_3 [1]), 
        .B(MCInst1_MC0_v2_3 [1]), .ZN(MCInst1_MC0_r3Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst1_MC0_r3Inst_XORInst_0_1_U1  ( .A(MCInst1_MC0_v0_3 [1]), .B(
        MCInst1_MC0_v1_3 [1]), .Z(MCInst1_MC0_r3Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst1_MC0_r3Inst_XORInst_0_2_U3  ( .A(
        MCInst1_MC0_r3Inst_XORInst_0_2_n5 ), .B(
        MCInst1_MC0_r3Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[14]) );
  XNOR2_X1 MCInst1_MC0_r3Inst_XORInst_0_2_U2  ( .A(MCInst1_MC0_v3_3 [2]), 
        .B(MCInst1_MC0_v2_3 [2]), .ZN(MCInst1_MC0_r3Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst1_MC0_r3Inst_XORInst_0_2_U1  ( .A(MCInst1_MC0_v0_0 [3]), .B(
        MCInst1_MC0_v1_3 [2]), .Z(MCInst1_MC0_r3Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst1_MC0_r3Inst_XORInst_0_3_U3  ( .A(
        MCInst1_MC0_r3Inst_XORInst_0_3_n5 ), .B(
        MCInst1_MC0_r3Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[15]) );
  XNOR2_X1 MCInst1_MC0_r3Inst_XORInst_0_3_U2  ( .A(MCInst1_MC0_v3_3 [3]), 
        .B(MCInst1_MC0_v2_3 [3]), .ZN(MCInst1_MC0_r3Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst1_MC0_r3Inst_XORInst_0_3_U1  ( .A(MCInst1_MC0_v0_3 [3]), .B(
        MCInst1_MC0_v1_3 [3]), .Z(MCInst1_MC0_r3Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst1_MC1_v0_2Inst_0_U4  ( .A(MCInst1_MC1_v0_2Inst_0_n2 ), .B(
        MCInst1_MC1_v0_0 [3]), .ZN(MCInst1_MC1_v0_2 [0]) );
  XNOR2_X1 MCInst1_MC1_v0_2Inst_0_U3  ( .A(MCInst1_MC1_v0_3 [0]), .B(
        ShiftRowsOutput[56]), .ZN(MCInst1_MC1_v0_2Inst_0_n2 ) );
  XOR2_X1 MCInst1_MC1_v1_1Inst_0_U3  ( .A(MCInst1_MC1_v1_3 [3]), .B(
        MCInst1_MC1_v1_3 [0]), .Z(MCInst1_MC1_v1_1 [0]) );
  XNOR2_X1 MCInst1_MC1_v1_2Inst_0_U4  ( .A(MCInst1_MC1_v1_2Inst_0_n2 ), .B(
        MCInst1_MC1_v1_3 [3]), .ZN(MCInst1_MC1_v1_2 [0]) );
  XNOR2_X1 MCInst1_MC1_v1_2Inst_0_U3  ( .A(MCInst1_MC1_v1_3 [0]), .B(
        MCInst1_MC1_v1_3 [2]), .ZN(MCInst1_MC1_v1_2Inst_0_n2 ) );
  XOR2_X1 MCInst1_MC1_v2_1Inst_0_U3  ( .A(MCInst1_MC1_v2_3 [1]), .B(
        MCInst1_MC1_v2_0 [3]), .Z(MCInst1_MC1_v2_1 [0]) );
  XOR2_X1 MCInst1_MC1_v2_2Inst_0_U3  ( .A(MCInst1_MC1_v2_0 [2]), .B(
        MCInst1_MC1_v2_0 [0]), .Z(MCInst1_MC1_v2_2 [0]) );
  XNOR2_X1 MCInst1_MC1_v2_3Inst_0_U5  ( .A(MCInst1_MC1_v2_3Inst_0_n4 ), .B(
        MCInst1_MC1_v2_3Inst_0_n3 ), .ZN(MCInst1_MC1_v2_3 [0]) );
  XNOR2_X1 MCInst1_MC1_v2_3Inst_0_U4  ( .A(MCInst1_MC1_v2_0 [2]), .B(
        MCInst1_MC1_v2_3 [1]), .ZN(MCInst1_MC1_v2_3Inst_0_n3 ) );
  XOR2_X1 MCInst1_MC1_v2_3Inst_0_U3  ( .A(MCInst1_MC1_v2_0 [3]), .B(
        MCInst1_MC1_v2_0 [0]), .Z(MCInst1_MC1_v2_3Inst_0_n4 ) );
  XOR2_X1 MCInst1_MC1_v3_1Inst_0_U3  ( .A(MCInst1_MC1_v3_0 [3]), .B(
        MCInst1_MC1_v3_2 [2]), .Z(MCInst1_MC1_v3_1 [0]) );
  XOR2_X1 MCInst1_MC1_v3_2Inst_0_U3  ( .A(MCInst1_MC1_v3_2 [3]), .B(
        MCInst1_MC1_v3_0 [2]), .Z(MCInst1_MC1_v3_2 [0]) );
  XNOR2_X1 MCInst1_MC1_v3_3Inst_0_U4  ( .A(MCInst1_MC1_v3_3Inst_0_n2 ), .B(
        MCInst1_MC1_v3_0 [2]), .ZN(MCInst1_MC1_v3_3 [0]) );
  XNOR2_X1 MCInst1_MC1_v3_3Inst_0_U3  ( .A(MCInst1_MC1_v3_2 [2]), .B(
        MCInst1_MC1_v3_2 [3]), .ZN(MCInst1_MC1_v3_3Inst_0_n2 ) );
  XOR2_X1 MCInst1_MC1_v0_0Inst_1_U3  ( .A(MCInst1_MC1_v0_3 [3]), .B(
        MCInst1_MC1_v0_3 [0]), .Z(MCInst1_MC1_v0_0 [1]) );
  XOR2_X1 MCInst1_MC1_v0_1Inst_1_U3  ( .A(MCInst1_MC1_v0_0 [3]), .B(
        MCInst1_MC1_v0_3 [3]), .Z(MCInst1_MC1_v0_1 [1]) );
  XNOR2_X1 MCInst1_MC1_v0_2Inst_1_U4  ( .A(MCInst1_MC1_v0_2Inst_1_n2 ), .B(
        MCInst1_MC1_v0_3 [3]), .ZN(MCInst1_MC1_v0_2 [1]) );
  XNOR2_X1 MCInst1_MC1_v0_2Inst_1_U3  ( .A(MCInst1_MC1_v0_3 [0]), .B(
        ShiftRowsOutput[56]), .ZN(MCInst1_MC1_v0_2Inst_1_n2 ) );
  XOR2_X1 MCInst1_MC1_v0_3Inst_1_U3  ( .A(ShiftRowsOutput[56]), .B(
        MCInst1_MC1_v0_3 [0]), .Z(MCInst1_MC1_v0_3 [1]) );
  XOR2_X1 MCInst1_MC1_v1_1Inst_1_U3  ( .A(ShiftRowsOutput[40]), .B(
        MCInst1_MC1_v1_3 [3]), .Z(MCInst1_MC1_v1_1 [1]) );
  XOR2_X1 MCInst1_MC1_v1_2Inst_1_U3  ( .A(ShiftRowsOutput[40]), .B(
        MCInst1_MC1_v1_3 [2]), .Z(MCInst1_MC1_v1_2 [1]) );
  XOR2_X1 MCInst1_MC1_v1_3Inst_1_U3  ( .A(ShiftRowsOutput[40]), .B(
        MCInst1_MC1_v1_3 [0]), .Z(MCInst1_MC1_v1_3 [1]) );
  XOR2_X1 MCInst1_MC1_v2_0Inst_1_U3  ( .A(MCInst1_MC1_v2_3 [1]), .B(
        MCInst1_MC1_v2_0 [0]), .Z(MCInst1_MC1_v2_0 [1]) );
  XNOR2_X1 MCInst1_MC1_v2_1Inst_1_U4  ( .A(MCInst1_MC1_v2_1Inst_1_n2 ), .B(
        MCInst1_MC1_v2_0 [3]), .ZN(MCInst1_MC1_v2_1 [1]) );
  XNOR2_X1 MCInst1_MC1_v2_1Inst_1_U3  ( .A(MCInst1_MC1_v2_0 [0]), .B(
        MCInst1_MC1_v2_0 [2]), .ZN(MCInst1_MC1_v2_1Inst_1_n2 ) );
  XNOR2_X1 MCInst1_MC1_v2_2Inst_1_U5  ( .A(MCInst1_MC1_v2_2Inst_1_n4 ), .B(
        MCInst1_MC1_v2_2Inst_1_n3 ), .ZN(MCInst1_MC1_v2_2 [1]) );
  XNOR2_X1 MCInst1_MC1_v2_2Inst_1_U4  ( .A(MCInst1_MC1_v2_0 [2]), .B(
        MCInst1_MC1_v2_3 [1]), .ZN(MCInst1_MC1_v2_2Inst_1_n3 ) );
  XOR2_X1 MCInst1_MC1_v2_2Inst_1_U3  ( .A(MCInst1_MC1_v2_0 [3]), .B(
        MCInst1_MC1_v2_0 [0]), .Z(MCInst1_MC1_v2_2Inst_1_n4 ) );
  XOR2_X1 MCInst1_MC1_v3_0Inst_1_U3  ( .A(MCInst1_MC1_v3_2 [3]), .B(
        MCInst1_MC1_v3_2 [2]), .Z(MCInst1_MC1_v3_0 [1]) );
  XOR2_X1 MCInst1_MC1_v3_1Inst_1_U3  ( .A(MCInst1_MC1_v3_2 [3]), .B(
        MCInst1_MC1_v3_0 [3]), .Z(MCInst1_MC1_v3_1 [1]) );
  XNOR2_X1 MCInst1_MC1_v3_3Inst_1_U4  ( .A(MCInst1_MC1_v3_3Inst_1_n2 ), .B(
        MCInst1_MC1_v3_0 [3]), .ZN(MCInst1_MC1_v3_3 [1]) );
  XNOR2_X1 MCInst1_MC1_v3_3Inst_1_U3  ( .A(MCInst1_MC1_v3_2 [2]), .B(
        MCInst1_MC1_v3_2 [3]), .ZN(MCInst1_MC1_v3_3Inst_1_n2 ) );
  XOR2_X1 MCInst1_MC1_v0_0Inst_2_U3  ( .A(ShiftRowsOutput[56]), .B(
        MCInst1_MC1_v0_3 [0]), .Z(MCInst1_MC1_v0_0 [2]) );
  XOR2_X1 MCInst1_MC1_v0_1Inst_2_U3  ( .A(MCInst1_MC1_v0_3 [3]), .B(
        MCInst1_MC1_v0_3 [0]), .Z(MCInst1_MC1_v0_1 [2]) );
  XOR2_X1 MCInst1_MC1_v0_2Inst_2_U3  ( .A(MCInst1_MC1_v0_0 [3]), .B(
        MCInst1_MC1_v0_3 [0]), .Z(MCInst1_MC1_v0_2 [2]) );
  XNOR2_X1 MCInst1_MC1_v1_1Inst_2_U4  ( .A(MCInst1_MC1_v1_1Inst_2_n2 ), .B(
        MCInst1_MC1_v1_3 [2]), .ZN(MCInst1_MC1_v1_1 [2]) );
  XNOR2_X1 MCInst1_MC1_v1_1Inst_2_U3  ( .A(MCInst1_MC1_v1_3 [0]), .B(
        ShiftRowsOutput[40]), .ZN(MCInst1_MC1_v1_1Inst_2_n2 ) );
  XNOR2_X1 MCInst1_MC1_v1_2Inst_2_U4  ( .A(MCInst1_MC1_v1_2Inst_2_n2 ), .B(
        MCInst1_MC1_v1_3 [2]), .ZN(MCInst1_MC1_v1_2 [2]) );
  XNOR2_X1 MCInst1_MC1_v1_2Inst_2_U3  ( .A(MCInst1_MC1_v1_3 [3]), .B(
        ShiftRowsOutput[40]), .ZN(MCInst1_MC1_v1_2Inst_2_n2 ) );
  XNOR2_X1 MCInst1_MC1_v2_1Inst_2_U4  ( .A(MCInst1_MC1_v2_1Inst_2_n2 ), .B(
        MCInst1_MC1_v2_0 [3]), .ZN(MCInst1_MC1_v2_1 [2]) );
  XNOR2_X1 MCInst1_MC1_v2_1Inst_2_U3  ( .A(MCInst1_MC1_v2_0 [0]), .B(
        MCInst1_MC1_v2_3 [1]), .ZN(MCInst1_MC1_v2_1Inst_2_n2 ) );
  XNOR2_X1 MCInst1_MC1_v2_2Inst_2_U4  ( .A(MCInst1_MC1_v2_2Inst_2_n2 ), .B(
        MCInst1_MC1_v2_0 [3]), .ZN(MCInst1_MC1_v2_2 [2]) );
  XNOR2_X1 MCInst1_MC1_v2_2Inst_2_U3  ( .A(MCInst1_MC1_v2_0 [0]), .B(
        MCInst1_MC1_v2_0 [2]), .ZN(MCInst1_MC1_v2_2Inst_2_n2 ) );
  XOR2_X1 MCInst1_MC1_v2_3Inst_2_U3  ( .A(MCInst1_MC1_v2_3 [1]), .B(
        MCInst1_MC1_v2_0 [2]), .Z(MCInst1_MC1_v2_3 [2]) );
  XNOR2_X1 MCInst1_MC1_v3_1Inst_2_U4  ( .A(MCInst1_MC1_v3_1Inst_2_n2 ), .B(
        MCInst1_MC1_v3_0 [2]), .ZN(MCInst1_MC1_v3_1 [2]) );
  XNOR2_X1 MCInst1_MC1_v3_1Inst_2_U3  ( .A(MCInst1_MC1_v3_2 [2]), .B(
        MCInst1_MC1_v3_2 [3]), .ZN(MCInst1_MC1_v3_1Inst_2_n2 ) );
  XOR2_X1 MCInst1_MC1_v3_3Inst_2_U3  ( .A(MCInst1_MC1_v3_0 [2]), .B(
        MCInst1_MC1_v3_2 [2]), .Z(MCInst1_MC1_v3_3 [2]) );
  XOR2_X1 MCInst1_MC1_v0_1Inst_3_U3  ( .A(ShiftRowsOutput[56]), .B(
        MCInst1_MC1_v0_3 [0]), .Z(MCInst1_MC1_v0_1 [3]) );
  XOR2_X1 MCInst1_MC1_v0_2Inst_3_U3  ( .A(ShiftRowsOutput[56]), .B(
        MCInst1_MC1_v0_3 [3]), .Z(MCInst1_MC1_v0_2 [3]) );
  XOR2_X1 MCInst1_MC1_v1_1Inst_3_U3  ( .A(MCInst1_MC1_v1_3 [2]), .B(
        MCInst1_MC1_v1_3 [3]), .Z(MCInst1_MC1_v1_1 [3]) );
  XNOR2_X1 MCInst1_MC1_v1_2Inst_3_U5  ( .A(MCInst1_MC1_v1_2Inst_3_n4 ), .B(
        MCInst1_MC1_v1_2Inst_3_n3 ), .ZN(MCInst1_MC1_v1_2 [3]) );
  XNOR2_X1 MCInst1_MC1_v1_2Inst_3_U4  ( .A(MCInst1_MC1_v1_3 [2]), .B(
        ShiftRowsOutput[40]), .ZN(MCInst1_MC1_v1_2Inst_3_n3 ) );
  XOR2_X1 MCInst1_MC1_v1_2Inst_3_U3  ( .A(MCInst1_MC1_v1_3 [3]), .B(
        MCInst1_MC1_v1_3 [0]), .Z(MCInst1_MC1_v1_2Inst_3_n4 ) );
  XOR2_X1 MCInst1_MC1_v2_1Inst_3_U3  ( .A(MCInst1_MC1_v2_0 [2]), .B(
        MCInst1_MC1_v2_0 [0]), .Z(MCInst1_MC1_v2_1 [3]) );
  XNOR2_X1 MCInst1_MC1_v2_2Inst_3_U4  ( .A(MCInst1_MC1_v2_2Inst_3_n2 ), .B(
        MCInst1_MC1_v2_0 [3]), .ZN(MCInst1_MC1_v2_2 [3]) );
  XNOR2_X1 MCInst1_MC1_v2_2Inst_3_U3  ( .A(MCInst1_MC1_v2_0 [0]), .B(
        MCInst1_MC1_v2_3 [1]), .ZN(MCInst1_MC1_v2_2Inst_3_n2 ) );
  XNOR2_X1 MCInst1_MC1_v2_3Inst_3_U4  ( .A(MCInst1_MC1_v2_3Inst_3_n2 ), .B(
        MCInst1_MC1_v2_0 [2]), .ZN(MCInst1_MC1_v2_3 [3]) );
  XNOR2_X1 MCInst1_MC1_v2_3Inst_3_U3  ( .A(MCInst1_MC1_v2_0 [3]), .B(
        MCInst1_MC1_v2_3 [1]), .ZN(MCInst1_MC1_v2_3Inst_3_n2 ) );
  XOR2_X1 MCInst1_MC1_v3_1Inst_3_U3  ( .A(MCInst1_MC1_v3_0 [2]), .B(
        MCInst1_MC1_v3_0 [3]), .Z(MCInst1_MC1_v3_1 [3]) );
  XOR2_X1 MCInst1_MC1_v3_3Inst_3_U3  ( .A(MCInst1_MC1_v3_2 [3]), .B(
        MCInst1_MC1_v3_0 [3]), .Z(MCInst1_MC1_v3_3 [3]) );
  XNOR2_X1 MCInst1_MC1_r0Inst_XORInst_0_0_U3  ( .A(
        MCInst1_MC1_r0Inst_XORInst_0_0_n5 ), .B(
        MCInst1_MC1_r0Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[56]) );
  XNOR2_X1 MCInst1_MC1_r0Inst_XORInst_0_0_U2  ( .A(MCInst1_MC1_v3_2 [2]), 
        .B(MCInst1_MC1_v2_0 [0]), .ZN(MCInst1_MC1_r0Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst1_MC1_r0Inst_XORInst_0_0_U1  ( .A(MCInst1_MC1_v0_3 [3]), .B(
        ShiftRowsOutput[40]), .Z(MCInst1_MC1_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst1_MC1_r0Inst_XORInst_0_1_U3  ( .A(
        MCInst1_MC1_r0Inst_XORInst_0_1_n5 ), .B(
        MCInst1_MC1_r0Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[57]) );
  XNOR2_X1 MCInst1_MC1_r0Inst_XORInst_0_1_U2  ( .A(MCInst1_MC1_v3_0 [1]), 
        .B(MCInst1_MC1_v2_0 [1]), .ZN(MCInst1_MC1_r0Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst1_MC1_r0Inst_XORInst_0_1_U1  ( .A(MCInst1_MC1_v0_0 [1]), .B(
        MCInst1_MC1_v1_3 [2]), .Z(MCInst1_MC1_r0Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst1_MC1_r0Inst_XORInst_0_2_U3  ( .A(
        MCInst1_MC1_r0Inst_XORInst_0_2_n5 ), .B(
        MCInst1_MC1_r0Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[58]) );
  XNOR2_X1 MCInst1_MC1_r0Inst_XORInst_0_2_U2  ( .A(MCInst1_MC1_v3_0 [2]), 
        .B(MCInst1_MC1_v2_0 [2]), .ZN(MCInst1_MC1_r0Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst1_MC1_r0Inst_XORInst_0_2_U1  ( .A(MCInst1_MC1_v0_0 [2]), .B(
        MCInst1_MC1_v1_3 [3]), .Z(MCInst1_MC1_r0Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst1_MC1_r0Inst_XORInst_0_3_U3  ( .A(
        MCInst1_MC1_r0Inst_XORInst_0_3_n5 ), .B(
        MCInst1_MC1_r0Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[59]) );
  XNOR2_X1 MCInst1_MC1_r0Inst_XORInst_0_3_U2  ( .A(MCInst1_MC1_v3_0 [3]), 
        .B(MCInst1_MC1_v2_0 [3]), .ZN(MCInst1_MC1_r0Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst1_MC1_r0Inst_XORInst_0_3_U1  ( .A(MCInst1_MC1_v0_0 [3]), .B(
        MCInst1_MC1_v1_3 [0]), .Z(MCInst1_MC1_r0Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst1_MC1_r1Inst_XORInst_0_0_U3  ( .A(
        MCInst1_MC1_r1Inst_XORInst_0_0_n5 ), .B(
        MCInst1_MC1_r1Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[40]) );
  XNOR2_X1 MCInst1_MC1_r1Inst_XORInst_0_0_U2  ( .A(MCInst1_MC1_v3_1 [0]), 
        .B(MCInst1_MC1_v2_1 [0]), .ZN(MCInst1_MC1_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst1_MC1_r1Inst_XORInst_0_0_U1  ( .A(MCInst1_MC1_v0_0 [3]), .B(
        MCInst1_MC1_v1_1 [0]), .Z(MCInst1_MC1_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst1_MC1_r1Inst_XORInst_0_1_U3  ( .A(
        MCInst1_MC1_r1Inst_XORInst_0_1_n5 ), .B(
        MCInst1_MC1_r1Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[41]) );
  XNOR2_X1 MCInst1_MC1_r1Inst_XORInst_0_1_U2  ( .A(MCInst1_MC1_v3_1 [1]), 
        .B(MCInst1_MC1_v2_1 [1]), .ZN(MCInst1_MC1_r1Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst1_MC1_r1Inst_XORInst_0_1_U1  ( .A(MCInst1_MC1_v0_1 [1]), .B(
        MCInst1_MC1_v1_1 [1]), .Z(MCInst1_MC1_r1Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst1_MC1_r1Inst_XORInst_0_2_U3  ( .A(
        MCInst1_MC1_r1Inst_XORInst_0_2_n5 ), .B(
        MCInst1_MC1_r1Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[42]) );
  XNOR2_X1 MCInst1_MC1_r1Inst_XORInst_0_2_U2  ( .A(MCInst1_MC1_v3_1 [2]), 
        .B(MCInst1_MC1_v2_1 [2]), .ZN(MCInst1_MC1_r1Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst1_MC1_r1Inst_XORInst_0_2_U1  ( .A(MCInst1_MC1_v0_1 [2]), .B(
        MCInst1_MC1_v1_1 [2]), .Z(MCInst1_MC1_r1Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst1_MC1_r1Inst_XORInst_0_3_U3  ( .A(
        MCInst1_MC1_r1Inst_XORInst_0_3_n5 ), .B(
        MCInst1_MC1_r1Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[43]) );
  XNOR2_X1 MCInst1_MC1_r1Inst_XORInst_0_3_U2  ( .A(MCInst1_MC1_v3_1 [3]), 
        .B(MCInst1_MC1_v2_1 [3]), .ZN(MCInst1_MC1_r1Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst1_MC1_r1Inst_XORInst_0_3_U1  ( .A(MCInst1_MC1_v0_1 [3]), .B(
        MCInst1_MC1_v1_1 [3]), .Z(MCInst1_MC1_r1Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst1_MC1_r2Inst_XORInst_0_0_U3  ( .A(
        MCInst1_MC1_r2Inst_XORInst_0_0_n5 ), .B(
        MCInst1_MC1_r2Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[24]) );
  XNOR2_X1 MCInst1_MC1_r2Inst_XORInst_0_0_U2  ( .A(MCInst1_MC1_v3_2 [0]), 
        .B(MCInst1_MC1_v2_2 [0]), .ZN(MCInst1_MC1_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst1_MC1_r2Inst_XORInst_0_0_U1  ( .A(MCInst1_MC1_v0_2 [0]), .B(
        MCInst1_MC1_v1_2 [0]), .Z(MCInst1_MC1_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst1_MC1_r2Inst_XORInst_0_1_U3  ( .A(
        MCInst1_MC1_r2Inst_XORInst_0_1_n5 ), .B(
        MCInst1_MC1_r2Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[25]) );
  XNOR2_X1 MCInst1_MC1_r2Inst_XORInst_0_1_U2  ( .A(MCInst1_MC1_v3_0 [3]), 
        .B(MCInst1_MC1_v2_2 [1]), .ZN(MCInst1_MC1_r2Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst1_MC1_r2Inst_XORInst_0_1_U1  ( .A(MCInst1_MC1_v0_2 [1]), .B(
        MCInst1_MC1_v1_2 [1]), .Z(MCInst1_MC1_r2Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst1_MC1_r2Inst_XORInst_0_2_U3  ( .A(
        MCInst1_MC1_r2Inst_XORInst_0_2_n5 ), .B(
        MCInst1_MC1_r2Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[26]) );
  XNOR2_X1 MCInst1_MC1_r2Inst_XORInst_0_2_U2  ( .A(MCInst1_MC1_v3_2 [2]), 
        .B(MCInst1_MC1_v2_2 [2]), .ZN(MCInst1_MC1_r2Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst1_MC1_r2Inst_XORInst_0_2_U1  ( .A(MCInst1_MC1_v0_2 [2]), .B(
        MCInst1_MC1_v1_2 [2]), .Z(MCInst1_MC1_r2Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst1_MC1_r2Inst_XORInst_0_3_U3  ( .A(
        MCInst1_MC1_r2Inst_XORInst_0_3_n5 ), .B(
        MCInst1_MC1_r2Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[27]) );
  XNOR2_X1 MCInst1_MC1_r2Inst_XORInst_0_3_U2  ( .A(MCInst1_MC1_v3_2 [3]), 
        .B(MCInst1_MC1_v2_2 [3]), .ZN(MCInst1_MC1_r2Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst1_MC1_r2Inst_XORInst_0_3_U1  ( .A(MCInst1_MC1_v0_2 [3]), .B(
        MCInst1_MC1_v1_2 [3]), .Z(MCInst1_MC1_r2Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst1_MC1_r3Inst_XORInst_0_0_U3  ( .A(
        MCInst1_MC1_r3Inst_XORInst_0_0_n5 ), .B(
        MCInst1_MC1_r3Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[8]) );
  XNOR2_X1 MCInst1_MC1_r3Inst_XORInst_0_0_U2  ( .A(MCInst1_MC1_v3_3 [0]), 
        .B(MCInst1_MC1_v2_3 [0]), .ZN(MCInst1_MC1_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst1_MC1_r3Inst_XORInst_0_0_U1  ( .A(MCInst1_MC1_v0_3 [0]), .B(
        MCInst1_MC1_v1_3 [0]), .Z(MCInst1_MC1_r3Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst1_MC1_r3Inst_XORInst_0_1_U3  ( .A(
        MCInst1_MC1_r3Inst_XORInst_0_1_n5 ), .B(
        MCInst1_MC1_r3Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[9]) );
  XNOR2_X1 MCInst1_MC1_r3Inst_XORInst_0_1_U2  ( .A(MCInst1_MC1_v3_3 [1]), 
        .B(MCInst1_MC1_v2_3 [1]), .ZN(MCInst1_MC1_r3Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst1_MC1_r3Inst_XORInst_0_1_U1  ( .A(MCInst1_MC1_v0_3 [1]), .B(
        MCInst1_MC1_v1_3 [1]), .Z(MCInst1_MC1_r3Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst1_MC1_r3Inst_XORInst_0_2_U3  ( .A(
        MCInst1_MC1_r3Inst_XORInst_0_2_n5 ), .B(
        MCInst1_MC1_r3Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[10]) );
  XNOR2_X1 MCInst1_MC1_r3Inst_XORInst_0_2_U2  ( .A(MCInst1_MC1_v3_3 [2]), 
        .B(MCInst1_MC1_v2_3 [2]), .ZN(MCInst1_MC1_r3Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst1_MC1_r3Inst_XORInst_0_2_U1  ( .A(MCInst1_MC1_v0_0 [3]), .B(
        MCInst1_MC1_v1_3 [2]), .Z(MCInst1_MC1_r3Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst1_MC1_r3Inst_XORInst_0_3_U3  ( .A(
        MCInst1_MC1_r3Inst_XORInst_0_3_n5 ), .B(
        MCInst1_MC1_r3Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[11]) );
  XNOR2_X1 MCInst1_MC1_r3Inst_XORInst_0_3_U2  ( .A(MCInst1_MC1_v3_3 [3]), 
        .B(MCInst1_MC1_v2_3 [3]), .ZN(MCInst1_MC1_r3Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst1_MC1_r3Inst_XORInst_0_3_U1  ( .A(MCInst1_MC1_v0_3 [3]), .B(
        MCInst1_MC1_v1_3 [3]), .Z(MCInst1_MC1_r3Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst1_MC2_v0_2Inst_0_U4  ( .A(MCInst1_MC2_v0_2Inst_0_n2 ), .B(
        MCInst1_MC2_v0_0 [3]), .ZN(MCInst1_MC2_v0_2 [0]) );
  XNOR2_X1 MCInst1_MC2_v0_2Inst_0_U3  ( .A(MCInst1_MC2_v0_3 [0]), .B(
        ShiftRowsOutput[52]), .ZN(MCInst1_MC2_v0_2Inst_0_n2 ) );
  XOR2_X1 MCInst1_MC2_v1_1Inst_0_U3  ( .A(MCInst1_MC2_v1_3 [3]), .B(
        MCInst1_MC2_v1_3 [0]), .Z(MCInst1_MC2_v1_1 [0]) );
  XNOR2_X1 MCInst1_MC2_v1_2Inst_0_U4  ( .A(MCInst1_MC2_v1_2Inst_0_n2 ), .B(
        MCInst1_MC2_v1_3 [3]), .ZN(MCInst1_MC2_v1_2 [0]) );
  XNOR2_X1 MCInst1_MC2_v1_2Inst_0_U3  ( .A(MCInst1_MC2_v1_3 [0]), .B(
        MCInst1_MC2_v1_3 [2]), .ZN(MCInst1_MC2_v1_2Inst_0_n2 ) );
  XOR2_X1 MCInst1_MC2_v2_1Inst_0_U3  ( .A(MCInst1_MC2_v2_3 [1]), .B(
        MCInst1_MC2_v2_0 [3]), .Z(MCInst1_MC2_v2_1 [0]) );
  XOR2_X1 MCInst1_MC2_v2_2Inst_0_U3  ( .A(MCInst1_MC2_v2_0 [2]), .B(
        MCInst1_MC2_v2_0 [0]), .Z(MCInst1_MC2_v2_2 [0]) );
  XNOR2_X1 MCInst1_MC2_v2_3Inst_0_U5  ( .A(MCInst1_MC2_v2_3Inst_0_n4 ), .B(
        MCInst1_MC2_v2_3Inst_0_n3 ), .ZN(MCInst1_MC2_v2_3 [0]) );
  XNOR2_X1 MCInst1_MC2_v2_3Inst_0_U4  ( .A(MCInst1_MC2_v2_0 [2]), .B(
        MCInst1_MC2_v2_3 [1]), .ZN(MCInst1_MC2_v2_3Inst_0_n3 ) );
  XOR2_X1 MCInst1_MC2_v2_3Inst_0_U3  ( .A(MCInst1_MC2_v2_0 [3]), .B(
        MCInst1_MC2_v2_0 [0]), .Z(MCInst1_MC2_v2_3Inst_0_n4 ) );
  XOR2_X1 MCInst1_MC2_v3_1Inst_0_U3  ( .A(MCInst1_MC2_v3_0 [3]), .B(
        MCInst1_MC2_v3_2 [2]), .Z(MCInst1_MC2_v3_1 [0]) );
  XOR2_X1 MCInst1_MC2_v3_2Inst_0_U3  ( .A(MCInst1_MC2_v3_2 [3]), .B(
        MCInst1_MC2_v3_0 [2]), .Z(MCInst1_MC2_v3_2 [0]) );
  XNOR2_X1 MCInst1_MC2_v3_3Inst_0_U4  ( .A(MCInst1_MC2_v3_3Inst_0_n2 ), .B(
        MCInst1_MC2_v3_0 [2]), .ZN(MCInst1_MC2_v3_3 [0]) );
  XNOR2_X1 MCInst1_MC2_v3_3Inst_0_U3  ( .A(MCInst1_MC2_v3_2 [2]), .B(
        MCInst1_MC2_v3_2 [3]), .ZN(MCInst1_MC2_v3_3Inst_0_n2 ) );
  XOR2_X1 MCInst1_MC2_v0_0Inst_1_U3  ( .A(MCInst1_MC2_v0_3 [3]), .B(
        MCInst1_MC2_v0_3 [0]), .Z(MCInst1_MC2_v0_0 [1]) );
  XOR2_X1 MCInst1_MC2_v0_1Inst_1_U3  ( .A(MCInst1_MC2_v0_0 [3]), .B(
        MCInst1_MC2_v0_3 [3]), .Z(MCInst1_MC2_v0_1 [1]) );
  XNOR2_X1 MCInst1_MC2_v0_2Inst_1_U4  ( .A(MCInst1_MC2_v0_2Inst_1_n2 ), .B(
        MCInst1_MC2_v0_3 [3]), .ZN(MCInst1_MC2_v0_2 [1]) );
  XNOR2_X1 MCInst1_MC2_v0_2Inst_1_U3  ( .A(MCInst1_MC2_v0_3 [0]), .B(
        ShiftRowsOutput[52]), .ZN(MCInst1_MC2_v0_2Inst_1_n2 ) );
  XOR2_X1 MCInst1_MC2_v0_3Inst_1_U3  ( .A(ShiftRowsOutput[52]), .B(
        MCInst1_MC2_v0_3 [0]), .Z(MCInst1_MC2_v0_3 [1]) );
  XOR2_X1 MCInst1_MC2_v1_1Inst_1_U3  ( .A(ShiftRowsOutput[36]), .B(
        MCInst1_MC2_v1_3 [3]), .Z(MCInst1_MC2_v1_1 [1]) );
  XOR2_X1 MCInst1_MC2_v1_2Inst_1_U3  ( .A(ShiftRowsOutput[36]), .B(
        MCInst1_MC2_v1_3 [2]), .Z(MCInst1_MC2_v1_2 [1]) );
  XOR2_X1 MCInst1_MC2_v1_3Inst_1_U3  ( .A(ShiftRowsOutput[36]), .B(
        MCInst1_MC2_v1_3 [0]), .Z(MCInst1_MC2_v1_3 [1]) );
  XOR2_X1 MCInst1_MC2_v2_0Inst_1_U3  ( .A(MCInst1_MC2_v2_3 [1]), .B(
        MCInst1_MC2_v2_0 [0]), .Z(MCInst1_MC2_v2_0 [1]) );
  XNOR2_X1 MCInst1_MC2_v2_1Inst_1_U4  ( .A(MCInst1_MC2_v2_1Inst_1_n2 ), .B(
        MCInst1_MC2_v2_0 [3]), .ZN(MCInst1_MC2_v2_1 [1]) );
  XNOR2_X1 MCInst1_MC2_v2_1Inst_1_U3  ( .A(MCInst1_MC2_v2_0 [0]), .B(
        MCInst1_MC2_v2_0 [2]), .ZN(MCInst1_MC2_v2_1Inst_1_n2 ) );
  XNOR2_X1 MCInst1_MC2_v2_2Inst_1_U5  ( .A(MCInst1_MC2_v2_2Inst_1_n4 ), .B(
        MCInst1_MC2_v2_2Inst_1_n3 ), .ZN(MCInst1_MC2_v2_2 [1]) );
  XNOR2_X1 MCInst1_MC2_v2_2Inst_1_U4  ( .A(MCInst1_MC2_v2_0 [2]), .B(
        MCInst1_MC2_v2_3 [1]), .ZN(MCInst1_MC2_v2_2Inst_1_n3 ) );
  XOR2_X1 MCInst1_MC2_v2_2Inst_1_U3  ( .A(MCInst1_MC2_v2_0 [3]), .B(
        MCInst1_MC2_v2_0 [0]), .Z(MCInst1_MC2_v2_2Inst_1_n4 ) );
  XOR2_X1 MCInst1_MC2_v3_0Inst_1_U3  ( .A(MCInst1_MC2_v3_2 [3]), .B(
        MCInst1_MC2_v3_2 [2]), .Z(MCInst1_MC2_v3_0 [1]) );
  XOR2_X1 MCInst1_MC2_v3_1Inst_1_U3  ( .A(MCInst1_MC2_v3_2 [3]), .B(
        MCInst1_MC2_v3_0 [3]), .Z(MCInst1_MC2_v3_1 [1]) );
  XNOR2_X1 MCInst1_MC2_v3_3Inst_1_U4  ( .A(MCInst1_MC2_v3_3Inst_1_n2 ), .B(
        MCInst1_MC2_v3_0 [3]), .ZN(MCInst1_MC2_v3_3 [1]) );
  XNOR2_X1 MCInst1_MC2_v3_3Inst_1_U3  ( .A(MCInst1_MC2_v3_2 [2]), .B(
        MCInst1_MC2_v3_2 [3]), .ZN(MCInst1_MC2_v3_3Inst_1_n2 ) );
  XOR2_X1 MCInst1_MC2_v0_0Inst_2_U3  ( .A(ShiftRowsOutput[52]), .B(
        MCInst1_MC2_v0_3 [0]), .Z(MCInst1_MC2_v0_0 [2]) );
  XOR2_X1 MCInst1_MC2_v0_1Inst_2_U3  ( .A(MCInst1_MC2_v0_3 [3]), .B(
        MCInst1_MC2_v0_3 [0]), .Z(MCInst1_MC2_v0_1 [2]) );
  XOR2_X1 MCInst1_MC2_v0_2Inst_2_U3  ( .A(MCInst1_MC2_v0_0 [3]), .B(
        MCInst1_MC2_v0_3 [0]), .Z(MCInst1_MC2_v0_2 [2]) );
  XNOR2_X1 MCInst1_MC2_v1_1Inst_2_U4  ( .A(MCInst1_MC2_v1_1Inst_2_n2 ), .B(
        MCInst1_MC2_v1_3 [2]), .ZN(MCInst1_MC2_v1_1 [2]) );
  XNOR2_X1 MCInst1_MC2_v1_1Inst_2_U3  ( .A(MCInst1_MC2_v1_3 [0]), .B(
        ShiftRowsOutput[36]), .ZN(MCInst1_MC2_v1_1Inst_2_n2 ) );
  XNOR2_X1 MCInst1_MC2_v1_2Inst_2_U4  ( .A(MCInst1_MC2_v1_2Inst_2_n2 ), .B(
        MCInst1_MC2_v1_3 [2]), .ZN(MCInst1_MC2_v1_2 [2]) );
  XNOR2_X1 MCInst1_MC2_v1_2Inst_2_U3  ( .A(MCInst1_MC2_v1_3 [3]), .B(
        ShiftRowsOutput[36]), .ZN(MCInst1_MC2_v1_2Inst_2_n2 ) );
  XNOR2_X1 MCInst1_MC2_v2_1Inst_2_U4  ( .A(MCInst1_MC2_v2_1Inst_2_n2 ), .B(
        MCInst1_MC2_v2_0 [3]), .ZN(MCInst1_MC2_v2_1 [2]) );
  XNOR2_X1 MCInst1_MC2_v2_1Inst_2_U3  ( .A(MCInst1_MC2_v2_0 [0]), .B(
        MCInst1_MC2_v2_3 [1]), .ZN(MCInst1_MC2_v2_1Inst_2_n2 ) );
  XNOR2_X1 MCInst1_MC2_v2_2Inst_2_U4  ( .A(MCInst1_MC2_v2_2Inst_2_n2 ), .B(
        MCInst1_MC2_v2_0 [3]), .ZN(MCInst1_MC2_v2_2 [2]) );
  XNOR2_X1 MCInst1_MC2_v2_2Inst_2_U3  ( .A(MCInst1_MC2_v2_0 [0]), .B(
        MCInst1_MC2_v2_0 [2]), .ZN(MCInst1_MC2_v2_2Inst_2_n2 ) );
  XOR2_X1 MCInst1_MC2_v2_3Inst_2_U3  ( .A(MCInst1_MC2_v2_3 [1]), .B(
        MCInst1_MC2_v2_0 [2]), .Z(MCInst1_MC2_v2_3 [2]) );
  XNOR2_X1 MCInst1_MC2_v3_1Inst_2_U4  ( .A(MCInst1_MC2_v3_1Inst_2_n2 ), .B(
        MCInst1_MC2_v3_0 [2]), .ZN(MCInst1_MC2_v3_1 [2]) );
  XNOR2_X1 MCInst1_MC2_v3_1Inst_2_U3  ( .A(MCInst1_MC2_v3_2 [2]), .B(
        MCInst1_MC2_v3_2 [3]), .ZN(MCInst1_MC2_v3_1Inst_2_n2 ) );
  XOR2_X1 MCInst1_MC2_v3_3Inst_2_U3  ( .A(MCInst1_MC2_v3_0 [2]), .B(
        MCInst1_MC2_v3_2 [2]), .Z(MCInst1_MC2_v3_3 [2]) );
  XOR2_X1 MCInst1_MC2_v0_1Inst_3_U3  ( .A(ShiftRowsOutput[52]), .B(
        MCInst1_MC2_v0_3 [0]), .Z(MCInst1_MC2_v0_1 [3]) );
  XOR2_X1 MCInst1_MC2_v0_2Inst_3_U3  ( .A(ShiftRowsOutput[52]), .B(
        MCInst1_MC2_v0_3 [3]), .Z(MCInst1_MC2_v0_2 [3]) );
  XOR2_X1 MCInst1_MC2_v1_1Inst_3_U3  ( .A(MCInst1_MC2_v1_3 [2]), .B(
        MCInst1_MC2_v1_3 [3]), .Z(MCInst1_MC2_v1_1 [3]) );
  XNOR2_X1 MCInst1_MC2_v1_2Inst_3_U5  ( .A(MCInst1_MC2_v1_2Inst_3_n4 ), .B(
        MCInst1_MC2_v1_2Inst_3_n3 ), .ZN(MCInst1_MC2_v1_2 [3]) );
  XNOR2_X1 MCInst1_MC2_v1_2Inst_3_U4  ( .A(MCInst1_MC2_v1_3 [2]), .B(
        ShiftRowsOutput[36]), .ZN(MCInst1_MC2_v1_2Inst_3_n3 ) );
  XOR2_X1 MCInst1_MC2_v1_2Inst_3_U3  ( .A(MCInst1_MC2_v1_3 [3]), .B(
        MCInst1_MC2_v1_3 [0]), .Z(MCInst1_MC2_v1_2Inst_3_n4 ) );
  XOR2_X1 MCInst1_MC2_v2_1Inst_3_U3  ( .A(MCInst1_MC2_v2_0 [2]), .B(
        MCInst1_MC2_v2_0 [0]), .Z(MCInst1_MC2_v2_1 [3]) );
  XNOR2_X1 MCInst1_MC2_v2_2Inst_3_U4  ( .A(MCInst1_MC2_v2_2Inst_3_n2 ), .B(
        MCInst1_MC2_v2_0 [3]), .ZN(MCInst1_MC2_v2_2 [3]) );
  XNOR2_X1 MCInst1_MC2_v2_2Inst_3_U3  ( .A(MCInst1_MC2_v2_0 [0]), .B(
        MCInst1_MC2_v2_3 [1]), .ZN(MCInst1_MC2_v2_2Inst_3_n2 ) );
  XNOR2_X1 MCInst1_MC2_v2_3Inst_3_U4  ( .A(MCInst1_MC2_v2_3Inst_3_n2 ), .B(
        MCInst1_MC2_v2_0 [2]), .ZN(MCInst1_MC2_v2_3 [3]) );
  XNOR2_X1 MCInst1_MC2_v2_3Inst_3_U3  ( .A(MCInst1_MC2_v2_0 [3]), .B(
        MCInst1_MC2_v2_3 [1]), .ZN(MCInst1_MC2_v2_3Inst_3_n2 ) );
  XOR2_X1 MCInst1_MC2_v3_1Inst_3_U3  ( .A(MCInst1_MC2_v3_0 [2]), .B(
        MCInst1_MC2_v3_0 [3]), .Z(MCInst1_MC2_v3_1 [3]) );
  XOR2_X1 MCInst1_MC2_v3_3Inst_3_U3  ( .A(MCInst1_MC2_v3_2 [3]), .B(
        MCInst1_MC2_v3_0 [3]), .Z(MCInst1_MC2_v3_3 [3]) );
  XNOR2_X1 MCInst1_MC2_r0Inst_XORInst_0_0_U3  ( .A(
        MCInst1_MC2_r0Inst_XORInst_0_0_n5 ), .B(
        MCInst1_MC2_r0Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[52]) );
  XNOR2_X1 MCInst1_MC2_r0Inst_XORInst_0_0_U2  ( .A(MCInst1_MC2_v3_2 [2]), 
        .B(MCInst1_MC2_v2_0 [0]), .ZN(MCInst1_MC2_r0Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst1_MC2_r0Inst_XORInst_0_0_U1  ( .A(MCInst1_MC2_v0_3 [3]), .B(
        ShiftRowsOutput[36]), .Z(MCInst1_MC2_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst1_MC2_r0Inst_XORInst_0_1_U3  ( .A(
        MCInst1_MC2_r0Inst_XORInst_0_1_n5 ), .B(
        MCInst1_MC2_r0Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[53]) );
  XNOR2_X1 MCInst1_MC2_r0Inst_XORInst_0_1_U2  ( .A(MCInst1_MC2_v3_0 [1]), 
        .B(MCInst1_MC2_v2_0 [1]), .ZN(MCInst1_MC2_r0Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst1_MC2_r0Inst_XORInst_0_1_U1  ( .A(MCInst1_MC2_v0_0 [1]), .B(
        MCInst1_MC2_v1_3 [2]), .Z(MCInst1_MC2_r0Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst1_MC2_r0Inst_XORInst_0_2_U3  ( .A(
        MCInst1_MC2_r0Inst_XORInst_0_2_n5 ), .B(
        MCInst1_MC2_r0Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[54]) );
  XNOR2_X1 MCInst1_MC2_r0Inst_XORInst_0_2_U2  ( .A(MCInst1_MC2_v3_0 [2]), 
        .B(MCInst1_MC2_v2_0 [2]), .ZN(MCInst1_MC2_r0Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst1_MC2_r0Inst_XORInst_0_2_U1  ( .A(MCInst1_MC2_v0_0 [2]), .B(
        MCInst1_MC2_v1_3 [3]), .Z(MCInst1_MC2_r0Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst1_MC2_r0Inst_XORInst_0_3_U3  ( .A(
        MCInst1_MC2_r0Inst_XORInst_0_3_n5 ), .B(
        MCInst1_MC2_r0Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[55]) );
  XNOR2_X1 MCInst1_MC2_r0Inst_XORInst_0_3_U2  ( .A(MCInst1_MC2_v3_0 [3]), 
        .B(MCInst1_MC2_v2_0 [3]), .ZN(MCInst1_MC2_r0Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst1_MC2_r0Inst_XORInst_0_3_U1  ( .A(MCInst1_MC2_v0_0 [3]), .B(
        MCInst1_MC2_v1_3 [0]), .Z(MCInst1_MC2_r0Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst1_MC2_r1Inst_XORInst_0_0_U3  ( .A(
        MCInst1_MC2_r1Inst_XORInst_0_0_n5 ), .B(
        MCInst1_MC2_r1Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[36]) );
  XNOR2_X1 MCInst1_MC2_r1Inst_XORInst_0_0_U2  ( .A(MCInst1_MC2_v3_1 [0]), 
        .B(MCInst1_MC2_v2_1 [0]), .ZN(MCInst1_MC2_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst1_MC2_r1Inst_XORInst_0_0_U1  ( .A(MCInst1_MC2_v0_0 [3]), .B(
        MCInst1_MC2_v1_1 [0]), .Z(MCInst1_MC2_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst1_MC2_r1Inst_XORInst_0_1_U3  ( .A(
        MCInst1_MC2_r1Inst_XORInst_0_1_n5 ), .B(
        MCInst1_MC2_r1Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[37]) );
  XNOR2_X1 MCInst1_MC2_r1Inst_XORInst_0_1_U2  ( .A(MCInst1_MC2_v3_1 [1]), 
        .B(MCInst1_MC2_v2_1 [1]), .ZN(MCInst1_MC2_r1Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst1_MC2_r1Inst_XORInst_0_1_U1  ( .A(MCInst1_MC2_v0_1 [1]), .B(
        MCInst1_MC2_v1_1 [1]), .Z(MCInst1_MC2_r1Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst1_MC2_r1Inst_XORInst_0_2_U3  ( .A(
        MCInst1_MC2_r1Inst_XORInst_0_2_n5 ), .B(
        MCInst1_MC2_r1Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[38]) );
  XNOR2_X1 MCInst1_MC2_r1Inst_XORInst_0_2_U2  ( .A(MCInst1_MC2_v3_1 [2]), 
        .B(MCInst1_MC2_v2_1 [2]), .ZN(MCInst1_MC2_r1Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst1_MC2_r1Inst_XORInst_0_2_U1  ( .A(MCInst1_MC2_v0_1 [2]), .B(
        MCInst1_MC2_v1_1 [2]), .Z(MCInst1_MC2_r1Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst1_MC2_r1Inst_XORInst_0_3_U3  ( .A(
        MCInst1_MC2_r1Inst_XORInst_0_3_n5 ), .B(
        MCInst1_MC2_r1Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[39]) );
  XNOR2_X1 MCInst1_MC2_r1Inst_XORInst_0_3_U2  ( .A(MCInst1_MC2_v3_1 [3]), 
        .B(MCInst1_MC2_v2_1 [3]), .ZN(MCInst1_MC2_r1Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst1_MC2_r1Inst_XORInst_0_3_U1  ( .A(MCInst1_MC2_v0_1 [3]), .B(
        MCInst1_MC2_v1_1 [3]), .Z(MCInst1_MC2_r1Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst1_MC2_r2Inst_XORInst_0_0_U3  ( .A(
        MCInst1_MC2_r2Inst_XORInst_0_0_n5 ), .B(
        MCInst1_MC2_r2Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[20]) );
  XNOR2_X1 MCInst1_MC2_r2Inst_XORInst_0_0_U2  ( .A(MCInst1_MC2_v3_2 [0]), 
        .B(MCInst1_MC2_v2_2 [0]), .ZN(MCInst1_MC2_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst1_MC2_r2Inst_XORInst_0_0_U1  ( .A(MCInst1_MC2_v0_2 [0]), .B(
        MCInst1_MC2_v1_2 [0]), .Z(MCInst1_MC2_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst1_MC2_r2Inst_XORInst_0_1_U3  ( .A(
        MCInst1_MC2_r2Inst_XORInst_0_1_n5 ), .B(
        MCInst1_MC2_r2Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[21]) );
  XNOR2_X1 MCInst1_MC2_r2Inst_XORInst_0_1_U2  ( .A(MCInst1_MC2_v3_0 [3]), 
        .B(MCInst1_MC2_v2_2 [1]), .ZN(MCInst1_MC2_r2Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst1_MC2_r2Inst_XORInst_0_1_U1  ( .A(MCInst1_MC2_v0_2 [1]), .B(
        MCInst1_MC2_v1_2 [1]), .Z(MCInst1_MC2_r2Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst1_MC2_r2Inst_XORInst_0_2_U3  ( .A(
        MCInst1_MC2_r2Inst_XORInst_0_2_n5 ), .B(
        MCInst1_MC2_r2Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[22]) );
  XNOR2_X1 MCInst1_MC2_r2Inst_XORInst_0_2_U2  ( .A(MCInst1_MC2_v3_2 [2]), 
        .B(MCInst1_MC2_v2_2 [2]), .ZN(MCInst1_MC2_r2Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst1_MC2_r2Inst_XORInst_0_2_U1  ( .A(MCInst1_MC2_v0_2 [2]), .B(
        MCInst1_MC2_v1_2 [2]), .Z(MCInst1_MC2_r2Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst1_MC2_r2Inst_XORInst_0_3_U3  ( .A(
        MCInst1_MC2_r2Inst_XORInst_0_3_n5 ), .B(
        MCInst1_MC2_r2Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[23]) );
  XNOR2_X1 MCInst1_MC2_r2Inst_XORInst_0_3_U2  ( .A(MCInst1_MC2_v3_2 [3]), 
        .B(MCInst1_MC2_v2_2 [3]), .ZN(MCInst1_MC2_r2Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst1_MC2_r2Inst_XORInst_0_3_U1  ( .A(MCInst1_MC2_v0_2 [3]), .B(
        MCInst1_MC2_v1_2 [3]), .Z(MCInst1_MC2_r2Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst1_MC2_r3Inst_XORInst_0_0_U3  ( .A(
        MCInst1_MC2_r3Inst_XORInst_0_0_n5 ), .B(
        MCInst1_MC2_r3Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[4]) );
  XNOR2_X1 MCInst1_MC2_r3Inst_XORInst_0_0_U2  ( .A(MCInst1_MC2_v3_3 [0]), 
        .B(MCInst1_MC2_v2_3 [0]), .ZN(MCInst1_MC2_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst1_MC2_r3Inst_XORInst_0_0_U1  ( .A(MCInst1_MC2_v0_3 [0]), .B(
        MCInst1_MC2_v1_3 [0]), .Z(MCInst1_MC2_r3Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst1_MC2_r3Inst_XORInst_0_1_U3  ( .A(
        MCInst1_MC2_r3Inst_XORInst_0_1_n5 ), .B(
        MCInst1_MC2_r3Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[5]) );
  XNOR2_X1 MCInst1_MC2_r3Inst_XORInst_0_1_U2  ( .A(MCInst1_MC2_v3_3 [1]), 
        .B(MCInst1_MC2_v2_3 [1]), .ZN(MCInst1_MC2_r3Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst1_MC2_r3Inst_XORInst_0_1_U1  ( .A(MCInst1_MC2_v0_3 [1]), .B(
        MCInst1_MC2_v1_3 [1]), .Z(MCInst1_MC2_r3Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst1_MC2_r3Inst_XORInst_0_2_U3  ( .A(
        MCInst1_MC2_r3Inst_XORInst_0_2_n5 ), .B(
        MCInst1_MC2_r3Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[6]) );
  XNOR2_X1 MCInst1_MC2_r3Inst_XORInst_0_2_U2  ( .A(MCInst1_MC2_v3_3 [2]), 
        .B(MCInst1_MC2_v2_3 [2]), .ZN(MCInst1_MC2_r3Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst1_MC2_r3Inst_XORInst_0_2_U1  ( .A(MCInst1_MC2_v0_0 [3]), .B(
        MCInst1_MC2_v1_3 [2]), .Z(MCInst1_MC2_r3Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst1_MC2_r3Inst_XORInst_0_3_U3  ( .A(
        MCInst1_MC2_r3Inst_XORInst_0_3_n5 ), .B(
        MCInst1_MC2_r3Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[7]) );
  XNOR2_X1 MCInst1_MC2_r3Inst_XORInst_0_3_U2  ( .A(MCInst1_MC2_v3_3 [3]), 
        .B(MCInst1_MC2_v2_3 [3]), .ZN(MCInst1_MC2_r3Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst1_MC2_r3Inst_XORInst_0_3_U1  ( .A(MCInst1_MC2_v0_3 [3]), .B(
        MCInst1_MC2_v1_3 [3]), .Z(MCInst1_MC2_r3Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst1_MC3_v0_2Inst_0_U4  ( .A(MCInst1_MC3_v0_2Inst_0_n2 ), .B(
        MCInst1_MC3_v0_0 [3]), .ZN(MCInst1_MC3_v0_2 [0]) );
  XNOR2_X1 MCInst1_MC3_v0_2Inst_0_U3  ( .A(MCInst1_MC3_v0_3 [0]), .B(
        ShiftRowsOutput[48]), .ZN(MCInst1_MC3_v0_2Inst_0_n2 ) );
  XOR2_X1 MCInst1_MC3_v1_1Inst_0_U3  ( .A(MCInst1_MC3_v1_3 [3]), .B(
        MCInst1_MC3_v1_3 [0]), .Z(MCInst1_MC3_v1_1 [0]) );
  XNOR2_X1 MCInst1_MC3_v1_2Inst_0_U4  ( .A(MCInst1_MC3_v1_2Inst_0_n2 ), .B(
        MCInst1_MC3_v1_3 [3]), .ZN(MCInst1_MC3_v1_2 [0]) );
  XNOR2_X1 MCInst1_MC3_v1_2Inst_0_U3  ( .A(MCInst1_MC3_v1_3 [0]), .B(
        MCInst1_MC3_v1_3 [2]), .ZN(MCInst1_MC3_v1_2Inst_0_n2 ) );
  XOR2_X1 MCInst1_MC3_v2_1Inst_0_U3  ( .A(MCInst1_MC3_v2_3 [1]), .B(
        MCInst1_MC3_v2_0 [3]), .Z(MCInst1_MC3_v2_1 [0]) );
  XOR2_X1 MCInst1_MC3_v2_2Inst_0_U3  ( .A(MCInst1_MC3_v2_0 [2]), .B(
        MCInst1_MC3_v2_0 [0]), .Z(MCInst1_MC3_v2_2 [0]) );
  XNOR2_X1 MCInst1_MC3_v2_3Inst_0_U5  ( .A(MCInst1_MC3_v2_3Inst_0_n4 ), .B(
        MCInst1_MC3_v2_3Inst_0_n3 ), .ZN(MCInst1_MC3_v2_3 [0]) );
  XNOR2_X1 MCInst1_MC3_v2_3Inst_0_U4  ( .A(MCInst1_MC3_v2_0 [2]), .B(
        MCInst1_MC3_v2_3 [1]), .ZN(MCInst1_MC3_v2_3Inst_0_n3 ) );
  XOR2_X1 MCInst1_MC3_v2_3Inst_0_U3  ( .A(MCInst1_MC3_v2_0 [3]), .B(
        MCInst1_MC3_v2_0 [0]), .Z(MCInst1_MC3_v2_3Inst_0_n4 ) );
  XOR2_X1 MCInst1_MC3_v3_1Inst_0_U3  ( .A(MCInst1_MC3_v3_0 [3]), .B(
        MCInst1_MC3_v3_2 [2]), .Z(MCInst1_MC3_v3_1 [0]) );
  XOR2_X1 MCInst1_MC3_v3_2Inst_0_U3  ( .A(MCInst1_MC3_v3_2 [3]), .B(
        MCInst1_MC3_v3_0 [2]), .Z(MCInst1_MC3_v3_2 [0]) );
  XNOR2_X1 MCInst1_MC3_v3_3Inst_0_U4  ( .A(MCInst1_MC3_v3_3Inst_0_n2 ), .B(
        MCInst1_MC3_v3_0 [2]), .ZN(MCInst1_MC3_v3_3 [0]) );
  XNOR2_X1 MCInst1_MC3_v3_3Inst_0_U3  ( .A(MCInst1_MC3_v3_2 [2]), .B(
        MCInst1_MC3_v3_2 [3]), .ZN(MCInst1_MC3_v3_3Inst_0_n2 ) );
  XOR2_X1 MCInst1_MC3_v0_0Inst_1_U3  ( .A(MCInst1_MC3_v0_3 [3]), .B(
        MCInst1_MC3_v0_3 [0]), .Z(MCInst1_MC3_v0_0 [1]) );
  XOR2_X1 MCInst1_MC3_v0_1Inst_1_U3  ( .A(MCInst1_MC3_v0_0 [3]), .B(
        MCInst1_MC3_v0_3 [3]), .Z(MCInst1_MC3_v0_1 [1]) );
  XNOR2_X1 MCInst1_MC3_v0_2Inst_1_U4  ( .A(MCInst1_MC3_v0_2Inst_1_n2 ), .B(
        MCInst1_MC3_v0_3 [3]), .ZN(MCInst1_MC3_v0_2 [1]) );
  XNOR2_X1 MCInst1_MC3_v0_2Inst_1_U3  ( .A(MCInst1_MC3_v0_3 [0]), .B(
        ShiftRowsOutput[48]), .ZN(MCInst1_MC3_v0_2Inst_1_n2 ) );
  XOR2_X1 MCInst1_MC3_v0_3Inst_1_U3  ( .A(ShiftRowsOutput[48]), .B(
        MCInst1_MC3_v0_3 [0]), .Z(MCInst1_MC3_v0_3 [1]) );
  XOR2_X1 MCInst1_MC3_v1_1Inst_1_U3  ( .A(ShiftRowsOutput[32]), .B(
        MCInst1_MC3_v1_3 [3]), .Z(MCInst1_MC3_v1_1 [1]) );
  XOR2_X1 MCInst1_MC3_v1_2Inst_1_U3  ( .A(ShiftRowsOutput[32]), .B(
        MCInst1_MC3_v1_3 [2]), .Z(MCInst1_MC3_v1_2 [1]) );
  XOR2_X1 MCInst1_MC3_v1_3Inst_1_U3  ( .A(ShiftRowsOutput[32]), .B(
        MCInst1_MC3_v1_3 [0]), .Z(MCInst1_MC3_v1_3 [1]) );
  XOR2_X1 MCInst1_MC3_v2_0Inst_1_U3  ( .A(MCInst1_MC3_v2_3 [1]), .B(
        MCInst1_MC3_v2_0 [0]), .Z(MCInst1_MC3_v2_0 [1]) );
  XNOR2_X1 MCInst1_MC3_v2_1Inst_1_U4  ( .A(MCInst1_MC3_v2_1Inst_1_n2 ), .B(
        MCInst1_MC3_v2_0 [3]), .ZN(MCInst1_MC3_v2_1 [1]) );
  XNOR2_X1 MCInst1_MC3_v2_1Inst_1_U3  ( .A(MCInst1_MC3_v2_0 [0]), .B(
        MCInst1_MC3_v2_0 [2]), .ZN(MCInst1_MC3_v2_1Inst_1_n2 ) );
  XNOR2_X1 MCInst1_MC3_v2_2Inst_1_U5  ( .A(MCInst1_MC3_v2_2Inst_1_n4 ), .B(
        MCInst1_MC3_v2_2Inst_1_n3 ), .ZN(MCInst1_MC3_v2_2 [1]) );
  XNOR2_X1 MCInst1_MC3_v2_2Inst_1_U4  ( .A(MCInst1_MC3_v2_0 [2]), .B(
        MCInst1_MC3_v2_3 [1]), .ZN(MCInst1_MC3_v2_2Inst_1_n3 ) );
  XOR2_X1 MCInst1_MC3_v2_2Inst_1_U3  ( .A(MCInst1_MC3_v2_0 [3]), .B(
        MCInst1_MC3_v2_0 [0]), .Z(MCInst1_MC3_v2_2Inst_1_n4 ) );
  XOR2_X1 MCInst1_MC3_v3_0Inst_1_U3  ( .A(MCInst1_MC3_v3_2 [3]), .B(
        MCInst1_MC3_v3_2 [2]), .Z(MCInst1_MC3_v3_0 [1]) );
  XOR2_X1 MCInst1_MC3_v3_1Inst_1_U3  ( .A(MCInst1_MC3_v3_2 [3]), .B(
        MCInst1_MC3_v3_0 [3]), .Z(MCInst1_MC3_v3_1 [1]) );
  XNOR2_X1 MCInst1_MC3_v3_3Inst_1_U4  ( .A(MCInst1_MC3_v3_3Inst_1_n2 ), .B(
        MCInst1_MC3_v3_0 [3]), .ZN(MCInst1_MC3_v3_3 [1]) );
  XNOR2_X1 MCInst1_MC3_v3_3Inst_1_U3  ( .A(MCInst1_MC3_v3_2 [2]), .B(
        MCInst1_MC3_v3_2 [3]), .ZN(MCInst1_MC3_v3_3Inst_1_n2 ) );
  XOR2_X1 MCInst1_MC3_v0_0Inst_2_U3  ( .A(ShiftRowsOutput[48]), .B(
        MCInst1_MC3_v0_3 [0]), .Z(MCInst1_MC3_v0_0 [2]) );
  XOR2_X1 MCInst1_MC3_v0_1Inst_2_U3  ( .A(MCInst1_MC3_v0_3 [3]), .B(
        MCInst1_MC3_v0_3 [0]), .Z(MCInst1_MC3_v0_1 [2]) );
  XOR2_X1 MCInst1_MC3_v0_2Inst_2_U3  ( .A(MCInst1_MC3_v0_0 [3]), .B(
        MCInst1_MC3_v0_3 [0]), .Z(MCInst1_MC3_v0_2 [2]) );
  XNOR2_X1 MCInst1_MC3_v1_1Inst_2_U4  ( .A(MCInst1_MC3_v1_1Inst_2_n2 ), .B(
        MCInst1_MC3_v1_3 [2]), .ZN(MCInst1_MC3_v1_1 [2]) );
  XNOR2_X1 MCInst1_MC3_v1_1Inst_2_U3  ( .A(MCInst1_MC3_v1_3 [0]), .B(
        ShiftRowsOutput[32]), .ZN(MCInst1_MC3_v1_1Inst_2_n2 ) );
  XNOR2_X1 MCInst1_MC3_v1_2Inst_2_U4  ( .A(MCInst1_MC3_v1_2Inst_2_n2 ), .B(
        MCInst1_MC3_v1_3 [2]), .ZN(MCInst1_MC3_v1_2 [2]) );
  XNOR2_X1 MCInst1_MC3_v1_2Inst_2_U3  ( .A(MCInst1_MC3_v1_3 [3]), .B(
        ShiftRowsOutput[32]), .ZN(MCInst1_MC3_v1_2Inst_2_n2 ) );
  XNOR2_X1 MCInst1_MC3_v2_1Inst_2_U4  ( .A(MCInst1_MC3_v2_1Inst_2_n2 ), .B(
        MCInst1_MC3_v2_0 [3]), .ZN(MCInst1_MC3_v2_1 [2]) );
  XNOR2_X1 MCInst1_MC3_v2_1Inst_2_U3  ( .A(MCInst1_MC3_v2_0 [0]), .B(
        MCInst1_MC3_v2_3 [1]), .ZN(MCInst1_MC3_v2_1Inst_2_n2 ) );
  XNOR2_X1 MCInst1_MC3_v2_2Inst_2_U4  ( .A(MCInst1_MC3_v2_2Inst_2_n2 ), .B(
        MCInst1_MC3_v2_0 [3]), .ZN(MCInst1_MC3_v2_2 [2]) );
  XNOR2_X1 MCInst1_MC3_v2_2Inst_2_U3  ( .A(MCInst1_MC3_v2_0 [0]), .B(
        MCInst1_MC3_v2_0 [2]), .ZN(MCInst1_MC3_v2_2Inst_2_n2 ) );
  XOR2_X1 MCInst1_MC3_v2_3Inst_2_U3  ( .A(MCInst1_MC3_v2_3 [1]), .B(
        MCInst1_MC3_v2_0 [2]), .Z(MCInst1_MC3_v2_3 [2]) );
  XNOR2_X1 MCInst1_MC3_v3_1Inst_2_U4  ( .A(MCInst1_MC3_v3_1Inst_2_n2 ), .B(
        MCInst1_MC3_v3_0 [2]), .ZN(MCInst1_MC3_v3_1 [2]) );
  XNOR2_X1 MCInst1_MC3_v3_1Inst_2_U3  ( .A(MCInst1_MC3_v3_2 [2]), .B(
        MCInst1_MC3_v3_2 [3]), .ZN(MCInst1_MC3_v3_1Inst_2_n2 ) );
  XOR2_X1 MCInst1_MC3_v3_3Inst_2_U3  ( .A(MCInst1_MC3_v3_0 [2]), .B(
        MCInst1_MC3_v3_2 [2]), .Z(MCInst1_MC3_v3_3 [2]) );
  XOR2_X1 MCInst1_MC3_v0_1Inst_3_U3  ( .A(ShiftRowsOutput[48]), .B(
        MCInst1_MC3_v0_3 [0]), .Z(MCInst1_MC3_v0_1 [3]) );
  XOR2_X1 MCInst1_MC3_v0_2Inst_3_U3  ( .A(ShiftRowsOutput[48]), .B(
        MCInst1_MC3_v0_3 [3]), .Z(MCInst1_MC3_v0_2 [3]) );
  XOR2_X1 MCInst1_MC3_v1_1Inst_3_U3  ( .A(MCInst1_MC3_v1_3 [2]), .B(
        MCInst1_MC3_v1_3 [3]), .Z(MCInst1_MC3_v1_1 [3]) );
  XNOR2_X1 MCInst1_MC3_v1_2Inst_3_U5  ( .A(MCInst1_MC3_v1_2Inst_3_n4 ), .B(
        MCInst1_MC3_v1_2Inst_3_n3 ), .ZN(MCInst1_MC3_v1_2 [3]) );
  XNOR2_X1 MCInst1_MC3_v1_2Inst_3_U4  ( .A(MCInst1_MC3_v1_3 [2]), .B(
        ShiftRowsOutput[32]), .ZN(MCInst1_MC3_v1_2Inst_3_n3 ) );
  XOR2_X1 MCInst1_MC3_v1_2Inst_3_U3  ( .A(MCInst1_MC3_v1_3 [3]), .B(
        MCInst1_MC3_v1_3 [0]), .Z(MCInst1_MC3_v1_2Inst_3_n4 ) );
  XOR2_X1 MCInst1_MC3_v2_1Inst_3_U3  ( .A(MCInst1_MC3_v2_0 [2]), .B(
        MCInst1_MC3_v2_0 [0]), .Z(MCInst1_MC3_v2_1 [3]) );
  XNOR2_X1 MCInst1_MC3_v2_2Inst_3_U4  ( .A(MCInst1_MC3_v2_2Inst_3_n2 ), .B(
        MCInst1_MC3_v2_0 [3]), .ZN(MCInst1_MC3_v2_2 [3]) );
  XNOR2_X1 MCInst1_MC3_v2_2Inst_3_U3  ( .A(MCInst1_MC3_v2_0 [0]), .B(
        MCInst1_MC3_v2_3 [1]), .ZN(MCInst1_MC3_v2_2Inst_3_n2 ) );
  XNOR2_X1 MCInst1_MC3_v2_3Inst_3_U4  ( .A(MCInst1_MC3_v2_3Inst_3_n2 ), .B(
        MCInst1_MC3_v2_0 [2]), .ZN(MCInst1_MC3_v2_3 [3]) );
  XNOR2_X1 MCInst1_MC3_v2_3Inst_3_U3  ( .A(MCInst1_MC3_v2_0 [3]), .B(
        MCInst1_MC3_v2_3 [1]), .ZN(MCInst1_MC3_v2_3Inst_3_n2 ) );
  XOR2_X1 MCInst1_MC3_v3_1Inst_3_U3  ( .A(MCInst1_MC3_v3_0 [2]), .B(
        MCInst1_MC3_v3_0 [3]), .Z(MCInst1_MC3_v3_1 [3]) );
  XOR2_X1 MCInst1_MC3_v3_3Inst_3_U3  ( .A(MCInst1_MC3_v3_2 [3]), .B(
        MCInst1_MC3_v3_0 [3]), .Z(MCInst1_MC3_v3_3 [3]) );
  XNOR2_X1 MCInst1_MC3_r0Inst_XORInst_0_0_U3  ( .A(
        MCInst1_MC3_r0Inst_XORInst_0_0_n5 ), .B(
        MCInst1_MC3_r0Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[48]) );
  XNOR2_X1 MCInst1_MC3_r0Inst_XORInst_0_0_U2  ( .A(MCInst1_MC3_v3_2 [2]), 
        .B(MCInst1_MC3_v2_0 [0]), .ZN(MCInst1_MC3_r0Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst1_MC3_r0Inst_XORInst_0_0_U1  ( .A(MCInst1_MC3_v0_3 [3]), .B(
        ShiftRowsOutput[32]), .Z(MCInst1_MC3_r0Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst1_MC3_r0Inst_XORInst_0_1_U3  ( .A(
        MCInst1_MC3_r0Inst_XORInst_0_1_n5 ), .B(
        MCInst1_MC3_r0Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[49]) );
  XNOR2_X1 MCInst1_MC3_r0Inst_XORInst_0_1_U2  ( .A(MCInst1_MC3_v3_0 [1]), 
        .B(MCInst1_MC3_v2_0 [1]), .ZN(MCInst1_MC3_r0Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst1_MC3_r0Inst_XORInst_0_1_U1  ( .A(MCInst1_MC3_v0_0 [1]), .B(
        MCInst1_MC3_v1_3 [2]), .Z(MCInst1_MC3_r0Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst1_MC3_r0Inst_XORInst_0_2_U3  ( .A(
        MCInst1_MC3_r0Inst_XORInst_0_2_n5 ), .B(
        MCInst1_MC3_r0Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[50]) );
  XNOR2_X1 MCInst1_MC3_r0Inst_XORInst_0_2_U2  ( .A(MCInst1_MC3_v3_0 [2]), 
        .B(MCInst1_MC3_v2_0 [2]), .ZN(MCInst1_MC3_r0Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst1_MC3_r0Inst_XORInst_0_2_U1  ( .A(MCInst1_MC3_v0_0 [2]), .B(
        MCInst1_MC3_v1_3 [3]), .Z(MCInst1_MC3_r0Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst1_MC3_r0Inst_XORInst_0_3_U3  ( .A(
        MCInst1_MC3_r0Inst_XORInst_0_3_n5 ), .B(
        MCInst1_MC3_r0Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[51]) );
  XNOR2_X1 MCInst1_MC3_r0Inst_XORInst_0_3_U2  ( .A(MCInst1_MC3_v3_0 [3]), 
        .B(MCInst1_MC3_v2_0 [3]), .ZN(MCInst1_MC3_r0Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst1_MC3_r0Inst_XORInst_0_3_U1  ( .A(MCInst1_MC3_v0_0 [3]), .B(
        MCInst1_MC3_v1_3 [0]), .Z(MCInst1_MC3_r0Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst1_MC3_r1Inst_XORInst_0_0_U3  ( .A(
        MCInst1_MC3_r1Inst_XORInst_0_0_n5 ), .B(
        MCInst1_MC3_r1Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[32]) );
  XNOR2_X1 MCInst1_MC3_r1Inst_XORInst_0_0_U2  ( .A(MCInst1_MC3_v3_1 [0]), 
        .B(MCInst1_MC3_v2_1 [0]), .ZN(MCInst1_MC3_r1Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst1_MC3_r1Inst_XORInst_0_0_U1  ( .A(MCInst1_MC3_v0_0 [3]), .B(
        MCInst1_MC3_v1_1 [0]), .Z(MCInst1_MC3_r1Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst1_MC3_r1Inst_XORInst_0_1_U3  ( .A(
        MCInst1_MC3_r1Inst_XORInst_0_1_n5 ), .B(
        MCInst1_MC3_r1Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[33]) );
  XNOR2_X1 MCInst1_MC3_r1Inst_XORInst_0_1_U2  ( .A(MCInst1_MC3_v3_1 [1]), 
        .B(MCInst1_MC3_v2_1 [1]), .ZN(MCInst1_MC3_r1Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst1_MC3_r1Inst_XORInst_0_1_U1  ( .A(MCInst1_MC3_v0_1 [1]), .B(
        MCInst1_MC3_v1_1 [1]), .Z(MCInst1_MC3_r1Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst1_MC3_r1Inst_XORInst_0_2_U3  ( .A(
        MCInst1_MC3_r1Inst_XORInst_0_2_n5 ), .B(
        MCInst1_MC3_r1Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[34]) );
  XNOR2_X1 MCInst1_MC3_r1Inst_XORInst_0_2_U2  ( .A(MCInst1_MC3_v3_1 [2]), 
        .B(MCInst1_MC3_v2_1 [2]), .ZN(MCInst1_MC3_r1Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst1_MC3_r1Inst_XORInst_0_2_U1  ( .A(MCInst1_MC3_v0_1 [2]), .B(
        MCInst1_MC3_v1_1 [2]), .Z(MCInst1_MC3_r1Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst1_MC3_r1Inst_XORInst_0_3_U3  ( .A(
        MCInst1_MC3_r1Inst_XORInst_0_3_n5 ), .B(
        MCInst1_MC3_r1Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[35]) );
  XNOR2_X1 MCInst1_MC3_r1Inst_XORInst_0_3_U2  ( .A(MCInst1_MC3_v3_1 [3]), 
        .B(MCInst1_MC3_v2_1 [3]), .ZN(MCInst1_MC3_r1Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst1_MC3_r1Inst_XORInst_0_3_U1  ( .A(MCInst1_MC3_v0_1 [3]), .B(
        MCInst1_MC3_v1_1 [3]), .Z(MCInst1_MC3_r1Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst1_MC3_r2Inst_XORInst_0_0_U3  ( .A(
        MCInst1_MC3_r2Inst_XORInst_0_0_n5 ), .B(
        MCInst1_MC3_r2Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[16]) );
  XNOR2_X1 MCInst1_MC3_r2Inst_XORInst_0_0_U2  ( .A(MCInst1_MC3_v3_2 [0]), 
        .B(MCInst1_MC3_v2_2 [0]), .ZN(MCInst1_MC3_r2Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst1_MC3_r2Inst_XORInst_0_0_U1  ( .A(MCInst1_MC3_v0_2 [0]), .B(
        MCInst1_MC3_v1_2 [0]), .Z(MCInst1_MC3_r2Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst1_MC3_r2Inst_XORInst_0_1_U3  ( .A(
        MCInst1_MC3_r2Inst_XORInst_0_1_n5 ), .B(
        MCInst1_MC3_r2Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[17]) );
  XNOR2_X1 MCInst1_MC3_r2Inst_XORInst_0_1_U2  ( .A(MCInst1_MC3_v3_0 [3]), 
        .B(MCInst1_MC3_v2_2 [1]), .ZN(MCInst1_MC3_r2Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst1_MC3_r2Inst_XORInst_0_1_U1  ( .A(MCInst1_MC3_v0_2 [1]), .B(
        MCInst1_MC3_v1_2 [1]), .Z(MCInst1_MC3_r2Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst1_MC3_r2Inst_XORInst_0_2_U3  ( .A(
        MCInst1_MC3_r2Inst_XORInst_0_2_n5 ), .B(
        MCInst1_MC3_r2Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[18]) );
  XNOR2_X1 MCInst1_MC3_r2Inst_XORInst_0_2_U2  ( .A(MCInst1_MC3_v3_2 [2]), 
        .B(MCInst1_MC3_v2_2 [2]), .ZN(MCInst1_MC3_r2Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst1_MC3_r2Inst_XORInst_0_2_U1  ( .A(MCInst1_MC3_v0_2 [2]), .B(
        MCInst1_MC3_v1_2 [2]), .Z(MCInst1_MC3_r2Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst1_MC3_r2Inst_XORInst_0_3_U3  ( .A(
        MCInst1_MC3_r2Inst_XORInst_0_3_n5 ), .B(
        MCInst1_MC3_r2Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[19]) );
  XNOR2_X1 MCInst1_MC3_r2Inst_XORInst_0_3_U2  ( .A(MCInst1_MC3_v3_2 [3]), 
        .B(MCInst1_MC3_v2_2 [3]), .ZN(MCInst1_MC3_r2Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst1_MC3_r2Inst_XORInst_0_3_U1  ( .A(MCInst1_MC3_v0_2 [3]), .B(
        MCInst1_MC3_v1_2 [3]), .Z(MCInst1_MC3_r2Inst_XORInst_0_3_n5 ) );
  XNOR2_X1 MCInst1_MC3_r3Inst_XORInst_0_0_U3  ( .A(
        MCInst1_MC3_r3Inst_XORInst_0_0_n5 ), .B(
        MCInst1_MC3_r3Inst_XORInst_0_0_n4 ), .ZN(Ciphertext[0]) );
  XNOR2_X1 MCInst1_MC3_r3Inst_XORInst_0_0_U2  ( .A(MCInst1_MC3_v3_3 [0]), 
        .B(MCInst1_MC3_v2_3 [0]), .ZN(MCInst1_MC3_r3Inst_XORInst_0_0_n4 ) );
  XOR2_X1 MCInst1_MC3_r3Inst_XORInst_0_0_U1  ( .A(MCInst1_MC3_v0_3 [0]), .B(
        MCInst1_MC3_v1_3 [0]), .Z(MCInst1_MC3_r3Inst_XORInst_0_0_n5 ) );
  XNOR2_X1 MCInst1_MC3_r3Inst_XORInst_0_1_U3  ( .A(
        MCInst1_MC3_r3Inst_XORInst_0_1_n5 ), .B(
        MCInst1_MC3_r3Inst_XORInst_0_1_n4 ), .ZN(Ciphertext[1]) );
  XNOR2_X1 MCInst1_MC3_r3Inst_XORInst_0_1_U2  ( .A(MCInst1_MC3_v3_3 [1]), 
        .B(MCInst1_MC3_v2_3 [1]), .ZN(MCInst1_MC3_r3Inst_XORInst_0_1_n4 ) );
  XOR2_X1 MCInst1_MC3_r3Inst_XORInst_0_1_U1  ( .A(MCInst1_MC3_v0_3 [1]), .B(
        MCInst1_MC3_v1_3 [1]), .Z(MCInst1_MC3_r3Inst_XORInst_0_1_n5 ) );
  XNOR2_X1 MCInst1_MC3_r3Inst_XORInst_0_2_U3  ( .A(
        MCInst1_MC3_r3Inst_XORInst_0_2_n5 ), .B(
        MCInst1_MC3_r3Inst_XORInst_0_2_n4 ), .ZN(Ciphertext[2]) );
  XNOR2_X1 MCInst1_MC3_r3Inst_XORInst_0_2_U2  ( .A(MCInst1_MC3_v3_3 [2]), 
        .B(MCInst1_MC3_v2_3 [2]), .ZN(MCInst1_MC3_r3Inst_XORInst_0_2_n4 ) );
  XOR2_X1 MCInst1_MC3_r3Inst_XORInst_0_2_U1  ( .A(MCInst1_MC3_v0_0 [3]), .B(
        MCInst1_MC3_v1_3 [2]), .Z(MCInst1_MC3_r3Inst_XORInst_0_2_n5 ) );
  XNOR2_X1 MCInst1_MC3_r3Inst_XORInst_0_3_U3  ( .A(
        MCInst1_MC3_r3Inst_XORInst_0_3_n5 ), .B(
        MCInst1_MC3_r3Inst_XORInst_0_3_n4 ), .ZN(Ciphertext[3]) );
  XNOR2_X1 MCInst1_MC3_r3Inst_XORInst_0_3_U2  ( .A(MCInst1_MC3_v3_3 [3]), 
        .B(MCInst1_MC3_v2_3 [3]), .ZN(MCInst1_MC3_r3Inst_XORInst_0_3_n4 ) );
  XOR2_X1 MCInst1_MC3_r3Inst_XORInst_0_3_U1  ( .A(MCInst1_MC3_v0_3 [3]), .B(
        MCInst1_MC3_v1_3 [3]), .Z(MCInst1_MC3_r3Inst_XORInst_0_3_n5 ) );
endmodule

